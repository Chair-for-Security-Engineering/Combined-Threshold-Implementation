// Generator : SpinalHDL v1.7.3    git head : aeaeece704fe43c766e0d36a93f2ecbb8a9f2003
// Component : AES_Round
// Git hash  : db593c14fe8e83f0a4a5d43cf13325e631d65148

`timescale 1ns/1ps

module Round_AES_TI_d1 (
  input      [0:0]    port_state_in_0_0_0,
  input      [0:0]    port_state_in_0_0_1,
  input      [0:0]    port_state_in_0_0_2,
  input      [0:0]    port_state_in_0_0_3,
  input      [0:0]    port_state_in_0_0_4,
  input      [0:0]    port_state_in_0_0_5,
  input      [0:0]    port_state_in_0_0_6,
  input      [0:0]    port_state_in_0_0_7,
  input      [0:0]    port_state_in_0_1_0,
  input      [0:0]    port_state_in_0_1_1,
  input      [0:0]    port_state_in_0_1_2,
  input      [0:0]    port_state_in_0_1_3,
  input      [0:0]    port_state_in_0_1_4,
  input      [0:0]    port_state_in_0_1_5,
  input      [0:0]    port_state_in_0_1_6,
  input      [0:0]    port_state_in_0_1_7,
  input      [0:0]    port_state_in_0_2_0,
  input      [0:0]    port_state_in_0_2_1,
  input      [0:0]    port_state_in_0_2_2,
  input      [0:0]    port_state_in_0_2_3,
  input      [0:0]    port_state_in_0_2_4,
  input      [0:0]    port_state_in_0_2_5,
  input      [0:0]    port_state_in_0_2_6,
  input      [0:0]    port_state_in_0_2_7,
  input      [0:0]    port_state_in_0_3_0,
  input      [0:0]    port_state_in_0_3_1,
  input      [0:0]    port_state_in_0_3_2,
  input      [0:0]    port_state_in_0_3_3,
  input      [0:0]    port_state_in_0_3_4,
  input      [0:0]    port_state_in_0_3_5,
  input      [0:0]    port_state_in_0_3_6,
  input      [0:0]    port_state_in_0_3_7,
  input      [0:0]    port_state_in_1_0_0,
  input      [0:0]    port_state_in_1_0_1,
  input      [0:0]    port_state_in_1_0_2,
  input      [0:0]    port_state_in_1_0_3,
  input      [0:0]    port_state_in_1_0_4,
  input      [0:0]    port_state_in_1_0_5,
  input      [0:0]    port_state_in_1_0_6,
  input      [0:0]    port_state_in_1_0_7,
  input      [0:0]    port_state_in_1_1_0,
  input      [0:0]    port_state_in_1_1_1,
  input      [0:0]    port_state_in_1_1_2,
  input      [0:0]    port_state_in_1_1_3,
  input      [0:0]    port_state_in_1_1_4,
  input      [0:0]    port_state_in_1_1_5,
  input      [0:0]    port_state_in_1_1_6,
  input      [0:0]    port_state_in_1_1_7,
  input      [0:0]    port_state_in_1_2_0,
  input      [0:0]    port_state_in_1_2_1,
  input      [0:0]    port_state_in_1_2_2,
  input      [0:0]    port_state_in_1_2_3,
  input      [0:0]    port_state_in_1_2_4,
  input      [0:0]    port_state_in_1_2_5,
  input      [0:0]    port_state_in_1_2_6,
  input      [0:0]    port_state_in_1_2_7,
  input      [0:0]    port_state_in_1_3_0,
  input      [0:0]    port_state_in_1_3_1,
  input      [0:0]    port_state_in_1_3_2,
  input      [0:0]    port_state_in_1_3_3,
  input      [0:0]    port_state_in_1_3_4,
  input      [0:0]    port_state_in_1_3_5,
  input      [0:0]    port_state_in_1_3_6,
  input      [0:0]    port_state_in_1_3_7,
  input      [0:0]    port_state_in_2_0_0,
  input      [0:0]    port_state_in_2_0_1,
  input      [0:0]    port_state_in_2_0_2,
  input      [0:0]    port_state_in_2_0_3,
  input      [0:0]    port_state_in_2_0_4,
  input      [0:0]    port_state_in_2_0_5,
  input      [0:0]    port_state_in_2_0_6,
  input      [0:0]    port_state_in_2_0_7,
  input      [0:0]    port_state_in_2_1_0,
  input      [0:0]    port_state_in_2_1_1,
  input      [0:0]    port_state_in_2_1_2,
  input      [0:0]    port_state_in_2_1_3,
  input      [0:0]    port_state_in_2_1_4,
  input      [0:0]    port_state_in_2_1_5,
  input      [0:0]    port_state_in_2_1_6,
  input      [0:0]    port_state_in_2_1_7,
  input      [0:0]    port_state_in_2_2_0,
  input      [0:0]    port_state_in_2_2_1,
  input      [0:0]    port_state_in_2_2_2,
  input      [0:0]    port_state_in_2_2_3,
  input      [0:0]    port_state_in_2_2_4,
  input      [0:0]    port_state_in_2_2_5,
  input      [0:0]    port_state_in_2_2_6,
  input      [0:0]    port_state_in_2_2_7,
  input      [0:0]    port_state_in_2_3_0,
  input      [0:0]    port_state_in_2_3_1,
  input      [0:0]    port_state_in_2_3_2,
  input      [0:0]    port_state_in_2_3_3,
  input      [0:0]    port_state_in_2_3_4,
  input      [0:0]    port_state_in_2_3_5,
  input      [0:0]    port_state_in_2_3_6,
  input      [0:0]    port_state_in_2_3_7,
  input      [0:0]    port_state_in_3_0_0,
  input      [0:0]    port_state_in_3_0_1,
  input      [0:0]    port_state_in_3_0_2,
  input      [0:0]    port_state_in_3_0_3,
  input      [0:0]    port_state_in_3_0_4,
  input      [0:0]    port_state_in_3_0_5,
  input      [0:0]    port_state_in_3_0_6,
  input      [0:0]    port_state_in_3_0_7,
  input      [0:0]    port_state_in_3_1_0,
  input      [0:0]    port_state_in_3_1_1,
  input      [0:0]    port_state_in_3_1_2,
  input      [0:0]    port_state_in_3_1_3,
  input      [0:0]    port_state_in_3_1_4,
  input      [0:0]    port_state_in_3_1_5,
  input      [0:0]    port_state_in_3_1_6,
  input      [0:0]    port_state_in_3_1_7,
  input      [0:0]    port_state_in_3_2_0,
  input      [0:0]    port_state_in_3_2_1,
  input      [0:0]    port_state_in_3_2_2,
  input      [0:0]    port_state_in_3_2_3,
  input      [0:0]    port_state_in_3_2_4,
  input      [0:0]    port_state_in_3_2_5,
  input      [0:0]    port_state_in_3_2_6,
  input      [0:0]    port_state_in_3_2_7,
  input      [0:0]    port_state_in_3_3_0,
  input      [0:0]    port_state_in_3_3_1,
  input      [0:0]    port_state_in_3_3_2,
  input      [0:0]    port_state_in_3_3_3,
  input      [0:0]    port_state_in_3_3_4,
  input      [0:0]    port_state_in_3_3_5,
  input      [0:0]    port_state_in_3_3_6,
  input      [0:0]    port_state_in_3_3_7,
  input      [0:0]    port_state_in_4_0_0,
  input      [0:0]    port_state_in_4_0_1,
  input      [0:0]    port_state_in_4_0_2,
  input      [0:0]    port_state_in_4_0_3,
  input      [0:0]    port_state_in_4_0_4,
  input      [0:0]    port_state_in_4_0_5,
  input      [0:0]    port_state_in_4_0_6,
  input      [0:0]    port_state_in_4_0_7,
  input      [0:0]    port_state_in_4_1_0,
  input      [0:0]    port_state_in_4_1_1,
  input      [0:0]    port_state_in_4_1_2,
  input      [0:0]    port_state_in_4_1_3,
  input      [0:0]    port_state_in_4_1_4,
  input      [0:0]    port_state_in_4_1_5,
  input      [0:0]    port_state_in_4_1_6,
  input      [0:0]    port_state_in_4_1_7,
  input      [0:0]    port_state_in_4_2_0,
  input      [0:0]    port_state_in_4_2_1,
  input      [0:0]    port_state_in_4_2_2,
  input      [0:0]    port_state_in_4_2_3,
  input      [0:0]    port_state_in_4_2_4,
  input      [0:0]    port_state_in_4_2_5,
  input      [0:0]    port_state_in_4_2_6,
  input      [0:0]    port_state_in_4_2_7,
  input      [0:0]    port_state_in_4_3_0,
  input      [0:0]    port_state_in_4_3_1,
  input      [0:0]    port_state_in_4_3_2,
  input      [0:0]    port_state_in_4_3_3,
  input      [0:0]    port_state_in_4_3_4,
  input      [0:0]    port_state_in_4_3_5,
  input      [0:0]    port_state_in_4_3_6,
  input      [0:0]    port_state_in_4_3_7,
  input      [0:0]    port_state_in_5_0_0,
  input      [0:0]    port_state_in_5_0_1,
  input      [0:0]    port_state_in_5_0_2,
  input      [0:0]    port_state_in_5_0_3,
  input      [0:0]    port_state_in_5_0_4,
  input      [0:0]    port_state_in_5_0_5,
  input      [0:0]    port_state_in_5_0_6,
  input      [0:0]    port_state_in_5_0_7,
  input      [0:0]    port_state_in_5_1_0,
  input      [0:0]    port_state_in_5_1_1,
  input      [0:0]    port_state_in_5_1_2,
  input      [0:0]    port_state_in_5_1_3,
  input      [0:0]    port_state_in_5_1_4,
  input      [0:0]    port_state_in_5_1_5,
  input      [0:0]    port_state_in_5_1_6,
  input      [0:0]    port_state_in_5_1_7,
  input      [0:0]    port_state_in_5_2_0,
  input      [0:0]    port_state_in_5_2_1,
  input      [0:0]    port_state_in_5_2_2,
  input      [0:0]    port_state_in_5_2_3,
  input      [0:0]    port_state_in_5_2_4,
  input      [0:0]    port_state_in_5_2_5,
  input      [0:0]    port_state_in_5_2_6,
  input      [0:0]    port_state_in_5_2_7,
  input      [0:0]    port_state_in_5_3_0,
  input      [0:0]    port_state_in_5_3_1,
  input      [0:0]    port_state_in_5_3_2,
  input      [0:0]    port_state_in_5_3_3,
  input      [0:0]    port_state_in_5_3_4,
  input      [0:0]    port_state_in_5_3_5,
  input      [0:0]    port_state_in_5_3_6,
  input      [0:0]    port_state_in_5_3_7,
  input      [0:0]    port_state_in_6_0_0,
  input      [0:0]    port_state_in_6_0_1,
  input      [0:0]    port_state_in_6_0_2,
  input      [0:0]    port_state_in_6_0_3,
  input      [0:0]    port_state_in_6_0_4,
  input      [0:0]    port_state_in_6_0_5,
  input      [0:0]    port_state_in_6_0_6,
  input      [0:0]    port_state_in_6_0_7,
  input      [0:0]    port_state_in_6_1_0,
  input      [0:0]    port_state_in_6_1_1,
  input      [0:0]    port_state_in_6_1_2,
  input      [0:0]    port_state_in_6_1_3,
  input      [0:0]    port_state_in_6_1_4,
  input      [0:0]    port_state_in_6_1_5,
  input      [0:0]    port_state_in_6_1_6,
  input      [0:0]    port_state_in_6_1_7,
  input      [0:0]    port_state_in_6_2_0,
  input      [0:0]    port_state_in_6_2_1,
  input      [0:0]    port_state_in_6_2_2,
  input      [0:0]    port_state_in_6_2_3,
  input      [0:0]    port_state_in_6_2_4,
  input      [0:0]    port_state_in_6_2_5,
  input      [0:0]    port_state_in_6_2_6,
  input      [0:0]    port_state_in_6_2_7,
  input      [0:0]    port_state_in_6_3_0,
  input      [0:0]    port_state_in_6_3_1,
  input      [0:0]    port_state_in_6_3_2,
  input      [0:0]    port_state_in_6_3_3,
  input      [0:0]    port_state_in_6_3_4,
  input      [0:0]    port_state_in_6_3_5,
  input      [0:0]    port_state_in_6_3_6,
  input      [0:0]    port_state_in_6_3_7,
  input      [0:0]    port_state_in_7_0_0,
  input      [0:0]    port_state_in_7_0_1,
  input      [0:0]    port_state_in_7_0_2,
  input      [0:0]    port_state_in_7_0_3,
  input      [0:0]    port_state_in_7_0_4,
  input      [0:0]    port_state_in_7_0_5,
  input      [0:0]    port_state_in_7_0_6,
  input      [0:0]    port_state_in_7_0_7,
  input      [0:0]    port_state_in_7_1_0,
  input      [0:0]    port_state_in_7_1_1,
  input      [0:0]    port_state_in_7_1_2,
  input      [0:0]    port_state_in_7_1_3,
  input      [0:0]    port_state_in_7_1_4,
  input      [0:0]    port_state_in_7_1_5,
  input      [0:0]    port_state_in_7_1_6,
  input      [0:0]    port_state_in_7_1_7,
  input      [0:0]    port_state_in_7_2_0,
  input      [0:0]    port_state_in_7_2_1,
  input      [0:0]    port_state_in_7_2_2,
  input      [0:0]    port_state_in_7_2_3,
  input      [0:0]    port_state_in_7_2_4,
  input      [0:0]    port_state_in_7_2_5,
  input      [0:0]    port_state_in_7_2_6,
  input      [0:0]    port_state_in_7_2_7,
  input      [0:0]    port_state_in_7_3_0,
  input      [0:0]    port_state_in_7_3_1,
  input      [0:0]    port_state_in_7_3_2,
  input      [0:0]    port_state_in_7_3_3,
  input      [0:0]    port_state_in_7_3_4,
  input      [0:0]    port_state_in_7_3_5,
  input      [0:0]    port_state_in_7_3_6,
  input      [0:0]    port_state_in_7_3_7,
  input      [0:0]    port_state_in_8_0_0,
  input      [0:0]    port_state_in_8_0_1,
  input      [0:0]    port_state_in_8_0_2,
  input      [0:0]    port_state_in_8_0_3,
  input      [0:0]    port_state_in_8_0_4,
  input      [0:0]    port_state_in_8_0_5,
  input      [0:0]    port_state_in_8_0_6,
  input      [0:0]    port_state_in_8_0_7,
  input      [0:0]    port_state_in_8_1_0,
  input      [0:0]    port_state_in_8_1_1,
  input      [0:0]    port_state_in_8_1_2,
  input      [0:0]    port_state_in_8_1_3,
  input      [0:0]    port_state_in_8_1_4,
  input      [0:0]    port_state_in_8_1_5,
  input      [0:0]    port_state_in_8_1_6,
  input      [0:0]    port_state_in_8_1_7,
  input      [0:0]    port_state_in_8_2_0,
  input      [0:0]    port_state_in_8_2_1,
  input      [0:0]    port_state_in_8_2_2,
  input      [0:0]    port_state_in_8_2_3,
  input      [0:0]    port_state_in_8_2_4,
  input      [0:0]    port_state_in_8_2_5,
  input      [0:0]    port_state_in_8_2_6,
  input      [0:0]    port_state_in_8_2_7,
  input      [0:0]    port_state_in_8_3_0,
  input      [0:0]    port_state_in_8_3_1,
  input      [0:0]    port_state_in_8_3_2,
  input      [0:0]    port_state_in_8_3_3,
  input      [0:0]    port_state_in_8_3_4,
  input      [0:0]    port_state_in_8_3_5,
  input      [0:0]    port_state_in_8_3_6,
  input      [0:0]    port_state_in_8_3_7,
  input      [0:0]    port_state_in_9_0_0,
  input      [0:0]    port_state_in_9_0_1,
  input      [0:0]    port_state_in_9_0_2,
  input      [0:0]    port_state_in_9_0_3,
  input      [0:0]    port_state_in_9_0_4,
  input      [0:0]    port_state_in_9_0_5,
  input      [0:0]    port_state_in_9_0_6,
  input      [0:0]    port_state_in_9_0_7,
  input      [0:0]    port_state_in_9_1_0,
  input      [0:0]    port_state_in_9_1_1,
  input      [0:0]    port_state_in_9_1_2,
  input      [0:0]    port_state_in_9_1_3,
  input      [0:0]    port_state_in_9_1_4,
  input      [0:0]    port_state_in_9_1_5,
  input      [0:0]    port_state_in_9_1_6,
  input      [0:0]    port_state_in_9_1_7,
  input      [0:0]    port_state_in_9_2_0,
  input      [0:0]    port_state_in_9_2_1,
  input      [0:0]    port_state_in_9_2_2,
  input      [0:0]    port_state_in_9_2_3,
  input      [0:0]    port_state_in_9_2_4,
  input      [0:0]    port_state_in_9_2_5,
  input      [0:0]    port_state_in_9_2_6,
  input      [0:0]    port_state_in_9_2_7,
  input      [0:0]    port_state_in_9_3_0,
  input      [0:0]    port_state_in_9_3_1,
  input      [0:0]    port_state_in_9_3_2,
  input      [0:0]    port_state_in_9_3_3,
  input      [0:0]    port_state_in_9_3_4,
  input      [0:0]    port_state_in_9_3_5,
  input      [0:0]    port_state_in_9_3_6,
  input      [0:0]    port_state_in_9_3_7,
  input      [0:0]    port_state_in_10_0_0,
  input      [0:0]    port_state_in_10_0_1,
  input      [0:0]    port_state_in_10_0_2,
  input      [0:0]    port_state_in_10_0_3,
  input      [0:0]    port_state_in_10_0_4,
  input      [0:0]    port_state_in_10_0_5,
  input      [0:0]    port_state_in_10_0_6,
  input      [0:0]    port_state_in_10_0_7,
  input      [0:0]    port_state_in_10_1_0,
  input      [0:0]    port_state_in_10_1_1,
  input      [0:0]    port_state_in_10_1_2,
  input      [0:0]    port_state_in_10_1_3,
  input      [0:0]    port_state_in_10_1_4,
  input      [0:0]    port_state_in_10_1_5,
  input      [0:0]    port_state_in_10_1_6,
  input      [0:0]    port_state_in_10_1_7,
  input      [0:0]    port_state_in_10_2_0,
  input      [0:0]    port_state_in_10_2_1,
  input      [0:0]    port_state_in_10_2_2,
  input      [0:0]    port_state_in_10_2_3,
  input      [0:0]    port_state_in_10_2_4,
  input      [0:0]    port_state_in_10_2_5,
  input      [0:0]    port_state_in_10_2_6,
  input      [0:0]    port_state_in_10_2_7,
  input      [0:0]    port_state_in_10_3_0,
  input      [0:0]    port_state_in_10_3_1,
  input      [0:0]    port_state_in_10_3_2,
  input      [0:0]    port_state_in_10_3_3,
  input      [0:0]    port_state_in_10_3_4,
  input      [0:0]    port_state_in_10_3_5,
  input      [0:0]    port_state_in_10_3_6,
  input      [0:0]    port_state_in_10_3_7,
  input      [0:0]    port_state_in_11_0_0,
  input      [0:0]    port_state_in_11_0_1,
  input      [0:0]    port_state_in_11_0_2,
  input      [0:0]    port_state_in_11_0_3,
  input      [0:0]    port_state_in_11_0_4,
  input      [0:0]    port_state_in_11_0_5,
  input      [0:0]    port_state_in_11_0_6,
  input      [0:0]    port_state_in_11_0_7,
  input      [0:0]    port_state_in_11_1_0,
  input      [0:0]    port_state_in_11_1_1,
  input      [0:0]    port_state_in_11_1_2,
  input      [0:0]    port_state_in_11_1_3,
  input      [0:0]    port_state_in_11_1_4,
  input      [0:0]    port_state_in_11_1_5,
  input      [0:0]    port_state_in_11_1_6,
  input      [0:0]    port_state_in_11_1_7,
  input      [0:0]    port_state_in_11_2_0,
  input      [0:0]    port_state_in_11_2_1,
  input      [0:0]    port_state_in_11_2_2,
  input      [0:0]    port_state_in_11_2_3,
  input      [0:0]    port_state_in_11_2_4,
  input      [0:0]    port_state_in_11_2_5,
  input      [0:0]    port_state_in_11_2_6,
  input      [0:0]    port_state_in_11_2_7,
  input      [0:0]    port_state_in_11_3_0,
  input      [0:0]    port_state_in_11_3_1,
  input      [0:0]    port_state_in_11_3_2,
  input      [0:0]    port_state_in_11_3_3,
  input      [0:0]    port_state_in_11_3_4,
  input      [0:0]    port_state_in_11_3_5,
  input      [0:0]    port_state_in_11_3_6,
  input      [0:0]    port_state_in_11_3_7,
  input      [0:0]    port_state_in_12_0_0,
  input      [0:0]    port_state_in_12_0_1,
  input      [0:0]    port_state_in_12_0_2,
  input      [0:0]    port_state_in_12_0_3,
  input      [0:0]    port_state_in_12_0_4,
  input      [0:0]    port_state_in_12_0_5,
  input      [0:0]    port_state_in_12_0_6,
  input      [0:0]    port_state_in_12_0_7,
  input      [0:0]    port_state_in_12_1_0,
  input      [0:0]    port_state_in_12_1_1,
  input      [0:0]    port_state_in_12_1_2,
  input      [0:0]    port_state_in_12_1_3,
  input      [0:0]    port_state_in_12_1_4,
  input      [0:0]    port_state_in_12_1_5,
  input      [0:0]    port_state_in_12_1_6,
  input      [0:0]    port_state_in_12_1_7,
  input      [0:0]    port_state_in_12_2_0,
  input      [0:0]    port_state_in_12_2_1,
  input      [0:0]    port_state_in_12_2_2,
  input      [0:0]    port_state_in_12_2_3,
  input      [0:0]    port_state_in_12_2_4,
  input      [0:0]    port_state_in_12_2_5,
  input      [0:0]    port_state_in_12_2_6,
  input      [0:0]    port_state_in_12_2_7,
  input      [0:0]    port_state_in_12_3_0,
  input      [0:0]    port_state_in_12_3_1,
  input      [0:0]    port_state_in_12_3_2,
  input      [0:0]    port_state_in_12_3_3,
  input      [0:0]    port_state_in_12_3_4,
  input      [0:0]    port_state_in_12_3_5,
  input      [0:0]    port_state_in_12_3_6,
  input      [0:0]    port_state_in_12_3_7,
  input      [0:0]    port_state_in_13_0_0,
  input      [0:0]    port_state_in_13_0_1,
  input      [0:0]    port_state_in_13_0_2,
  input      [0:0]    port_state_in_13_0_3,
  input      [0:0]    port_state_in_13_0_4,
  input      [0:0]    port_state_in_13_0_5,
  input      [0:0]    port_state_in_13_0_6,
  input      [0:0]    port_state_in_13_0_7,
  input      [0:0]    port_state_in_13_1_0,
  input      [0:0]    port_state_in_13_1_1,
  input      [0:0]    port_state_in_13_1_2,
  input      [0:0]    port_state_in_13_1_3,
  input      [0:0]    port_state_in_13_1_4,
  input      [0:0]    port_state_in_13_1_5,
  input      [0:0]    port_state_in_13_1_6,
  input      [0:0]    port_state_in_13_1_7,
  input      [0:0]    port_state_in_13_2_0,
  input      [0:0]    port_state_in_13_2_1,
  input      [0:0]    port_state_in_13_2_2,
  input      [0:0]    port_state_in_13_2_3,
  input      [0:0]    port_state_in_13_2_4,
  input      [0:0]    port_state_in_13_2_5,
  input      [0:0]    port_state_in_13_2_6,
  input      [0:0]    port_state_in_13_2_7,
  input      [0:0]    port_state_in_13_3_0,
  input      [0:0]    port_state_in_13_3_1,
  input      [0:0]    port_state_in_13_3_2,
  input      [0:0]    port_state_in_13_3_3,
  input      [0:0]    port_state_in_13_3_4,
  input      [0:0]    port_state_in_13_3_5,
  input      [0:0]    port_state_in_13_3_6,
  input      [0:0]    port_state_in_13_3_7,
  input      [0:0]    port_state_in_14_0_0,
  input      [0:0]    port_state_in_14_0_1,
  input      [0:0]    port_state_in_14_0_2,
  input      [0:0]    port_state_in_14_0_3,
  input      [0:0]    port_state_in_14_0_4,
  input      [0:0]    port_state_in_14_0_5,
  input      [0:0]    port_state_in_14_0_6,
  input      [0:0]    port_state_in_14_0_7,
  input      [0:0]    port_state_in_14_1_0,
  input      [0:0]    port_state_in_14_1_1,
  input      [0:0]    port_state_in_14_1_2,
  input      [0:0]    port_state_in_14_1_3,
  input      [0:0]    port_state_in_14_1_4,
  input      [0:0]    port_state_in_14_1_5,
  input      [0:0]    port_state_in_14_1_6,
  input      [0:0]    port_state_in_14_1_7,
  input      [0:0]    port_state_in_14_2_0,
  input      [0:0]    port_state_in_14_2_1,
  input      [0:0]    port_state_in_14_2_2,
  input      [0:0]    port_state_in_14_2_3,
  input      [0:0]    port_state_in_14_2_4,
  input      [0:0]    port_state_in_14_2_5,
  input      [0:0]    port_state_in_14_2_6,
  input      [0:0]    port_state_in_14_2_7,
  input      [0:0]    port_state_in_14_3_0,
  input      [0:0]    port_state_in_14_3_1,
  input      [0:0]    port_state_in_14_3_2,
  input      [0:0]    port_state_in_14_3_3,
  input      [0:0]    port_state_in_14_3_4,
  input      [0:0]    port_state_in_14_3_5,
  input      [0:0]    port_state_in_14_3_6,
  input      [0:0]    port_state_in_14_3_7,
  input      [0:0]    port_state_in_15_0_0,
  input      [0:0]    port_state_in_15_0_1,
  input      [0:0]    port_state_in_15_0_2,
  input      [0:0]    port_state_in_15_0_3,
  input      [0:0]    port_state_in_15_0_4,
  input      [0:0]    port_state_in_15_0_5,
  input      [0:0]    port_state_in_15_0_6,
  input      [0:0]    port_state_in_15_0_7,
  input      [0:0]    port_state_in_15_1_0,
  input      [0:0]    port_state_in_15_1_1,
  input      [0:0]    port_state_in_15_1_2,
  input      [0:0]    port_state_in_15_1_3,
  input      [0:0]    port_state_in_15_1_4,
  input      [0:0]    port_state_in_15_1_5,
  input      [0:0]    port_state_in_15_1_6,
  input      [0:0]    port_state_in_15_1_7,
  input      [0:0]    port_state_in_15_2_0,
  input      [0:0]    port_state_in_15_2_1,
  input      [0:0]    port_state_in_15_2_2,
  input      [0:0]    port_state_in_15_2_3,
  input      [0:0]    port_state_in_15_2_4,
  input      [0:0]    port_state_in_15_2_5,
  input      [0:0]    port_state_in_15_2_6,
  input      [0:0]    port_state_in_15_2_7,
  input      [0:0]    port_state_in_15_3_0,
  input      [0:0]    port_state_in_15_3_1,
  input      [0:0]    port_state_in_15_3_2,
  input      [0:0]    port_state_in_15_3_3,
  input      [0:0]    port_state_in_15_3_4,
  input      [0:0]    port_state_in_15_3_5,
  input      [0:0]    port_state_in_15_3_6,
  input      [0:0]    port_state_in_15_3_7,
  input      [0:0]    port_key_0_0_0,
  input      [0:0]    port_key_0_0_1,
  input      [0:0]    port_key_0_0_2,
  input      [0:0]    port_key_0_0_3,
  input      [0:0]    port_key_0_0_4,
  input      [0:0]    port_key_0_0_5,
  input      [0:0]    port_key_0_0_6,
  input      [0:0]    port_key_0_0_7,
  input      [0:0]    port_key_0_1_0,
  input      [0:0]    port_key_0_1_1,
  input      [0:0]    port_key_0_1_2,
  input      [0:0]    port_key_0_1_3,
  input      [0:0]    port_key_0_1_4,
  input      [0:0]    port_key_0_1_5,
  input      [0:0]    port_key_0_1_6,
  input      [0:0]    port_key_0_1_7,
  input      [0:0]    port_key_0_2_0,
  input      [0:0]    port_key_0_2_1,
  input      [0:0]    port_key_0_2_2,
  input      [0:0]    port_key_0_2_3,
  input      [0:0]    port_key_0_2_4,
  input      [0:0]    port_key_0_2_5,
  input      [0:0]    port_key_0_2_6,
  input      [0:0]    port_key_0_2_7,
  input      [0:0]    port_key_0_3_0,
  input      [0:0]    port_key_0_3_1,
  input      [0:0]    port_key_0_3_2,
  input      [0:0]    port_key_0_3_3,
  input      [0:0]    port_key_0_3_4,
  input      [0:0]    port_key_0_3_5,
  input      [0:0]    port_key_0_3_6,
  input      [0:0]    port_key_0_3_7,
  input      [0:0]    port_key_1_0_0,
  input      [0:0]    port_key_1_0_1,
  input      [0:0]    port_key_1_0_2,
  input      [0:0]    port_key_1_0_3,
  input      [0:0]    port_key_1_0_4,
  input      [0:0]    port_key_1_0_5,
  input      [0:0]    port_key_1_0_6,
  input      [0:0]    port_key_1_0_7,
  input      [0:0]    port_key_1_1_0,
  input      [0:0]    port_key_1_1_1,
  input      [0:0]    port_key_1_1_2,
  input      [0:0]    port_key_1_1_3,
  input      [0:0]    port_key_1_1_4,
  input      [0:0]    port_key_1_1_5,
  input      [0:0]    port_key_1_1_6,
  input      [0:0]    port_key_1_1_7,
  input      [0:0]    port_key_1_2_0,
  input      [0:0]    port_key_1_2_1,
  input      [0:0]    port_key_1_2_2,
  input      [0:0]    port_key_1_2_3,
  input      [0:0]    port_key_1_2_4,
  input      [0:0]    port_key_1_2_5,
  input      [0:0]    port_key_1_2_6,
  input      [0:0]    port_key_1_2_7,
  input      [0:0]    port_key_1_3_0,
  input      [0:0]    port_key_1_3_1,
  input      [0:0]    port_key_1_3_2,
  input      [0:0]    port_key_1_3_3,
  input      [0:0]    port_key_1_3_4,
  input      [0:0]    port_key_1_3_5,
  input      [0:0]    port_key_1_3_6,
  input      [0:0]    port_key_1_3_7,
  input      [0:0]    port_key_2_0_0,
  input      [0:0]    port_key_2_0_1,
  input      [0:0]    port_key_2_0_2,
  input      [0:0]    port_key_2_0_3,
  input      [0:0]    port_key_2_0_4,
  input      [0:0]    port_key_2_0_5,
  input      [0:0]    port_key_2_0_6,
  input      [0:0]    port_key_2_0_7,
  input      [0:0]    port_key_2_1_0,
  input      [0:0]    port_key_2_1_1,
  input      [0:0]    port_key_2_1_2,
  input      [0:0]    port_key_2_1_3,
  input      [0:0]    port_key_2_1_4,
  input      [0:0]    port_key_2_1_5,
  input      [0:0]    port_key_2_1_6,
  input      [0:0]    port_key_2_1_7,
  input      [0:0]    port_key_2_2_0,
  input      [0:0]    port_key_2_2_1,
  input      [0:0]    port_key_2_2_2,
  input      [0:0]    port_key_2_2_3,
  input      [0:0]    port_key_2_2_4,
  input      [0:0]    port_key_2_2_5,
  input      [0:0]    port_key_2_2_6,
  input      [0:0]    port_key_2_2_7,
  input      [0:0]    port_key_2_3_0,
  input      [0:0]    port_key_2_3_1,
  input      [0:0]    port_key_2_3_2,
  input      [0:0]    port_key_2_3_3,
  input      [0:0]    port_key_2_3_4,
  input      [0:0]    port_key_2_3_5,
  input      [0:0]    port_key_2_3_6,
  input      [0:0]    port_key_2_3_7,
  input      [0:0]    port_key_3_0_0,
  input      [0:0]    port_key_3_0_1,
  input      [0:0]    port_key_3_0_2,
  input      [0:0]    port_key_3_0_3,
  input      [0:0]    port_key_3_0_4,
  input      [0:0]    port_key_3_0_5,
  input      [0:0]    port_key_3_0_6,
  input      [0:0]    port_key_3_0_7,
  input      [0:0]    port_key_3_1_0,
  input      [0:0]    port_key_3_1_1,
  input      [0:0]    port_key_3_1_2,
  input      [0:0]    port_key_3_1_3,
  input      [0:0]    port_key_3_1_4,
  input      [0:0]    port_key_3_1_5,
  input      [0:0]    port_key_3_1_6,
  input      [0:0]    port_key_3_1_7,
  input      [0:0]    port_key_3_2_0,
  input      [0:0]    port_key_3_2_1,
  input      [0:0]    port_key_3_2_2,
  input      [0:0]    port_key_3_2_3,
  input      [0:0]    port_key_3_2_4,
  input      [0:0]    port_key_3_2_5,
  input      [0:0]    port_key_3_2_6,
  input      [0:0]    port_key_3_2_7,
  input      [0:0]    port_key_3_3_0,
  input      [0:0]    port_key_3_3_1,
  input      [0:0]    port_key_3_3_2,
  input      [0:0]    port_key_3_3_3,
  input      [0:0]    port_key_3_3_4,
  input      [0:0]    port_key_3_3_5,
  input      [0:0]    port_key_3_3_6,
  input      [0:0]    port_key_3_3_7,
  input      [0:0]    port_key_4_0_0,
  input      [0:0]    port_key_4_0_1,
  input      [0:0]    port_key_4_0_2,
  input      [0:0]    port_key_4_0_3,
  input      [0:0]    port_key_4_0_4,
  input      [0:0]    port_key_4_0_5,
  input      [0:0]    port_key_4_0_6,
  input      [0:0]    port_key_4_0_7,
  input      [0:0]    port_key_4_1_0,
  input      [0:0]    port_key_4_1_1,
  input      [0:0]    port_key_4_1_2,
  input      [0:0]    port_key_4_1_3,
  input      [0:0]    port_key_4_1_4,
  input      [0:0]    port_key_4_1_5,
  input      [0:0]    port_key_4_1_6,
  input      [0:0]    port_key_4_1_7,
  input      [0:0]    port_key_4_2_0,
  input      [0:0]    port_key_4_2_1,
  input      [0:0]    port_key_4_2_2,
  input      [0:0]    port_key_4_2_3,
  input      [0:0]    port_key_4_2_4,
  input      [0:0]    port_key_4_2_5,
  input      [0:0]    port_key_4_2_6,
  input      [0:0]    port_key_4_2_7,
  input      [0:0]    port_key_4_3_0,
  input      [0:0]    port_key_4_3_1,
  input      [0:0]    port_key_4_3_2,
  input      [0:0]    port_key_4_3_3,
  input      [0:0]    port_key_4_3_4,
  input      [0:0]    port_key_4_3_5,
  input      [0:0]    port_key_4_3_6,
  input      [0:0]    port_key_4_3_7,
  input      [0:0]    port_key_5_0_0,
  input      [0:0]    port_key_5_0_1,
  input      [0:0]    port_key_5_0_2,
  input      [0:0]    port_key_5_0_3,
  input      [0:0]    port_key_5_0_4,
  input      [0:0]    port_key_5_0_5,
  input      [0:0]    port_key_5_0_6,
  input      [0:0]    port_key_5_0_7,
  input      [0:0]    port_key_5_1_0,
  input      [0:0]    port_key_5_1_1,
  input      [0:0]    port_key_5_1_2,
  input      [0:0]    port_key_5_1_3,
  input      [0:0]    port_key_5_1_4,
  input      [0:0]    port_key_5_1_5,
  input      [0:0]    port_key_5_1_6,
  input      [0:0]    port_key_5_1_7,
  input      [0:0]    port_key_5_2_0,
  input      [0:0]    port_key_5_2_1,
  input      [0:0]    port_key_5_2_2,
  input      [0:0]    port_key_5_2_3,
  input      [0:0]    port_key_5_2_4,
  input      [0:0]    port_key_5_2_5,
  input      [0:0]    port_key_5_2_6,
  input      [0:0]    port_key_5_2_7,
  input      [0:0]    port_key_5_3_0,
  input      [0:0]    port_key_5_3_1,
  input      [0:0]    port_key_5_3_2,
  input      [0:0]    port_key_5_3_3,
  input      [0:0]    port_key_5_3_4,
  input      [0:0]    port_key_5_3_5,
  input      [0:0]    port_key_5_3_6,
  input      [0:0]    port_key_5_3_7,
  input      [0:0]    port_key_6_0_0,
  input      [0:0]    port_key_6_0_1,
  input      [0:0]    port_key_6_0_2,
  input      [0:0]    port_key_6_0_3,
  input      [0:0]    port_key_6_0_4,
  input      [0:0]    port_key_6_0_5,
  input      [0:0]    port_key_6_0_6,
  input      [0:0]    port_key_6_0_7,
  input      [0:0]    port_key_6_1_0,
  input      [0:0]    port_key_6_1_1,
  input      [0:0]    port_key_6_1_2,
  input      [0:0]    port_key_6_1_3,
  input      [0:0]    port_key_6_1_4,
  input      [0:0]    port_key_6_1_5,
  input      [0:0]    port_key_6_1_6,
  input      [0:0]    port_key_6_1_7,
  input      [0:0]    port_key_6_2_0,
  input      [0:0]    port_key_6_2_1,
  input      [0:0]    port_key_6_2_2,
  input      [0:0]    port_key_6_2_3,
  input      [0:0]    port_key_6_2_4,
  input      [0:0]    port_key_6_2_5,
  input      [0:0]    port_key_6_2_6,
  input      [0:0]    port_key_6_2_7,
  input      [0:0]    port_key_6_3_0,
  input      [0:0]    port_key_6_3_1,
  input      [0:0]    port_key_6_3_2,
  input      [0:0]    port_key_6_3_3,
  input      [0:0]    port_key_6_3_4,
  input      [0:0]    port_key_6_3_5,
  input      [0:0]    port_key_6_3_6,
  input      [0:0]    port_key_6_3_7,
  input      [0:0]    port_key_7_0_0,
  input      [0:0]    port_key_7_0_1,
  input      [0:0]    port_key_7_0_2,
  input      [0:0]    port_key_7_0_3,
  input      [0:0]    port_key_7_0_4,
  input      [0:0]    port_key_7_0_5,
  input      [0:0]    port_key_7_0_6,
  input      [0:0]    port_key_7_0_7,
  input      [0:0]    port_key_7_1_0,
  input      [0:0]    port_key_7_1_1,
  input      [0:0]    port_key_7_1_2,
  input      [0:0]    port_key_7_1_3,
  input      [0:0]    port_key_7_1_4,
  input      [0:0]    port_key_7_1_5,
  input      [0:0]    port_key_7_1_6,
  input      [0:0]    port_key_7_1_7,
  input      [0:0]    port_key_7_2_0,
  input      [0:0]    port_key_7_2_1,
  input      [0:0]    port_key_7_2_2,
  input      [0:0]    port_key_7_2_3,
  input      [0:0]    port_key_7_2_4,
  input      [0:0]    port_key_7_2_5,
  input      [0:0]    port_key_7_2_6,
  input      [0:0]    port_key_7_2_7,
  input      [0:0]    port_key_7_3_0,
  input      [0:0]    port_key_7_3_1,
  input      [0:0]    port_key_7_3_2,
  input      [0:0]    port_key_7_3_3,
  input      [0:0]    port_key_7_3_4,
  input      [0:0]    port_key_7_3_5,
  input      [0:0]    port_key_7_3_6,
  input      [0:0]    port_key_7_3_7,
  input      [0:0]    port_key_8_0_0,
  input      [0:0]    port_key_8_0_1,
  input      [0:0]    port_key_8_0_2,
  input      [0:0]    port_key_8_0_3,
  input      [0:0]    port_key_8_0_4,
  input      [0:0]    port_key_8_0_5,
  input      [0:0]    port_key_8_0_6,
  input      [0:0]    port_key_8_0_7,
  input      [0:0]    port_key_8_1_0,
  input      [0:0]    port_key_8_1_1,
  input      [0:0]    port_key_8_1_2,
  input      [0:0]    port_key_8_1_3,
  input      [0:0]    port_key_8_1_4,
  input      [0:0]    port_key_8_1_5,
  input      [0:0]    port_key_8_1_6,
  input      [0:0]    port_key_8_1_7,
  input      [0:0]    port_key_8_2_0,
  input      [0:0]    port_key_8_2_1,
  input      [0:0]    port_key_8_2_2,
  input      [0:0]    port_key_8_2_3,
  input      [0:0]    port_key_8_2_4,
  input      [0:0]    port_key_8_2_5,
  input      [0:0]    port_key_8_2_6,
  input      [0:0]    port_key_8_2_7,
  input      [0:0]    port_key_8_3_0,
  input      [0:0]    port_key_8_3_1,
  input      [0:0]    port_key_8_3_2,
  input      [0:0]    port_key_8_3_3,
  input      [0:0]    port_key_8_3_4,
  input      [0:0]    port_key_8_3_5,
  input      [0:0]    port_key_8_3_6,
  input      [0:0]    port_key_8_3_7,
  input      [0:0]    port_key_9_0_0,
  input      [0:0]    port_key_9_0_1,
  input      [0:0]    port_key_9_0_2,
  input      [0:0]    port_key_9_0_3,
  input      [0:0]    port_key_9_0_4,
  input      [0:0]    port_key_9_0_5,
  input      [0:0]    port_key_9_0_6,
  input      [0:0]    port_key_9_0_7,
  input      [0:0]    port_key_9_1_0,
  input      [0:0]    port_key_9_1_1,
  input      [0:0]    port_key_9_1_2,
  input      [0:0]    port_key_9_1_3,
  input      [0:0]    port_key_9_1_4,
  input      [0:0]    port_key_9_1_5,
  input      [0:0]    port_key_9_1_6,
  input      [0:0]    port_key_9_1_7,
  input      [0:0]    port_key_9_2_0,
  input      [0:0]    port_key_9_2_1,
  input      [0:0]    port_key_9_2_2,
  input      [0:0]    port_key_9_2_3,
  input      [0:0]    port_key_9_2_4,
  input      [0:0]    port_key_9_2_5,
  input      [0:0]    port_key_9_2_6,
  input      [0:0]    port_key_9_2_7,
  input      [0:0]    port_key_9_3_0,
  input      [0:0]    port_key_9_3_1,
  input      [0:0]    port_key_9_3_2,
  input      [0:0]    port_key_9_3_3,
  input      [0:0]    port_key_9_3_4,
  input      [0:0]    port_key_9_3_5,
  input      [0:0]    port_key_9_3_6,
  input      [0:0]    port_key_9_3_7,
  input      [0:0]    port_key_10_0_0,
  input      [0:0]    port_key_10_0_1,
  input      [0:0]    port_key_10_0_2,
  input      [0:0]    port_key_10_0_3,
  input      [0:0]    port_key_10_0_4,
  input      [0:0]    port_key_10_0_5,
  input      [0:0]    port_key_10_0_6,
  input      [0:0]    port_key_10_0_7,
  input      [0:0]    port_key_10_1_0,
  input      [0:0]    port_key_10_1_1,
  input      [0:0]    port_key_10_1_2,
  input      [0:0]    port_key_10_1_3,
  input      [0:0]    port_key_10_1_4,
  input      [0:0]    port_key_10_1_5,
  input      [0:0]    port_key_10_1_6,
  input      [0:0]    port_key_10_1_7,
  input      [0:0]    port_key_10_2_0,
  input      [0:0]    port_key_10_2_1,
  input      [0:0]    port_key_10_2_2,
  input      [0:0]    port_key_10_2_3,
  input      [0:0]    port_key_10_2_4,
  input      [0:0]    port_key_10_2_5,
  input      [0:0]    port_key_10_2_6,
  input      [0:0]    port_key_10_2_7,
  input      [0:0]    port_key_10_3_0,
  input      [0:0]    port_key_10_3_1,
  input      [0:0]    port_key_10_3_2,
  input      [0:0]    port_key_10_3_3,
  input      [0:0]    port_key_10_3_4,
  input      [0:0]    port_key_10_3_5,
  input      [0:0]    port_key_10_3_6,
  input      [0:0]    port_key_10_3_7,
  input      [0:0]    port_key_11_0_0,
  input      [0:0]    port_key_11_0_1,
  input      [0:0]    port_key_11_0_2,
  input      [0:0]    port_key_11_0_3,
  input      [0:0]    port_key_11_0_4,
  input      [0:0]    port_key_11_0_5,
  input      [0:0]    port_key_11_0_6,
  input      [0:0]    port_key_11_0_7,
  input      [0:0]    port_key_11_1_0,
  input      [0:0]    port_key_11_1_1,
  input      [0:0]    port_key_11_1_2,
  input      [0:0]    port_key_11_1_3,
  input      [0:0]    port_key_11_1_4,
  input      [0:0]    port_key_11_1_5,
  input      [0:0]    port_key_11_1_6,
  input      [0:0]    port_key_11_1_7,
  input      [0:0]    port_key_11_2_0,
  input      [0:0]    port_key_11_2_1,
  input      [0:0]    port_key_11_2_2,
  input      [0:0]    port_key_11_2_3,
  input      [0:0]    port_key_11_2_4,
  input      [0:0]    port_key_11_2_5,
  input      [0:0]    port_key_11_2_6,
  input      [0:0]    port_key_11_2_7,
  input      [0:0]    port_key_11_3_0,
  input      [0:0]    port_key_11_3_1,
  input      [0:0]    port_key_11_3_2,
  input      [0:0]    port_key_11_3_3,
  input      [0:0]    port_key_11_3_4,
  input      [0:0]    port_key_11_3_5,
  input      [0:0]    port_key_11_3_6,
  input      [0:0]    port_key_11_3_7,
  input      [0:0]    port_key_12_0_0,
  input      [0:0]    port_key_12_0_1,
  input      [0:0]    port_key_12_0_2,
  input      [0:0]    port_key_12_0_3,
  input      [0:0]    port_key_12_0_4,
  input      [0:0]    port_key_12_0_5,
  input      [0:0]    port_key_12_0_6,
  input      [0:0]    port_key_12_0_7,
  input      [0:0]    port_key_12_1_0,
  input      [0:0]    port_key_12_1_1,
  input      [0:0]    port_key_12_1_2,
  input      [0:0]    port_key_12_1_3,
  input      [0:0]    port_key_12_1_4,
  input      [0:0]    port_key_12_1_5,
  input      [0:0]    port_key_12_1_6,
  input      [0:0]    port_key_12_1_7,
  input      [0:0]    port_key_12_2_0,
  input      [0:0]    port_key_12_2_1,
  input      [0:0]    port_key_12_2_2,
  input      [0:0]    port_key_12_2_3,
  input      [0:0]    port_key_12_2_4,
  input      [0:0]    port_key_12_2_5,
  input      [0:0]    port_key_12_2_6,
  input      [0:0]    port_key_12_2_7,
  input      [0:0]    port_key_12_3_0,
  input      [0:0]    port_key_12_3_1,
  input      [0:0]    port_key_12_3_2,
  input      [0:0]    port_key_12_3_3,
  input      [0:0]    port_key_12_3_4,
  input      [0:0]    port_key_12_3_5,
  input      [0:0]    port_key_12_3_6,
  input      [0:0]    port_key_12_3_7,
  input      [0:0]    port_key_13_0_0,
  input      [0:0]    port_key_13_0_1,
  input      [0:0]    port_key_13_0_2,
  input      [0:0]    port_key_13_0_3,
  input      [0:0]    port_key_13_0_4,
  input      [0:0]    port_key_13_0_5,
  input      [0:0]    port_key_13_0_6,
  input      [0:0]    port_key_13_0_7,
  input      [0:0]    port_key_13_1_0,
  input      [0:0]    port_key_13_1_1,
  input      [0:0]    port_key_13_1_2,
  input      [0:0]    port_key_13_1_3,
  input      [0:0]    port_key_13_1_4,
  input      [0:0]    port_key_13_1_5,
  input      [0:0]    port_key_13_1_6,
  input      [0:0]    port_key_13_1_7,
  input      [0:0]    port_key_13_2_0,
  input      [0:0]    port_key_13_2_1,
  input      [0:0]    port_key_13_2_2,
  input      [0:0]    port_key_13_2_3,
  input      [0:0]    port_key_13_2_4,
  input      [0:0]    port_key_13_2_5,
  input      [0:0]    port_key_13_2_6,
  input      [0:0]    port_key_13_2_7,
  input      [0:0]    port_key_13_3_0,
  input      [0:0]    port_key_13_3_1,
  input      [0:0]    port_key_13_3_2,
  input      [0:0]    port_key_13_3_3,
  input      [0:0]    port_key_13_3_4,
  input      [0:0]    port_key_13_3_5,
  input      [0:0]    port_key_13_3_6,
  input      [0:0]    port_key_13_3_7,
  input      [0:0]    port_key_14_0_0,
  input      [0:0]    port_key_14_0_1,
  input      [0:0]    port_key_14_0_2,
  input      [0:0]    port_key_14_0_3,
  input      [0:0]    port_key_14_0_4,
  input      [0:0]    port_key_14_0_5,
  input      [0:0]    port_key_14_0_6,
  input      [0:0]    port_key_14_0_7,
  input      [0:0]    port_key_14_1_0,
  input      [0:0]    port_key_14_1_1,
  input      [0:0]    port_key_14_1_2,
  input      [0:0]    port_key_14_1_3,
  input      [0:0]    port_key_14_1_4,
  input      [0:0]    port_key_14_1_5,
  input      [0:0]    port_key_14_1_6,
  input      [0:0]    port_key_14_1_7,
  input      [0:0]    port_key_14_2_0,
  input      [0:0]    port_key_14_2_1,
  input      [0:0]    port_key_14_2_2,
  input      [0:0]    port_key_14_2_3,
  input      [0:0]    port_key_14_2_4,
  input      [0:0]    port_key_14_2_5,
  input      [0:0]    port_key_14_2_6,
  input      [0:0]    port_key_14_2_7,
  input      [0:0]    port_key_14_3_0,
  input      [0:0]    port_key_14_3_1,
  input      [0:0]    port_key_14_3_2,
  input      [0:0]    port_key_14_3_3,
  input      [0:0]    port_key_14_3_4,
  input      [0:0]    port_key_14_3_5,
  input      [0:0]    port_key_14_3_6,
  input      [0:0]    port_key_14_3_7,
  input      [0:0]    port_key_15_0_0,
  input      [0:0]    port_key_15_0_1,
  input      [0:0]    port_key_15_0_2,
  input      [0:0]    port_key_15_0_3,
  input      [0:0]    port_key_15_0_4,
  input      [0:0]    port_key_15_0_5,
  input      [0:0]    port_key_15_0_6,
  input      [0:0]    port_key_15_0_7,
  input      [0:0]    port_key_15_1_0,
  input      [0:0]    port_key_15_1_1,
  input      [0:0]    port_key_15_1_2,
  input      [0:0]    port_key_15_1_3,
  input      [0:0]    port_key_15_1_4,
  input      [0:0]    port_key_15_1_5,
  input      [0:0]    port_key_15_1_6,
  input      [0:0]    port_key_15_1_7,
  input      [0:0]    port_key_15_2_0,
  input      [0:0]    port_key_15_2_1,
  input      [0:0]    port_key_15_2_2,
  input      [0:0]    port_key_15_2_3,
  input      [0:0]    port_key_15_2_4,
  input      [0:0]    port_key_15_2_5,
  input      [0:0]    port_key_15_2_6,
  input      [0:0]    port_key_15_2_7,
  input      [0:0]    port_key_15_3_0,
  input      [0:0]    port_key_15_3_1,
  input      [0:0]    port_key_15_3_2,
  input      [0:0]    port_key_15_3_3,
  input      [0:0]    port_key_15_3_4,
  input      [0:0]    port_key_15_3_5,
  input      [0:0]    port_key_15_3_6,
  input      [0:0]    port_key_15_3_7,
  output     [0:0]    port_state_out_0_0_0,
  output     [0:0]    port_state_out_0_0_1,
  output     [0:0]    port_state_out_0_0_2,
  output     [0:0]    port_state_out_0_0_3,
  output     [0:0]    port_state_out_0_0_4,
  output     [0:0]    port_state_out_0_0_5,
  output     [0:0]    port_state_out_0_0_6,
  output     [0:0]    port_state_out_0_0_7,
  output     [0:0]    port_state_out_0_1_0,
  output     [0:0]    port_state_out_0_1_1,
  output     [0:0]    port_state_out_0_1_2,
  output     [0:0]    port_state_out_0_1_3,
  output     [0:0]    port_state_out_0_1_4,
  output     [0:0]    port_state_out_0_1_5,
  output     [0:0]    port_state_out_0_1_6,
  output     [0:0]    port_state_out_0_1_7,
  output     [0:0]    port_state_out_0_2_0,
  output     [0:0]    port_state_out_0_2_1,
  output     [0:0]    port_state_out_0_2_2,
  output     [0:0]    port_state_out_0_2_3,
  output     [0:0]    port_state_out_0_2_4,
  output     [0:0]    port_state_out_0_2_5,
  output     [0:0]    port_state_out_0_2_6,
  output     [0:0]    port_state_out_0_2_7,
  output     [0:0]    port_state_out_0_3_0,
  output     [0:0]    port_state_out_0_3_1,
  output     [0:0]    port_state_out_0_3_2,
  output     [0:0]    port_state_out_0_3_3,
  output     [0:0]    port_state_out_0_3_4,
  output     [0:0]    port_state_out_0_3_5,
  output     [0:0]    port_state_out_0_3_6,
  output     [0:0]    port_state_out_0_3_7,
  output     [0:0]    port_state_out_1_0_0,
  output     [0:0]    port_state_out_1_0_1,
  output     [0:0]    port_state_out_1_0_2,
  output     [0:0]    port_state_out_1_0_3,
  output     [0:0]    port_state_out_1_0_4,
  output     [0:0]    port_state_out_1_0_5,
  output     [0:0]    port_state_out_1_0_6,
  output     [0:0]    port_state_out_1_0_7,
  output     [0:0]    port_state_out_1_1_0,
  output     [0:0]    port_state_out_1_1_1,
  output     [0:0]    port_state_out_1_1_2,
  output     [0:0]    port_state_out_1_1_3,
  output     [0:0]    port_state_out_1_1_4,
  output     [0:0]    port_state_out_1_1_5,
  output     [0:0]    port_state_out_1_1_6,
  output     [0:0]    port_state_out_1_1_7,
  output     [0:0]    port_state_out_1_2_0,
  output     [0:0]    port_state_out_1_2_1,
  output     [0:0]    port_state_out_1_2_2,
  output     [0:0]    port_state_out_1_2_3,
  output     [0:0]    port_state_out_1_2_4,
  output     [0:0]    port_state_out_1_2_5,
  output     [0:0]    port_state_out_1_2_6,
  output     [0:0]    port_state_out_1_2_7,
  output     [0:0]    port_state_out_1_3_0,
  output     [0:0]    port_state_out_1_3_1,
  output     [0:0]    port_state_out_1_3_2,
  output     [0:0]    port_state_out_1_3_3,
  output     [0:0]    port_state_out_1_3_4,
  output     [0:0]    port_state_out_1_3_5,
  output     [0:0]    port_state_out_1_3_6,
  output     [0:0]    port_state_out_1_3_7,
  output     [0:0]    port_state_out_2_0_0,
  output     [0:0]    port_state_out_2_0_1,
  output     [0:0]    port_state_out_2_0_2,
  output     [0:0]    port_state_out_2_0_3,
  output     [0:0]    port_state_out_2_0_4,
  output     [0:0]    port_state_out_2_0_5,
  output     [0:0]    port_state_out_2_0_6,
  output     [0:0]    port_state_out_2_0_7,
  output     [0:0]    port_state_out_2_1_0,
  output     [0:0]    port_state_out_2_1_1,
  output     [0:0]    port_state_out_2_1_2,
  output     [0:0]    port_state_out_2_1_3,
  output     [0:0]    port_state_out_2_1_4,
  output     [0:0]    port_state_out_2_1_5,
  output     [0:0]    port_state_out_2_1_6,
  output     [0:0]    port_state_out_2_1_7,
  output     [0:0]    port_state_out_2_2_0,
  output     [0:0]    port_state_out_2_2_1,
  output     [0:0]    port_state_out_2_2_2,
  output     [0:0]    port_state_out_2_2_3,
  output     [0:0]    port_state_out_2_2_4,
  output     [0:0]    port_state_out_2_2_5,
  output     [0:0]    port_state_out_2_2_6,
  output     [0:0]    port_state_out_2_2_7,
  output     [0:0]    port_state_out_2_3_0,
  output     [0:0]    port_state_out_2_3_1,
  output     [0:0]    port_state_out_2_3_2,
  output     [0:0]    port_state_out_2_3_3,
  output     [0:0]    port_state_out_2_3_4,
  output     [0:0]    port_state_out_2_3_5,
  output     [0:0]    port_state_out_2_3_6,
  output     [0:0]    port_state_out_2_3_7,
  output     [0:0]    port_state_out_3_0_0,
  output     [0:0]    port_state_out_3_0_1,
  output     [0:0]    port_state_out_3_0_2,
  output     [0:0]    port_state_out_3_0_3,
  output     [0:0]    port_state_out_3_0_4,
  output     [0:0]    port_state_out_3_0_5,
  output     [0:0]    port_state_out_3_0_6,
  output     [0:0]    port_state_out_3_0_7,
  output     [0:0]    port_state_out_3_1_0,
  output     [0:0]    port_state_out_3_1_1,
  output     [0:0]    port_state_out_3_1_2,
  output     [0:0]    port_state_out_3_1_3,
  output     [0:0]    port_state_out_3_1_4,
  output     [0:0]    port_state_out_3_1_5,
  output     [0:0]    port_state_out_3_1_6,
  output     [0:0]    port_state_out_3_1_7,
  output     [0:0]    port_state_out_3_2_0,
  output     [0:0]    port_state_out_3_2_1,
  output     [0:0]    port_state_out_3_2_2,
  output     [0:0]    port_state_out_3_2_3,
  output     [0:0]    port_state_out_3_2_4,
  output     [0:0]    port_state_out_3_2_5,
  output     [0:0]    port_state_out_3_2_6,
  output     [0:0]    port_state_out_3_2_7,
  output     [0:0]    port_state_out_3_3_0,
  output     [0:0]    port_state_out_3_3_1,
  output     [0:0]    port_state_out_3_3_2,
  output     [0:0]    port_state_out_3_3_3,
  output     [0:0]    port_state_out_3_3_4,
  output     [0:0]    port_state_out_3_3_5,
  output     [0:0]    port_state_out_3_3_6,
  output     [0:0]    port_state_out_3_3_7,
  output     [0:0]    port_state_out_4_0_0,
  output     [0:0]    port_state_out_4_0_1,
  output     [0:0]    port_state_out_4_0_2,
  output     [0:0]    port_state_out_4_0_3,
  output     [0:0]    port_state_out_4_0_4,
  output     [0:0]    port_state_out_4_0_5,
  output     [0:0]    port_state_out_4_0_6,
  output     [0:0]    port_state_out_4_0_7,
  output     [0:0]    port_state_out_4_1_0,
  output     [0:0]    port_state_out_4_1_1,
  output     [0:0]    port_state_out_4_1_2,
  output     [0:0]    port_state_out_4_1_3,
  output     [0:0]    port_state_out_4_1_4,
  output     [0:0]    port_state_out_4_1_5,
  output     [0:0]    port_state_out_4_1_6,
  output     [0:0]    port_state_out_4_1_7,
  output     [0:0]    port_state_out_4_2_0,
  output     [0:0]    port_state_out_4_2_1,
  output     [0:0]    port_state_out_4_2_2,
  output     [0:0]    port_state_out_4_2_3,
  output     [0:0]    port_state_out_4_2_4,
  output     [0:0]    port_state_out_4_2_5,
  output     [0:0]    port_state_out_4_2_6,
  output     [0:0]    port_state_out_4_2_7,
  output     [0:0]    port_state_out_4_3_0,
  output     [0:0]    port_state_out_4_3_1,
  output     [0:0]    port_state_out_4_3_2,
  output     [0:0]    port_state_out_4_3_3,
  output     [0:0]    port_state_out_4_3_4,
  output     [0:0]    port_state_out_4_3_5,
  output     [0:0]    port_state_out_4_3_6,
  output     [0:0]    port_state_out_4_3_7,
  output     [0:0]    port_state_out_5_0_0,
  output     [0:0]    port_state_out_5_0_1,
  output     [0:0]    port_state_out_5_0_2,
  output     [0:0]    port_state_out_5_0_3,
  output     [0:0]    port_state_out_5_0_4,
  output     [0:0]    port_state_out_5_0_5,
  output     [0:0]    port_state_out_5_0_6,
  output     [0:0]    port_state_out_5_0_7,
  output     [0:0]    port_state_out_5_1_0,
  output     [0:0]    port_state_out_5_1_1,
  output     [0:0]    port_state_out_5_1_2,
  output     [0:0]    port_state_out_5_1_3,
  output     [0:0]    port_state_out_5_1_4,
  output     [0:0]    port_state_out_5_1_5,
  output     [0:0]    port_state_out_5_1_6,
  output     [0:0]    port_state_out_5_1_7,
  output     [0:0]    port_state_out_5_2_0,
  output     [0:0]    port_state_out_5_2_1,
  output     [0:0]    port_state_out_5_2_2,
  output     [0:0]    port_state_out_5_2_3,
  output     [0:0]    port_state_out_5_2_4,
  output     [0:0]    port_state_out_5_2_5,
  output     [0:0]    port_state_out_5_2_6,
  output     [0:0]    port_state_out_5_2_7,
  output     [0:0]    port_state_out_5_3_0,
  output     [0:0]    port_state_out_5_3_1,
  output     [0:0]    port_state_out_5_3_2,
  output     [0:0]    port_state_out_5_3_3,
  output     [0:0]    port_state_out_5_3_4,
  output     [0:0]    port_state_out_5_3_5,
  output     [0:0]    port_state_out_5_3_6,
  output     [0:0]    port_state_out_5_3_7,
  output     [0:0]    port_state_out_6_0_0,
  output     [0:0]    port_state_out_6_0_1,
  output     [0:0]    port_state_out_6_0_2,
  output     [0:0]    port_state_out_6_0_3,
  output     [0:0]    port_state_out_6_0_4,
  output     [0:0]    port_state_out_6_0_5,
  output     [0:0]    port_state_out_6_0_6,
  output     [0:0]    port_state_out_6_0_7,
  output     [0:0]    port_state_out_6_1_0,
  output     [0:0]    port_state_out_6_1_1,
  output     [0:0]    port_state_out_6_1_2,
  output     [0:0]    port_state_out_6_1_3,
  output     [0:0]    port_state_out_6_1_4,
  output     [0:0]    port_state_out_6_1_5,
  output     [0:0]    port_state_out_6_1_6,
  output     [0:0]    port_state_out_6_1_7,
  output     [0:0]    port_state_out_6_2_0,
  output     [0:0]    port_state_out_6_2_1,
  output     [0:0]    port_state_out_6_2_2,
  output     [0:0]    port_state_out_6_2_3,
  output     [0:0]    port_state_out_6_2_4,
  output     [0:0]    port_state_out_6_2_5,
  output     [0:0]    port_state_out_6_2_6,
  output     [0:0]    port_state_out_6_2_7,
  output     [0:0]    port_state_out_6_3_0,
  output     [0:0]    port_state_out_6_3_1,
  output     [0:0]    port_state_out_6_3_2,
  output     [0:0]    port_state_out_6_3_3,
  output     [0:0]    port_state_out_6_3_4,
  output     [0:0]    port_state_out_6_3_5,
  output     [0:0]    port_state_out_6_3_6,
  output     [0:0]    port_state_out_6_3_7,
  output     [0:0]    port_state_out_7_0_0,
  output     [0:0]    port_state_out_7_0_1,
  output     [0:0]    port_state_out_7_0_2,
  output     [0:0]    port_state_out_7_0_3,
  output     [0:0]    port_state_out_7_0_4,
  output     [0:0]    port_state_out_7_0_5,
  output     [0:0]    port_state_out_7_0_6,
  output     [0:0]    port_state_out_7_0_7,
  output     [0:0]    port_state_out_7_1_0,
  output     [0:0]    port_state_out_7_1_1,
  output     [0:0]    port_state_out_7_1_2,
  output     [0:0]    port_state_out_7_1_3,
  output     [0:0]    port_state_out_7_1_4,
  output     [0:0]    port_state_out_7_1_5,
  output     [0:0]    port_state_out_7_1_6,
  output     [0:0]    port_state_out_7_1_7,
  output     [0:0]    port_state_out_7_2_0,
  output     [0:0]    port_state_out_7_2_1,
  output     [0:0]    port_state_out_7_2_2,
  output     [0:0]    port_state_out_7_2_3,
  output     [0:0]    port_state_out_7_2_4,
  output     [0:0]    port_state_out_7_2_5,
  output     [0:0]    port_state_out_7_2_6,
  output     [0:0]    port_state_out_7_2_7,
  output     [0:0]    port_state_out_7_3_0,
  output     [0:0]    port_state_out_7_3_1,
  output     [0:0]    port_state_out_7_3_2,
  output     [0:0]    port_state_out_7_3_3,
  output     [0:0]    port_state_out_7_3_4,
  output     [0:0]    port_state_out_7_3_5,
  output     [0:0]    port_state_out_7_3_6,
  output     [0:0]    port_state_out_7_3_7,
  output     [0:0]    port_state_out_8_0_0,
  output     [0:0]    port_state_out_8_0_1,
  output     [0:0]    port_state_out_8_0_2,
  output     [0:0]    port_state_out_8_0_3,
  output     [0:0]    port_state_out_8_0_4,
  output     [0:0]    port_state_out_8_0_5,
  output     [0:0]    port_state_out_8_0_6,
  output     [0:0]    port_state_out_8_0_7,
  output     [0:0]    port_state_out_8_1_0,
  output     [0:0]    port_state_out_8_1_1,
  output     [0:0]    port_state_out_8_1_2,
  output     [0:0]    port_state_out_8_1_3,
  output     [0:0]    port_state_out_8_1_4,
  output     [0:0]    port_state_out_8_1_5,
  output     [0:0]    port_state_out_8_1_6,
  output     [0:0]    port_state_out_8_1_7,
  output     [0:0]    port_state_out_8_2_0,
  output     [0:0]    port_state_out_8_2_1,
  output     [0:0]    port_state_out_8_2_2,
  output     [0:0]    port_state_out_8_2_3,
  output     [0:0]    port_state_out_8_2_4,
  output     [0:0]    port_state_out_8_2_5,
  output     [0:0]    port_state_out_8_2_6,
  output     [0:0]    port_state_out_8_2_7,
  output     [0:0]    port_state_out_8_3_0,
  output     [0:0]    port_state_out_8_3_1,
  output     [0:0]    port_state_out_8_3_2,
  output     [0:0]    port_state_out_8_3_3,
  output     [0:0]    port_state_out_8_3_4,
  output     [0:0]    port_state_out_8_3_5,
  output     [0:0]    port_state_out_8_3_6,
  output     [0:0]    port_state_out_8_3_7,
  output     [0:0]    port_state_out_9_0_0,
  output     [0:0]    port_state_out_9_0_1,
  output     [0:0]    port_state_out_9_0_2,
  output     [0:0]    port_state_out_9_0_3,
  output     [0:0]    port_state_out_9_0_4,
  output     [0:0]    port_state_out_9_0_5,
  output     [0:0]    port_state_out_9_0_6,
  output     [0:0]    port_state_out_9_0_7,
  output     [0:0]    port_state_out_9_1_0,
  output     [0:0]    port_state_out_9_1_1,
  output     [0:0]    port_state_out_9_1_2,
  output     [0:0]    port_state_out_9_1_3,
  output     [0:0]    port_state_out_9_1_4,
  output     [0:0]    port_state_out_9_1_5,
  output     [0:0]    port_state_out_9_1_6,
  output     [0:0]    port_state_out_9_1_7,
  output     [0:0]    port_state_out_9_2_0,
  output     [0:0]    port_state_out_9_2_1,
  output     [0:0]    port_state_out_9_2_2,
  output     [0:0]    port_state_out_9_2_3,
  output     [0:0]    port_state_out_9_2_4,
  output     [0:0]    port_state_out_9_2_5,
  output     [0:0]    port_state_out_9_2_6,
  output     [0:0]    port_state_out_9_2_7,
  output     [0:0]    port_state_out_9_3_0,
  output     [0:0]    port_state_out_9_3_1,
  output     [0:0]    port_state_out_9_3_2,
  output     [0:0]    port_state_out_9_3_3,
  output     [0:0]    port_state_out_9_3_4,
  output     [0:0]    port_state_out_9_3_5,
  output     [0:0]    port_state_out_9_3_6,
  output     [0:0]    port_state_out_9_3_7,
  output     [0:0]    port_state_out_10_0_0,
  output     [0:0]    port_state_out_10_0_1,
  output     [0:0]    port_state_out_10_0_2,
  output     [0:0]    port_state_out_10_0_3,
  output     [0:0]    port_state_out_10_0_4,
  output     [0:0]    port_state_out_10_0_5,
  output     [0:0]    port_state_out_10_0_6,
  output     [0:0]    port_state_out_10_0_7,
  output     [0:0]    port_state_out_10_1_0,
  output     [0:0]    port_state_out_10_1_1,
  output     [0:0]    port_state_out_10_1_2,
  output     [0:0]    port_state_out_10_1_3,
  output     [0:0]    port_state_out_10_1_4,
  output     [0:0]    port_state_out_10_1_5,
  output     [0:0]    port_state_out_10_1_6,
  output     [0:0]    port_state_out_10_1_7,
  output     [0:0]    port_state_out_10_2_0,
  output     [0:0]    port_state_out_10_2_1,
  output     [0:0]    port_state_out_10_2_2,
  output     [0:0]    port_state_out_10_2_3,
  output     [0:0]    port_state_out_10_2_4,
  output     [0:0]    port_state_out_10_2_5,
  output     [0:0]    port_state_out_10_2_6,
  output     [0:0]    port_state_out_10_2_7,
  output     [0:0]    port_state_out_10_3_0,
  output     [0:0]    port_state_out_10_3_1,
  output     [0:0]    port_state_out_10_3_2,
  output     [0:0]    port_state_out_10_3_3,
  output     [0:0]    port_state_out_10_3_4,
  output     [0:0]    port_state_out_10_3_5,
  output     [0:0]    port_state_out_10_3_6,
  output     [0:0]    port_state_out_10_3_7,
  output     [0:0]    port_state_out_11_0_0,
  output     [0:0]    port_state_out_11_0_1,
  output     [0:0]    port_state_out_11_0_2,
  output     [0:0]    port_state_out_11_0_3,
  output     [0:0]    port_state_out_11_0_4,
  output     [0:0]    port_state_out_11_0_5,
  output     [0:0]    port_state_out_11_0_6,
  output     [0:0]    port_state_out_11_0_7,
  output     [0:0]    port_state_out_11_1_0,
  output     [0:0]    port_state_out_11_1_1,
  output     [0:0]    port_state_out_11_1_2,
  output     [0:0]    port_state_out_11_1_3,
  output     [0:0]    port_state_out_11_1_4,
  output     [0:0]    port_state_out_11_1_5,
  output     [0:0]    port_state_out_11_1_6,
  output     [0:0]    port_state_out_11_1_7,
  output     [0:0]    port_state_out_11_2_0,
  output     [0:0]    port_state_out_11_2_1,
  output     [0:0]    port_state_out_11_2_2,
  output     [0:0]    port_state_out_11_2_3,
  output     [0:0]    port_state_out_11_2_4,
  output     [0:0]    port_state_out_11_2_5,
  output     [0:0]    port_state_out_11_2_6,
  output     [0:0]    port_state_out_11_2_7,
  output     [0:0]    port_state_out_11_3_0,
  output     [0:0]    port_state_out_11_3_1,
  output     [0:0]    port_state_out_11_3_2,
  output     [0:0]    port_state_out_11_3_3,
  output     [0:0]    port_state_out_11_3_4,
  output     [0:0]    port_state_out_11_3_5,
  output     [0:0]    port_state_out_11_3_6,
  output     [0:0]    port_state_out_11_3_7,
  output     [0:0]    port_state_out_12_0_0,
  output     [0:0]    port_state_out_12_0_1,
  output     [0:0]    port_state_out_12_0_2,
  output     [0:0]    port_state_out_12_0_3,
  output     [0:0]    port_state_out_12_0_4,
  output     [0:0]    port_state_out_12_0_5,
  output     [0:0]    port_state_out_12_0_6,
  output     [0:0]    port_state_out_12_0_7,
  output     [0:0]    port_state_out_12_1_0,
  output     [0:0]    port_state_out_12_1_1,
  output     [0:0]    port_state_out_12_1_2,
  output     [0:0]    port_state_out_12_1_3,
  output     [0:0]    port_state_out_12_1_4,
  output     [0:0]    port_state_out_12_1_5,
  output     [0:0]    port_state_out_12_1_6,
  output     [0:0]    port_state_out_12_1_7,
  output     [0:0]    port_state_out_12_2_0,
  output     [0:0]    port_state_out_12_2_1,
  output     [0:0]    port_state_out_12_2_2,
  output     [0:0]    port_state_out_12_2_3,
  output     [0:0]    port_state_out_12_2_4,
  output     [0:0]    port_state_out_12_2_5,
  output     [0:0]    port_state_out_12_2_6,
  output     [0:0]    port_state_out_12_2_7,
  output     [0:0]    port_state_out_12_3_0,
  output     [0:0]    port_state_out_12_3_1,
  output     [0:0]    port_state_out_12_3_2,
  output     [0:0]    port_state_out_12_3_3,
  output     [0:0]    port_state_out_12_3_4,
  output     [0:0]    port_state_out_12_3_5,
  output     [0:0]    port_state_out_12_3_6,
  output     [0:0]    port_state_out_12_3_7,
  output     [0:0]    port_state_out_13_0_0,
  output     [0:0]    port_state_out_13_0_1,
  output     [0:0]    port_state_out_13_0_2,
  output     [0:0]    port_state_out_13_0_3,
  output     [0:0]    port_state_out_13_0_4,
  output     [0:0]    port_state_out_13_0_5,
  output     [0:0]    port_state_out_13_0_6,
  output     [0:0]    port_state_out_13_0_7,
  output     [0:0]    port_state_out_13_1_0,
  output     [0:0]    port_state_out_13_1_1,
  output     [0:0]    port_state_out_13_1_2,
  output     [0:0]    port_state_out_13_1_3,
  output     [0:0]    port_state_out_13_1_4,
  output     [0:0]    port_state_out_13_1_5,
  output     [0:0]    port_state_out_13_1_6,
  output     [0:0]    port_state_out_13_1_7,
  output     [0:0]    port_state_out_13_2_0,
  output     [0:0]    port_state_out_13_2_1,
  output     [0:0]    port_state_out_13_2_2,
  output     [0:0]    port_state_out_13_2_3,
  output     [0:0]    port_state_out_13_2_4,
  output     [0:0]    port_state_out_13_2_5,
  output     [0:0]    port_state_out_13_2_6,
  output     [0:0]    port_state_out_13_2_7,
  output     [0:0]    port_state_out_13_3_0,
  output     [0:0]    port_state_out_13_3_1,
  output     [0:0]    port_state_out_13_3_2,
  output     [0:0]    port_state_out_13_3_3,
  output     [0:0]    port_state_out_13_3_4,
  output     [0:0]    port_state_out_13_3_5,
  output     [0:0]    port_state_out_13_3_6,
  output     [0:0]    port_state_out_13_3_7,
  output     [0:0]    port_state_out_14_0_0,
  output     [0:0]    port_state_out_14_0_1,
  output     [0:0]    port_state_out_14_0_2,
  output     [0:0]    port_state_out_14_0_3,
  output     [0:0]    port_state_out_14_0_4,
  output     [0:0]    port_state_out_14_0_5,
  output     [0:0]    port_state_out_14_0_6,
  output     [0:0]    port_state_out_14_0_7,
  output     [0:0]    port_state_out_14_1_0,
  output     [0:0]    port_state_out_14_1_1,
  output     [0:0]    port_state_out_14_1_2,
  output     [0:0]    port_state_out_14_1_3,
  output     [0:0]    port_state_out_14_1_4,
  output     [0:0]    port_state_out_14_1_5,
  output     [0:0]    port_state_out_14_1_6,
  output     [0:0]    port_state_out_14_1_7,
  output     [0:0]    port_state_out_14_2_0,
  output     [0:0]    port_state_out_14_2_1,
  output     [0:0]    port_state_out_14_2_2,
  output     [0:0]    port_state_out_14_2_3,
  output     [0:0]    port_state_out_14_2_4,
  output     [0:0]    port_state_out_14_2_5,
  output     [0:0]    port_state_out_14_2_6,
  output     [0:0]    port_state_out_14_2_7,
  output     [0:0]    port_state_out_14_3_0,
  output     [0:0]    port_state_out_14_3_1,
  output     [0:0]    port_state_out_14_3_2,
  output     [0:0]    port_state_out_14_3_3,
  output     [0:0]    port_state_out_14_3_4,
  output     [0:0]    port_state_out_14_3_5,
  output     [0:0]    port_state_out_14_3_6,
  output     [0:0]    port_state_out_14_3_7,
  output     [0:0]    port_state_out_15_0_0,
  output     [0:0]    port_state_out_15_0_1,
  output     [0:0]    port_state_out_15_0_2,
  output     [0:0]    port_state_out_15_0_3,
  output     [0:0]    port_state_out_15_0_4,
  output     [0:0]    port_state_out_15_0_5,
  output     [0:0]    port_state_out_15_0_6,
  output     [0:0]    port_state_out_15_0_7,
  output     [0:0]    port_state_out_15_1_0,
  output     [0:0]    port_state_out_15_1_1,
  output     [0:0]    port_state_out_15_1_2,
  output     [0:0]    port_state_out_15_1_3,
  output     [0:0]    port_state_out_15_1_4,
  output     [0:0]    port_state_out_15_1_5,
  output     [0:0]    port_state_out_15_1_6,
  output     [0:0]    port_state_out_15_1_7,
  output     [0:0]    port_state_out_15_2_0,
  output     [0:0]    port_state_out_15_2_1,
  output     [0:0]    port_state_out_15_2_2,
  output     [0:0]    port_state_out_15_2_3,
  output     [0:0]    port_state_out_15_2_4,
  output     [0:0]    port_state_out_15_2_5,
  output     [0:0]    port_state_out_15_2_6,
  output     [0:0]    port_state_out_15_2_7,
  output     [0:0]    port_state_out_15_3_0,
  output     [0:0]    port_state_out_15_3_1,
  output     [0:0]    port_state_out_15_3_2,
  output     [0:0]    port_state_out_15_3_3,
  output     [0:0]    port_state_out_15_3_4,
  output     [0:0]    port_state_out_15_3_5,
  output     [0:0]    port_state_out_15_3_6,
  output     [0:0]    port_state_out_15_3_7,
  input               clk,
  input               reset
);

  wire       [0:0]    keyAdd_port_state_out_0_0_0;
  wire       [0:0]    keyAdd_port_state_out_0_0_1;
  wire       [0:0]    keyAdd_port_state_out_0_0_2;
  wire       [0:0]    keyAdd_port_state_out_0_0_3;
  wire       [0:0]    keyAdd_port_state_out_0_0_4;
  wire       [0:0]    keyAdd_port_state_out_0_0_5;
  wire       [0:0]    keyAdd_port_state_out_0_0_6;
  wire       [0:0]    keyAdd_port_state_out_0_0_7;
  wire       [0:0]    keyAdd_port_state_out_0_1_0;
  wire       [0:0]    keyAdd_port_state_out_0_1_1;
  wire       [0:0]    keyAdd_port_state_out_0_1_2;
  wire       [0:0]    keyAdd_port_state_out_0_1_3;
  wire       [0:0]    keyAdd_port_state_out_0_1_4;
  wire       [0:0]    keyAdd_port_state_out_0_1_5;
  wire       [0:0]    keyAdd_port_state_out_0_1_6;
  wire       [0:0]    keyAdd_port_state_out_0_1_7;
  wire       [0:0]    keyAdd_port_state_out_0_2_0;
  wire       [0:0]    keyAdd_port_state_out_0_2_1;
  wire       [0:0]    keyAdd_port_state_out_0_2_2;
  wire       [0:0]    keyAdd_port_state_out_0_2_3;
  wire       [0:0]    keyAdd_port_state_out_0_2_4;
  wire       [0:0]    keyAdd_port_state_out_0_2_5;
  wire       [0:0]    keyAdd_port_state_out_0_2_6;
  wire       [0:0]    keyAdd_port_state_out_0_2_7;
  wire       [0:0]    keyAdd_port_state_out_0_3_0;
  wire       [0:0]    keyAdd_port_state_out_0_3_1;
  wire       [0:0]    keyAdd_port_state_out_0_3_2;
  wire       [0:0]    keyAdd_port_state_out_0_3_3;
  wire       [0:0]    keyAdd_port_state_out_0_3_4;
  wire       [0:0]    keyAdd_port_state_out_0_3_5;
  wire       [0:0]    keyAdd_port_state_out_0_3_6;
  wire       [0:0]    keyAdd_port_state_out_0_3_7;
  wire       [0:0]    keyAdd_port_state_out_1_0_0;
  wire       [0:0]    keyAdd_port_state_out_1_0_1;
  wire       [0:0]    keyAdd_port_state_out_1_0_2;
  wire       [0:0]    keyAdd_port_state_out_1_0_3;
  wire       [0:0]    keyAdd_port_state_out_1_0_4;
  wire       [0:0]    keyAdd_port_state_out_1_0_5;
  wire       [0:0]    keyAdd_port_state_out_1_0_6;
  wire       [0:0]    keyAdd_port_state_out_1_0_7;
  wire       [0:0]    keyAdd_port_state_out_1_1_0;
  wire       [0:0]    keyAdd_port_state_out_1_1_1;
  wire       [0:0]    keyAdd_port_state_out_1_1_2;
  wire       [0:0]    keyAdd_port_state_out_1_1_3;
  wire       [0:0]    keyAdd_port_state_out_1_1_4;
  wire       [0:0]    keyAdd_port_state_out_1_1_5;
  wire       [0:0]    keyAdd_port_state_out_1_1_6;
  wire       [0:0]    keyAdd_port_state_out_1_1_7;
  wire       [0:0]    keyAdd_port_state_out_1_2_0;
  wire       [0:0]    keyAdd_port_state_out_1_2_1;
  wire       [0:0]    keyAdd_port_state_out_1_2_2;
  wire       [0:0]    keyAdd_port_state_out_1_2_3;
  wire       [0:0]    keyAdd_port_state_out_1_2_4;
  wire       [0:0]    keyAdd_port_state_out_1_2_5;
  wire       [0:0]    keyAdd_port_state_out_1_2_6;
  wire       [0:0]    keyAdd_port_state_out_1_2_7;
  wire       [0:0]    keyAdd_port_state_out_1_3_0;
  wire       [0:0]    keyAdd_port_state_out_1_3_1;
  wire       [0:0]    keyAdd_port_state_out_1_3_2;
  wire       [0:0]    keyAdd_port_state_out_1_3_3;
  wire       [0:0]    keyAdd_port_state_out_1_3_4;
  wire       [0:0]    keyAdd_port_state_out_1_3_5;
  wire       [0:0]    keyAdd_port_state_out_1_3_6;
  wire       [0:0]    keyAdd_port_state_out_1_3_7;
  wire       [0:0]    keyAdd_port_state_out_2_0_0;
  wire       [0:0]    keyAdd_port_state_out_2_0_1;
  wire       [0:0]    keyAdd_port_state_out_2_0_2;
  wire       [0:0]    keyAdd_port_state_out_2_0_3;
  wire       [0:0]    keyAdd_port_state_out_2_0_4;
  wire       [0:0]    keyAdd_port_state_out_2_0_5;
  wire       [0:0]    keyAdd_port_state_out_2_0_6;
  wire       [0:0]    keyAdd_port_state_out_2_0_7;
  wire       [0:0]    keyAdd_port_state_out_2_1_0;
  wire       [0:0]    keyAdd_port_state_out_2_1_1;
  wire       [0:0]    keyAdd_port_state_out_2_1_2;
  wire       [0:0]    keyAdd_port_state_out_2_1_3;
  wire       [0:0]    keyAdd_port_state_out_2_1_4;
  wire       [0:0]    keyAdd_port_state_out_2_1_5;
  wire       [0:0]    keyAdd_port_state_out_2_1_6;
  wire       [0:0]    keyAdd_port_state_out_2_1_7;
  wire       [0:0]    keyAdd_port_state_out_2_2_0;
  wire       [0:0]    keyAdd_port_state_out_2_2_1;
  wire       [0:0]    keyAdd_port_state_out_2_2_2;
  wire       [0:0]    keyAdd_port_state_out_2_2_3;
  wire       [0:0]    keyAdd_port_state_out_2_2_4;
  wire       [0:0]    keyAdd_port_state_out_2_2_5;
  wire       [0:0]    keyAdd_port_state_out_2_2_6;
  wire       [0:0]    keyAdd_port_state_out_2_2_7;
  wire       [0:0]    keyAdd_port_state_out_2_3_0;
  wire       [0:0]    keyAdd_port_state_out_2_3_1;
  wire       [0:0]    keyAdd_port_state_out_2_3_2;
  wire       [0:0]    keyAdd_port_state_out_2_3_3;
  wire       [0:0]    keyAdd_port_state_out_2_3_4;
  wire       [0:0]    keyAdd_port_state_out_2_3_5;
  wire       [0:0]    keyAdd_port_state_out_2_3_6;
  wire       [0:0]    keyAdd_port_state_out_2_3_7;
  wire       [0:0]    keyAdd_port_state_out_3_0_0;
  wire       [0:0]    keyAdd_port_state_out_3_0_1;
  wire       [0:0]    keyAdd_port_state_out_3_0_2;
  wire       [0:0]    keyAdd_port_state_out_3_0_3;
  wire       [0:0]    keyAdd_port_state_out_3_0_4;
  wire       [0:0]    keyAdd_port_state_out_3_0_5;
  wire       [0:0]    keyAdd_port_state_out_3_0_6;
  wire       [0:0]    keyAdd_port_state_out_3_0_7;
  wire       [0:0]    keyAdd_port_state_out_3_1_0;
  wire       [0:0]    keyAdd_port_state_out_3_1_1;
  wire       [0:0]    keyAdd_port_state_out_3_1_2;
  wire       [0:0]    keyAdd_port_state_out_3_1_3;
  wire       [0:0]    keyAdd_port_state_out_3_1_4;
  wire       [0:0]    keyAdd_port_state_out_3_1_5;
  wire       [0:0]    keyAdd_port_state_out_3_1_6;
  wire       [0:0]    keyAdd_port_state_out_3_1_7;
  wire       [0:0]    keyAdd_port_state_out_3_2_0;
  wire       [0:0]    keyAdd_port_state_out_3_2_1;
  wire       [0:0]    keyAdd_port_state_out_3_2_2;
  wire       [0:0]    keyAdd_port_state_out_3_2_3;
  wire       [0:0]    keyAdd_port_state_out_3_2_4;
  wire       [0:0]    keyAdd_port_state_out_3_2_5;
  wire       [0:0]    keyAdd_port_state_out_3_2_6;
  wire       [0:0]    keyAdd_port_state_out_3_2_7;
  wire       [0:0]    keyAdd_port_state_out_3_3_0;
  wire       [0:0]    keyAdd_port_state_out_3_3_1;
  wire       [0:0]    keyAdd_port_state_out_3_3_2;
  wire       [0:0]    keyAdd_port_state_out_3_3_3;
  wire       [0:0]    keyAdd_port_state_out_3_3_4;
  wire       [0:0]    keyAdd_port_state_out_3_3_5;
  wire       [0:0]    keyAdd_port_state_out_3_3_6;
  wire       [0:0]    keyAdd_port_state_out_3_3_7;
  wire       [0:0]    keyAdd_port_state_out_4_0_0;
  wire       [0:0]    keyAdd_port_state_out_4_0_1;
  wire       [0:0]    keyAdd_port_state_out_4_0_2;
  wire       [0:0]    keyAdd_port_state_out_4_0_3;
  wire       [0:0]    keyAdd_port_state_out_4_0_4;
  wire       [0:0]    keyAdd_port_state_out_4_0_5;
  wire       [0:0]    keyAdd_port_state_out_4_0_6;
  wire       [0:0]    keyAdd_port_state_out_4_0_7;
  wire       [0:0]    keyAdd_port_state_out_4_1_0;
  wire       [0:0]    keyAdd_port_state_out_4_1_1;
  wire       [0:0]    keyAdd_port_state_out_4_1_2;
  wire       [0:0]    keyAdd_port_state_out_4_1_3;
  wire       [0:0]    keyAdd_port_state_out_4_1_4;
  wire       [0:0]    keyAdd_port_state_out_4_1_5;
  wire       [0:0]    keyAdd_port_state_out_4_1_6;
  wire       [0:0]    keyAdd_port_state_out_4_1_7;
  wire       [0:0]    keyAdd_port_state_out_4_2_0;
  wire       [0:0]    keyAdd_port_state_out_4_2_1;
  wire       [0:0]    keyAdd_port_state_out_4_2_2;
  wire       [0:0]    keyAdd_port_state_out_4_2_3;
  wire       [0:0]    keyAdd_port_state_out_4_2_4;
  wire       [0:0]    keyAdd_port_state_out_4_2_5;
  wire       [0:0]    keyAdd_port_state_out_4_2_6;
  wire       [0:0]    keyAdd_port_state_out_4_2_7;
  wire       [0:0]    keyAdd_port_state_out_4_3_0;
  wire       [0:0]    keyAdd_port_state_out_4_3_1;
  wire       [0:0]    keyAdd_port_state_out_4_3_2;
  wire       [0:0]    keyAdd_port_state_out_4_3_3;
  wire       [0:0]    keyAdd_port_state_out_4_3_4;
  wire       [0:0]    keyAdd_port_state_out_4_3_5;
  wire       [0:0]    keyAdd_port_state_out_4_3_6;
  wire       [0:0]    keyAdd_port_state_out_4_3_7;
  wire       [0:0]    keyAdd_port_state_out_5_0_0;
  wire       [0:0]    keyAdd_port_state_out_5_0_1;
  wire       [0:0]    keyAdd_port_state_out_5_0_2;
  wire       [0:0]    keyAdd_port_state_out_5_0_3;
  wire       [0:0]    keyAdd_port_state_out_5_0_4;
  wire       [0:0]    keyAdd_port_state_out_5_0_5;
  wire       [0:0]    keyAdd_port_state_out_5_0_6;
  wire       [0:0]    keyAdd_port_state_out_5_0_7;
  wire       [0:0]    keyAdd_port_state_out_5_1_0;
  wire       [0:0]    keyAdd_port_state_out_5_1_1;
  wire       [0:0]    keyAdd_port_state_out_5_1_2;
  wire       [0:0]    keyAdd_port_state_out_5_1_3;
  wire       [0:0]    keyAdd_port_state_out_5_1_4;
  wire       [0:0]    keyAdd_port_state_out_5_1_5;
  wire       [0:0]    keyAdd_port_state_out_5_1_6;
  wire       [0:0]    keyAdd_port_state_out_5_1_7;
  wire       [0:0]    keyAdd_port_state_out_5_2_0;
  wire       [0:0]    keyAdd_port_state_out_5_2_1;
  wire       [0:0]    keyAdd_port_state_out_5_2_2;
  wire       [0:0]    keyAdd_port_state_out_5_2_3;
  wire       [0:0]    keyAdd_port_state_out_5_2_4;
  wire       [0:0]    keyAdd_port_state_out_5_2_5;
  wire       [0:0]    keyAdd_port_state_out_5_2_6;
  wire       [0:0]    keyAdd_port_state_out_5_2_7;
  wire       [0:0]    keyAdd_port_state_out_5_3_0;
  wire       [0:0]    keyAdd_port_state_out_5_3_1;
  wire       [0:0]    keyAdd_port_state_out_5_3_2;
  wire       [0:0]    keyAdd_port_state_out_5_3_3;
  wire       [0:0]    keyAdd_port_state_out_5_3_4;
  wire       [0:0]    keyAdd_port_state_out_5_3_5;
  wire       [0:0]    keyAdd_port_state_out_5_3_6;
  wire       [0:0]    keyAdd_port_state_out_5_3_7;
  wire       [0:0]    keyAdd_port_state_out_6_0_0;
  wire       [0:0]    keyAdd_port_state_out_6_0_1;
  wire       [0:0]    keyAdd_port_state_out_6_0_2;
  wire       [0:0]    keyAdd_port_state_out_6_0_3;
  wire       [0:0]    keyAdd_port_state_out_6_0_4;
  wire       [0:0]    keyAdd_port_state_out_6_0_5;
  wire       [0:0]    keyAdd_port_state_out_6_0_6;
  wire       [0:0]    keyAdd_port_state_out_6_0_7;
  wire       [0:0]    keyAdd_port_state_out_6_1_0;
  wire       [0:0]    keyAdd_port_state_out_6_1_1;
  wire       [0:0]    keyAdd_port_state_out_6_1_2;
  wire       [0:0]    keyAdd_port_state_out_6_1_3;
  wire       [0:0]    keyAdd_port_state_out_6_1_4;
  wire       [0:0]    keyAdd_port_state_out_6_1_5;
  wire       [0:0]    keyAdd_port_state_out_6_1_6;
  wire       [0:0]    keyAdd_port_state_out_6_1_7;
  wire       [0:0]    keyAdd_port_state_out_6_2_0;
  wire       [0:0]    keyAdd_port_state_out_6_2_1;
  wire       [0:0]    keyAdd_port_state_out_6_2_2;
  wire       [0:0]    keyAdd_port_state_out_6_2_3;
  wire       [0:0]    keyAdd_port_state_out_6_2_4;
  wire       [0:0]    keyAdd_port_state_out_6_2_5;
  wire       [0:0]    keyAdd_port_state_out_6_2_6;
  wire       [0:0]    keyAdd_port_state_out_6_2_7;
  wire       [0:0]    keyAdd_port_state_out_6_3_0;
  wire       [0:0]    keyAdd_port_state_out_6_3_1;
  wire       [0:0]    keyAdd_port_state_out_6_3_2;
  wire       [0:0]    keyAdd_port_state_out_6_3_3;
  wire       [0:0]    keyAdd_port_state_out_6_3_4;
  wire       [0:0]    keyAdd_port_state_out_6_3_5;
  wire       [0:0]    keyAdd_port_state_out_6_3_6;
  wire       [0:0]    keyAdd_port_state_out_6_3_7;
  wire       [0:0]    keyAdd_port_state_out_7_0_0;
  wire       [0:0]    keyAdd_port_state_out_7_0_1;
  wire       [0:0]    keyAdd_port_state_out_7_0_2;
  wire       [0:0]    keyAdd_port_state_out_7_0_3;
  wire       [0:0]    keyAdd_port_state_out_7_0_4;
  wire       [0:0]    keyAdd_port_state_out_7_0_5;
  wire       [0:0]    keyAdd_port_state_out_7_0_6;
  wire       [0:0]    keyAdd_port_state_out_7_0_7;
  wire       [0:0]    keyAdd_port_state_out_7_1_0;
  wire       [0:0]    keyAdd_port_state_out_7_1_1;
  wire       [0:0]    keyAdd_port_state_out_7_1_2;
  wire       [0:0]    keyAdd_port_state_out_7_1_3;
  wire       [0:0]    keyAdd_port_state_out_7_1_4;
  wire       [0:0]    keyAdd_port_state_out_7_1_5;
  wire       [0:0]    keyAdd_port_state_out_7_1_6;
  wire       [0:0]    keyAdd_port_state_out_7_1_7;
  wire       [0:0]    keyAdd_port_state_out_7_2_0;
  wire       [0:0]    keyAdd_port_state_out_7_2_1;
  wire       [0:0]    keyAdd_port_state_out_7_2_2;
  wire       [0:0]    keyAdd_port_state_out_7_2_3;
  wire       [0:0]    keyAdd_port_state_out_7_2_4;
  wire       [0:0]    keyAdd_port_state_out_7_2_5;
  wire       [0:0]    keyAdd_port_state_out_7_2_6;
  wire       [0:0]    keyAdd_port_state_out_7_2_7;
  wire       [0:0]    keyAdd_port_state_out_7_3_0;
  wire       [0:0]    keyAdd_port_state_out_7_3_1;
  wire       [0:0]    keyAdd_port_state_out_7_3_2;
  wire       [0:0]    keyAdd_port_state_out_7_3_3;
  wire       [0:0]    keyAdd_port_state_out_7_3_4;
  wire       [0:0]    keyAdd_port_state_out_7_3_5;
  wire       [0:0]    keyAdd_port_state_out_7_3_6;
  wire       [0:0]    keyAdd_port_state_out_7_3_7;
  wire       [0:0]    keyAdd_port_state_out_8_0_0;
  wire       [0:0]    keyAdd_port_state_out_8_0_1;
  wire       [0:0]    keyAdd_port_state_out_8_0_2;
  wire       [0:0]    keyAdd_port_state_out_8_0_3;
  wire       [0:0]    keyAdd_port_state_out_8_0_4;
  wire       [0:0]    keyAdd_port_state_out_8_0_5;
  wire       [0:0]    keyAdd_port_state_out_8_0_6;
  wire       [0:0]    keyAdd_port_state_out_8_0_7;
  wire       [0:0]    keyAdd_port_state_out_8_1_0;
  wire       [0:0]    keyAdd_port_state_out_8_1_1;
  wire       [0:0]    keyAdd_port_state_out_8_1_2;
  wire       [0:0]    keyAdd_port_state_out_8_1_3;
  wire       [0:0]    keyAdd_port_state_out_8_1_4;
  wire       [0:0]    keyAdd_port_state_out_8_1_5;
  wire       [0:0]    keyAdd_port_state_out_8_1_6;
  wire       [0:0]    keyAdd_port_state_out_8_1_7;
  wire       [0:0]    keyAdd_port_state_out_8_2_0;
  wire       [0:0]    keyAdd_port_state_out_8_2_1;
  wire       [0:0]    keyAdd_port_state_out_8_2_2;
  wire       [0:0]    keyAdd_port_state_out_8_2_3;
  wire       [0:0]    keyAdd_port_state_out_8_2_4;
  wire       [0:0]    keyAdd_port_state_out_8_2_5;
  wire       [0:0]    keyAdd_port_state_out_8_2_6;
  wire       [0:0]    keyAdd_port_state_out_8_2_7;
  wire       [0:0]    keyAdd_port_state_out_8_3_0;
  wire       [0:0]    keyAdd_port_state_out_8_3_1;
  wire       [0:0]    keyAdd_port_state_out_8_3_2;
  wire       [0:0]    keyAdd_port_state_out_8_3_3;
  wire       [0:0]    keyAdd_port_state_out_8_3_4;
  wire       [0:0]    keyAdd_port_state_out_8_3_5;
  wire       [0:0]    keyAdd_port_state_out_8_3_6;
  wire       [0:0]    keyAdd_port_state_out_8_3_7;
  wire       [0:0]    keyAdd_port_state_out_9_0_0;
  wire       [0:0]    keyAdd_port_state_out_9_0_1;
  wire       [0:0]    keyAdd_port_state_out_9_0_2;
  wire       [0:0]    keyAdd_port_state_out_9_0_3;
  wire       [0:0]    keyAdd_port_state_out_9_0_4;
  wire       [0:0]    keyAdd_port_state_out_9_0_5;
  wire       [0:0]    keyAdd_port_state_out_9_0_6;
  wire       [0:0]    keyAdd_port_state_out_9_0_7;
  wire       [0:0]    keyAdd_port_state_out_9_1_0;
  wire       [0:0]    keyAdd_port_state_out_9_1_1;
  wire       [0:0]    keyAdd_port_state_out_9_1_2;
  wire       [0:0]    keyAdd_port_state_out_9_1_3;
  wire       [0:0]    keyAdd_port_state_out_9_1_4;
  wire       [0:0]    keyAdd_port_state_out_9_1_5;
  wire       [0:0]    keyAdd_port_state_out_9_1_6;
  wire       [0:0]    keyAdd_port_state_out_9_1_7;
  wire       [0:0]    keyAdd_port_state_out_9_2_0;
  wire       [0:0]    keyAdd_port_state_out_9_2_1;
  wire       [0:0]    keyAdd_port_state_out_9_2_2;
  wire       [0:0]    keyAdd_port_state_out_9_2_3;
  wire       [0:0]    keyAdd_port_state_out_9_2_4;
  wire       [0:0]    keyAdd_port_state_out_9_2_5;
  wire       [0:0]    keyAdd_port_state_out_9_2_6;
  wire       [0:0]    keyAdd_port_state_out_9_2_7;
  wire       [0:0]    keyAdd_port_state_out_9_3_0;
  wire       [0:0]    keyAdd_port_state_out_9_3_1;
  wire       [0:0]    keyAdd_port_state_out_9_3_2;
  wire       [0:0]    keyAdd_port_state_out_9_3_3;
  wire       [0:0]    keyAdd_port_state_out_9_3_4;
  wire       [0:0]    keyAdd_port_state_out_9_3_5;
  wire       [0:0]    keyAdd_port_state_out_9_3_6;
  wire       [0:0]    keyAdd_port_state_out_9_3_7;
  wire       [0:0]    keyAdd_port_state_out_10_0_0;
  wire       [0:0]    keyAdd_port_state_out_10_0_1;
  wire       [0:0]    keyAdd_port_state_out_10_0_2;
  wire       [0:0]    keyAdd_port_state_out_10_0_3;
  wire       [0:0]    keyAdd_port_state_out_10_0_4;
  wire       [0:0]    keyAdd_port_state_out_10_0_5;
  wire       [0:0]    keyAdd_port_state_out_10_0_6;
  wire       [0:0]    keyAdd_port_state_out_10_0_7;
  wire       [0:0]    keyAdd_port_state_out_10_1_0;
  wire       [0:0]    keyAdd_port_state_out_10_1_1;
  wire       [0:0]    keyAdd_port_state_out_10_1_2;
  wire       [0:0]    keyAdd_port_state_out_10_1_3;
  wire       [0:0]    keyAdd_port_state_out_10_1_4;
  wire       [0:0]    keyAdd_port_state_out_10_1_5;
  wire       [0:0]    keyAdd_port_state_out_10_1_6;
  wire       [0:0]    keyAdd_port_state_out_10_1_7;
  wire       [0:0]    keyAdd_port_state_out_10_2_0;
  wire       [0:0]    keyAdd_port_state_out_10_2_1;
  wire       [0:0]    keyAdd_port_state_out_10_2_2;
  wire       [0:0]    keyAdd_port_state_out_10_2_3;
  wire       [0:0]    keyAdd_port_state_out_10_2_4;
  wire       [0:0]    keyAdd_port_state_out_10_2_5;
  wire       [0:0]    keyAdd_port_state_out_10_2_6;
  wire       [0:0]    keyAdd_port_state_out_10_2_7;
  wire       [0:0]    keyAdd_port_state_out_10_3_0;
  wire       [0:0]    keyAdd_port_state_out_10_3_1;
  wire       [0:0]    keyAdd_port_state_out_10_3_2;
  wire       [0:0]    keyAdd_port_state_out_10_3_3;
  wire       [0:0]    keyAdd_port_state_out_10_3_4;
  wire       [0:0]    keyAdd_port_state_out_10_3_5;
  wire       [0:0]    keyAdd_port_state_out_10_3_6;
  wire       [0:0]    keyAdd_port_state_out_10_3_7;
  wire       [0:0]    keyAdd_port_state_out_11_0_0;
  wire       [0:0]    keyAdd_port_state_out_11_0_1;
  wire       [0:0]    keyAdd_port_state_out_11_0_2;
  wire       [0:0]    keyAdd_port_state_out_11_0_3;
  wire       [0:0]    keyAdd_port_state_out_11_0_4;
  wire       [0:0]    keyAdd_port_state_out_11_0_5;
  wire       [0:0]    keyAdd_port_state_out_11_0_6;
  wire       [0:0]    keyAdd_port_state_out_11_0_7;
  wire       [0:0]    keyAdd_port_state_out_11_1_0;
  wire       [0:0]    keyAdd_port_state_out_11_1_1;
  wire       [0:0]    keyAdd_port_state_out_11_1_2;
  wire       [0:0]    keyAdd_port_state_out_11_1_3;
  wire       [0:0]    keyAdd_port_state_out_11_1_4;
  wire       [0:0]    keyAdd_port_state_out_11_1_5;
  wire       [0:0]    keyAdd_port_state_out_11_1_6;
  wire       [0:0]    keyAdd_port_state_out_11_1_7;
  wire       [0:0]    keyAdd_port_state_out_11_2_0;
  wire       [0:0]    keyAdd_port_state_out_11_2_1;
  wire       [0:0]    keyAdd_port_state_out_11_2_2;
  wire       [0:0]    keyAdd_port_state_out_11_2_3;
  wire       [0:0]    keyAdd_port_state_out_11_2_4;
  wire       [0:0]    keyAdd_port_state_out_11_2_5;
  wire       [0:0]    keyAdd_port_state_out_11_2_6;
  wire       [0:0]    keyAdd_port_state_out_11_2_7;
  wire       [0:0]    keyAdd_port_state_out_11_3_0;
  wire       [0:0]    keyAdd_port_state_out_11_3_1;
  wire       [0:0]    keyAdd_port_state_out_11_3_2;
  wire       [0:0]    keyAdd_port_state_out_11_3_3;
  wire       [0:0]    keyAdd_port_state_out_11_3_4;
  wire       [0:0]    keyAdd_port_state_out_11_3_5;
  wire       [0:0]    keyAdd_port_state_out_11_3_6;
  wire       [0:0]    keyAdd_port_state_out_11_3_7;
  wire       [0:0]    keyAdd_port_state_out_12_0_0;
  wire       [0:0]    keyAdd_port_state_out_12_0_1;
  wire       [0:0]    keyAdd_port_state_out_12_0_2;
  wire       [0:0]    keyAdd_port_state_out_12_0_3;
  wire       [0:0]    keyAdd_port_state_out_12_0_4;
  wire       [0:0]    keyAdd_port_state_out_12_0_5;
  wire       [0:0]    keyAdd_port_state_out_12_0_6;
  wire       [0:0]    keyAdd_port_state_out_12_0_7;
  wire       [0:0]    keyAdd_port_state_out_12_1_0;
  wire       [0:0]    keyAdd_port_state_out_12_1_1;
  wire       [0:0]    keyAdd_port_state_out_12_1_2;
  wire       [0:0]    keyAdd_port_state_out_12_1_3;
  wire       [0:0]    keyAdd_port_state_out_12_1_4;
  wire       [0:0]    keyAdd_port_state_out_12_1_5;
  wire       [0:0]    keyAdd_port_state_out_12_1_6;
  wire       [0:0]    keyAdd_port_state_out_12_1_7;
  wire       [0:0]    keyAdd_port_state_out_12_2_0;
  wire       [0:0]    keyAdd_port_state_out_12_2_1;
  wire       [0:0]    keyAdd_port_state_out_12_2_2;
  wire       [0:0]    keyAdd_port_state_out_12_2_3;
  wire       [0:0]    keyAdd_port_state_out_12_2_4;
  wire       [0:0]    keyAdd_port_state_out_12_2_5;
  wire       [0:0]    keyAdd_port_state_out_12_2_6;
  wire       [0:0]    keyAdd_port_state_out_12_2_7;
  wire       [0:0]    keyAdd_port_state_out_12_3_0;
  wire       [0:0]    keyAdd_port_state_out_12_3_1;
  wire       [0:0]    keyAdd_port_state_out_12_3_2;
  wire       [0:0]    keyAdd_port_state_out_12_3_3;
  wire       [0:0]    keyAdd_port_state_out_12_3_4;
  wire       [0:0]    keyAdd_port_state_out_12_3_5;
  wire       [0:0]    keyAdd_port_state_out_12_3_6;
  wire       [0:0]    keyAdd_port_state_out_12_3_7;
  wire       [0:0]    keyAdd_port_state_out_13_0_0;
  wire       [0:0]    keyAdd_port_state_out_13_0_1;
  wire       [0:0]    keyAdd_port_state_out_13_0_2;
  wire       [0:0]    keyAdd_port_state_out_13_0_3;
  wire       [0:0]    keyAdd_port_state_out_13_0_4;
  wire       [0:0]    keyAdd_port_state_out_13_0_5;
  wire       [0:0]    keyAdd_port_state_out_13_0_6;
  wire       [0:0]    keyAdd_port_state_out_13_0_7;
  wire       [0:0]    keyAdd_port_state_out_13_1_0;
  wire       [0:0]    keyAdd_port_state_out_13_1_1;
  wire       [0:0]    keyAdd_port_state_out_13_1_2;
  wire       [0:0]    keyAdd_port_state_out_13_1_3;
  wire       [0:0]    keyAdd_port_state_out_13_1_4;
  wire       [0:0]    keyAdd_port_state_out_13_1_5;
  wire       [0:0]    keyAdd_port_state_out_13_1_6;
  wire       [0:0]    keyAdd_port_state_out_13_1_7;
  wire       [0:0]    keyAdd_port_state_out_13_2_0;
  wire       [0:0]    keyAdd_port_state_out_13_2_1;
  wire       [0:0]    keyAdd_port_state_out_13_2_2;
  wire       [0:0]    keyAdd_port_state_out_13_2_3;
  wire       [0:0]    keyAdd_port_state_out_13_2_4;
  wire       [0:0]    keyAdd_port_state_out_13_2_5;
  wire       [0:0]    keyAdd_port_state_out_13_2_6;
  wire       [0:0]    keyAdd_port_state_out_13_2_7;
  wire       [0:0]    keyAdd_port_state_out_13_3_0;
  wire       [0:0]    keyAdd_port_state_out_13_3_1;
  wire       [0:0]    keyAdd_port_state_out_13_3_2;
  wire       [0:0]    keyAdd_port_state_out_13_3_3;
  wire       [0:0]    keyAdd_port_state_out_13_3_4;
  wire       [0:0]    keyAdd_port_state_out_13_3_5;
  wire       [0:0]    keyAdd_port_state_out_13_3_6;
  wire       [0:0]    keyAdd_port_state_out_13_3_7;
  wire       [0:0]    keyAdd_port_state_out_14_0_0;
  wire       [0:0]    keyAdd_port_state_out_14_0_1;
  wire       [0:0]    keyAdd_port_state_out_14_0_2;
  wire       [0:0]    keyAdd_port_state_out_14_0_3;
  wire       [0:0]    keyAdd_port_state_out_14_0_4;
  wire       [0:0]    keyAdd_port_state_out_14_0_5;
  wire       [0:0]    keyAdd_port_state_out_14_0_6;
  wire       [0:0]    keyAdd_port_state_out_14_0_7;
  wire       [0:0]    keyAdd_port_state_out_14_1_0;
  wire       [0:0]    keyAdd_port_state_out_14_1_1;
  wire       [0:0]    keyAdd_port_state_out_14_1_2;
  wire       [0:0]    keyAdd_port_state_out_14_1_3;
  wire       [0:0]    keyAdd_port_state_out_14_1_4;
  wire       [0:0]    keyAdd_port_state_out_14_1_5;
  wire       [0:0]    keyAdd_port_state_out_14_1_6;
  wire       [0:0]    keyAdd_port_state_out_14_1_7;
  wire       [0:0]    keyAdd_port_state_out_14_2_0;
  wire       [0:0]    keyAdd_port_state_out_14_2_1;
  wire       [0:0]    keyAdd_port_state_out_14_2_2;
  wire       [0:0]    keyAdd_port_state_out_14_2_3;
  wire       [0:0]    keyAdd_port_state_out_14_2_4;
  wire       [0:0]    keyAdd_port_state_out_14_2_5;
  wire       [0:0]    keyAdd_port_state_out_14_2_6;
  wire       [0:0]    keyAdd_port_state_out_14_2_7;
  wire       [0:0]    keyAdd_port_state_out_14_3_0;
  wire       [0:0]    keyAdd_port_state_out_14_3_1;
  wire       [0:0]    keyAdd_port_state_out_14_3_2;
  wire       [0:0]    keyAdd_port_state_out_14_3_3;
  wire       [0:0]    keyAdd_port_state_out_14_3_4;
  wire       [0:0]    keyAdd_port_state_out_14_3_5;
  wire       [0:0]    keyAdd_port_state_out_14_3_6;
  wire       [0:0]    keyAdd_port_state_out_14_3_7;
  wire       [0:0]    keyAdd_port_state_out_15_0_0;
  wire       [0:0]    keyAdd_port_state_out_15_0_1;
  wire       [0:0]    keyAdd_port_state_out_15_0_2;
  wire       [0:0]    keyAdd_port_state_out_15_0_3;
  wire       [0:0]    keyAdd_port_state_out_15_0_4;
  wire       [0:0]    keyAdd_port_state_out_15_0_5;
  wire       [0:0]    keyAdd_port_state_out_15_0_6;
  wire       [0:0]    keyAdd_port_state_out_15_0_7;
  wire       [0:0]    keyAdd_port_state_out_15_1_0;
  wire       [0:0]    keyAdd_port_state_out_15_1_1;
  wire       [0:0]    keyAdd_port_state_out_15_1_2;
  wire       [0:0]    keyAdd_port_state_out_15_1_3;
  wire       [0:0]    keyAdd_port_state_out_15_1_4;
  wire       [0:0]    keyAdd_port_state_out_15_1_5;
  wire       [0:0]    keyAdd_port_state_out_15_1_6;
  wire       [0:0]    keyAdd_port_state_out_15_1_7;
  wire       [0:0]    keyAdd_port_state_out_15_2_0;
  wire       [0:0]    keyAdd_port_state_out_15_2_1;
  wire       [0:0]    keyAdd_port_state_out_15_2_2;
  wire       [0:0]    keyAdd_port_state_out_15_2_3;
  wire       [0:0]    keyAdd_port_state_out_15_2_4;
  wire       [0:0]    keyAdd_port_state_out_15_2_5;
  wire       [0:0]    keyAdd_port_state_out_15_2_6;
  wire       [0:0]    keyAdd_port_state_out_15_2_7;
  wire       [0:0]    keyAdd_port_state_out_15_3_0;
  wire       [0:0]    keyAdd_port_state_out_15_3_1;
  wire       [0:0]    keyAdd_port_state_out_15_3_2;
  wire       [0:0]    keyAdd_port_state_out_15_3_3;
  wire       [0:0]    keyAdd_port_state_out_15_3_4;
  wire       [0:0]    keyAdd_port_state_out_15_3_5;
  wire       [0:0]    keyAdd_port_state_out_15_3_6;
  wire       [0:0]    keyAdd_port_state_out_15_3_7;
  wire       [0:0]    sbox_AES_BoyarPeralta_16_port_o_0_0;
  wire       [0:0]    sbox_AES_BoyarPeralta_16_port_o_0_1;
  wire       [0:0]    sbox_AES_BoyarPeralta_16_port_o_0_2;
  wire       [0:0]    sbox_AES_BoyarPeralta_16_port_o_0_3;
  wire       [0:0]    sbox_AES_BoyarPeralta_16_port_o_0_4;
  wire       [0:0]    sbox_AES_BoyarPeralta_16_port_o_0_5;
  wire       [0:0]    sbox_AES_BoyarPeralta_16_port_o_0_6;
  wire       [0:0]    sbox_AES_BoyarPeralta_16_port_o_0_7;
  wire       [0:0]    sbox_AES_BoyarPeralta_16_port_o_1_0;
  wire       [0:0]    sbox_AES_BoyarPeralta_16_port_o_1_1;
  wire       [0:0]    sbox_AES_BoyarPeralta_16_port_o_1_2;
  wire       [0:0]    sbox_AES_BoyarPeralta_16_port_o_1_3;
  wire       [0:0]    sbox_AES_BoyarPeralta_16_port_o_1_4;
  wire       [0:0]    sbox_AES_BoyarPeralta_16_port_o_1_5;
  wire       [0:0]    sbox_AES_BoyarPeralta_16_port_o_1_6;
  wire       [0:0]    sbox_AES_BoyarPeralta_16_port_o_1_7;
  wire       [0:0]    sbox_AES_BoyarPeralta_16_port_o_2_0;
  wire       [0:0]    sbox_AES_BoyarPeralta_16_port_o_2_1;
  wire       [0:0]    sbox_AES_BoyarPeralta_16_port_o_2_2;
  wire       [0:0]    sbox_AES_BoyarPeralta_16_port_o_2_3;
  wire       [0:0]    sbox_AES_BoyarPeralta_16_port_o_2_4;
  wire       [0:0]    sbox_AES_BoyarPeralta_16_port_o_2_5;
  wire       [0:0]    sbox_AES_BoyarPeralta_16_port_o_2_6;
  wire       [0:0]    sbox_AES_BoyarPeralta_16_port_o_2_7;
  wire       [0:0]    sbox_AES_BoyarPeralta_16_port_o_3_0;
  wire       [0:0]    sbox_AES_BoyarPeralta_16_port_o_3_1;
  wire       [0:0]    sbox_AES_BoyarPeralta_16_port_o_3_2;
  wire       [0:0]    sbox_AES_BoyarPeralta_16_port_o_3_3;
  wire       [0:0]    sbox_AES_BoyarPeralta_16_port_o_3_4;
  wire       [0:0]    sbox_AES_BoyarPeralta_16_port_o_3_5;
  wire       [0:0]    sbox_AES_BoyarPeralta_16_port_o_3_6;
  wire       [0:0]    sbox_AES_BoyarPeralta_16_port_o_3_7;
  wire       [0:0]    sbox_AES_BoyarPeralta_17_port_o_0_0;
  wire       [0:0]    sbox_AES_BoyarPeralta_17_port_o_0_1;
  wire       [0:0]    sbox_AES_BoyarPeralta_17_port_o_0_2;
  wire       [0:0]    sbox_AES_BoyarPeralta_17_port_o_0_3;
  wire       [0:0]    sbox_AES_BoyarPeralta_17_port_o_0_4;
  wire       [0:0]    sbox_AES_BoyarPeralta_17_port_o_0_5;
  wire       [0:0]    sbox_AES_BoyarPeralta_17_port_o_0_6;
  wire       [0:0]    sbox_AES_BoyarPeralta_17_port_o_0_7;
  wire       [0:0]    sbox_AES_BoyarPeralta_17_port_o_1_0;
  wire       [0:0]    sbox_AES_BoyarPeralta_17_port_o_1_1;
  wire       [0:0]    sbox_AES_BoyarPeralta_17_port_o_1_2;
  wire       [0:0]    sbox_AES_BoyarPeralta_17_port_o_1_3;
  wire       [0:0]    sbox_AES_BoyarPeralta_17_port_o_1_4;
  wire       [0:0]    sbox_AES_BoyarPeralta_17_port_o_1_5;
  wire       [0:0]    sbox_AES_BoyarPeralta_17_port_o_1_6;
  wire       [0:0]    sbox_AES_BoyarPeralta_17_port_o_1_7;
  wire       [0:0]    sbox_AES_BoyarPeralta_17_port_o_2_0;
  wire       [0:0]    sbox_AES_BoyarPeralta_17_port_o_2_1;
  wire       [0:0]    sbox_AES_BoyarPeralta_17_port_o_2_2;
  wire       [0:0]    sbox_AES_BoyarPeralta_17_port_o_2_3;
  wire       [0:0]    sbox_AES_BoyarPeralta_17_port_o_2_4;
  wire       [0:0]    sbox_AES_BoyarPeralta_17_port_o_2_5;
  wire       [0:0]    sbox_AES_BoyarPeralta_17_port_o_2_6;
  wire       [0:0]    sbox_AES_BoyarPeralta_17_port_o_2_7;
  wire       [0:0]    sbox_AES_BoyarPeralta_17_port_o_3_0;
  wire       [0:0]    sbox_AES_BoyarPeralta_17_port_o_3_1;
  wire       [0:0]    sbox_AES_BoyarPeralta_17_port_o_3_2;
  wire       [0:0]    sbox_AES_BoyarPeralta_17_port_o_3_3;
  wire       [0:0]    sbox_AES_BoyarPeralta_17_port_o_3_4;
  wire       [0:0]    sbox_AES_BoyarPeralta_17_port_o_3_5;
  wire       [0:0]    sbox_AES_BoyarPeralta_17_port_o_3_6;
  wire       [0:0]    sbox_AES_BoyarPeralta_17_port_o_3_7;
  wire       [0:0]    sbox_AES_BoyarPeralta_18_port_o_0_0;
  wire       [0:0]    sbox_AES_BoyarPeralta_18_port_o_0_1;
  wire       [0:0]    sbox_AES_BoyarPeralta_18_port_o_0_2;
  wire       [0:0]    sbox_AES_BoyarPeralta_18_port_o_0_3;
  wire       [0:0]    sbox_AES_BoyarPeralta_18_port_o_0_4;
  wire       [0:0]    sbox_AES_BoyarPeralta_18_port_o_0_5;
  wire       [0:0]    sbox_AES_BoyarPeralta_18_port_o_0_6;
  wire       [0:0]    sbox_AES_BoyarPeralta_18_port_o_0_7;
  wire       [0:0]    sbox_AES_BoyarPeralta_18_port_o_1_0;
  wire       [0:0]    sbox_AES_BoyarPeralta_18_port_o_1_1;
  wire       [0:0]    sbox_AES_BoyarPeralta_18_port_o_1_2;
  wire       [0:0]    sbox_AES_BoyarPeralta_18_port_o_1_3;
  wire       [0:0]    sbox_AES_BoyarPeralta_18_port_o_1_4;
  wire       [0:0]    sbox_AES_BoyarPeralta_18_port_o_1_5;
  wire       [0:0]    sbox_AES_BoyarPeralta_18_port_o_1_6;
  wire       [0:0]    sbox_AES_BoyarPeralta_18_port_o_1_7;
  wire       [0:0]    sbox_AES_BoyarPeralta_18_port_o_2_0;
  wire       [0:0]    sbox_AES_BoyarPeralta_18_port_o_2_1;
  wire       [0:0]    sbox_AES_BoyarPeralta_18_port_o_2_2;
  wire       [0:0]    sbox_AES_BoyarPeralta_18_port_o_2_3;
  wire       [0:0]    sbox_AES_BoyarPeralta_18_port_o_2_4;
  wire       [0:0]    sbox_AES_BoyarPeralta_18_port_o_2_5;
  wire       [0:0]    sbox_AES_BoyarPeralta_18_port_o_2_6;
  wire       [0:0]    sbox_AES_BoyarPeralta_18_port_o_2_7;
  wire       [0:0]    sbox_AES_BoyarPeralta_18_port_o_3_0;
  wire       [0:0]    sbox_AES_BoyarPeralta_18_port_o_3_1;
  wire       [0:0]    sbox_AES_BoyarPeralta_18_port_o_3_2;
  wire       [0:0]    sbox_AES_BoyarPeralta_18_port_o_3_3;
  wire       [0:0]    sbox_AES_BoyarPeralta_18_port_o_3_4;
  wire       [0:0]    sbox_AES_BoyarPeralta_18_port_o_3_5;
  wire       [0:0]    sbox_AES_BoyarPeralta_18_port_o_3_6;
  wire       [0:0]    sbox_AES_BoyarPeralta_18_port_o_3_7;
  wire       [0:0]    sbox_AES_BoyarPeralta_19_port_o_0_0;
  wire       [0:0]    sbox_AES_BoyarPeralta_19_port_o_0_1;
  wire       [0:0]    sbox_AES_BoyarPeralta_19_port_o_0_2;
  wire       [0:0]    sbox_AES_BoyarPeralta_19_port_o_0_3;
  wire       [0:0]    sbox_AES_BoyarPeralta_19_port_o_0_4;
  wire       [0:0]    sbox_AES_BoyarPeralta_19_port_o_0_5;
  wire       [0:0]    sbox_AES_BoyarPeralta_19_port_o_0_6;
  wire       [0:0]    sbox_AES_BoyarPeralta_19_port_o_0_7;
  wire       [0:0]    sbox_AES_BoyarPeralta_19_port_o_1_0;
  wire       [0:0]    sbox_AES_BoyarPeralta_19_port_o_1_1;
  wire       [0:0]    sbox_AES_BoyarPeralta_19_port_o_1_2;
  wire       [0:0]    sbox_AES_BoyarPeralta_19_port_o_1_3;
  wire       [0:0]    sbox_AES_BoyarPeralta_19_port_o_1_4;
  wire       [0:0]    sbox_AES_BoyarPeralta_19_port_o_1_5;
  wire       [0:0]    sbox_AES_BoyarPeralta_19_port_o_1_6;
  wire       [0:0]    sbox_AES_BoyarPeralta_19_port_o_1_7;
  wire       [0:0]    sbox_AES_BoyarPeralta_19_port_o_2_0;
  wire       [0:0]    sbox_AES_BoyarPeralta_19_port_o_2_1;
  wire       [0:0]    sbox_AES_BoyarPeralta_19_port_o_2_2;
  wire       [0:0]    sbox_AES_BoyarPeralta_19_port_o_2_3;
  wire       [0:0]    sbox_AES_BoyarPeralta_19_port_o_2_4;
  wire       [0:0]    sbox_AES_BoyarPeralta_19_port_o_2_5;
  wire       [0:0]    sbox_AES_BoyarPeralta_19_port_o_2_6;
  wire       [0:0]    sbox_AES_BoyarPeralta_19_port_o_2_7;
  wire       [0:0]    sbox_AES_BoyarPeralta_19_port_o_3_0;
  wire       [0:0]    sbox_AES_BoyarPeralta_19_port_o_3_1;
  wire       [0:0]    sbox_AES_BoyarPeralta_19_port_o_3_2;
  wire       [0:0]    sbox_AES_BoyarPeralta_19_port_o_3_3;
  wire       [0:0]    sbox_AES_BoyarPeralta_19_port_o_3_4;
  wire       [0:0]    sbox_AES_BoyarPeralta_19_port_o_3_5;
  wire       [0:0]    sbox_AES_BoyarPeralta_19_port_o_3_6;
  wire       [0:0]    sbox_AES_BoyarPeralta_19_port_o_3_7;
  wire       [0:0]    sbox_AES_BoyarPeralta_20_port_o_0_0;
  wire       [0:0]    sbox_AES_BoyarPeralta_20_port_o_0_1;
  wire       [0:0]    sbox_AES_BoyarPeralta_20_port_o_0_2;
  wire       [0:0]    sbox_AES_BoyarPeralta_20_port_o_0_3;
  wire       [0:0]    sbox_AES_BoyarPeralta_20_port_o_0_4;
  wire       [0:0]    sbox_AES_BoyarPeralta_20_port_o_0_5;
  wire       [0:0]    sbox_AES_BoyarPeralta_20_port_o_0_6;
  wire       [0:0]    sbox_AES_BoyarPeralta_20_port_o_0_7;
  wire       [0:0]    sbox_AES_BoyarPeralta_20_port_o_1_0;
  wire       [0:0]    sbox_AES_BoyarPeralta_20_port_o_1_1;
  wire       [0:0]    sbox_AES_BoyarPeralta_20_port_o_1_2;
  wire       [0:0]    sbox_AES_BoyarPeralta_20_port_o_1_3;
  wire       [0:0]    sbox_AES_BoyarPeralta_20_port_o_1_4;
  wire       [0:0]    sbox_AES_BoyarPeralta_20_port_o_1_5;
  wire       [0:0]    sbox_AES_BoyarPeralta_20_port_o_1_6;
  wire       [0:0]    sbox_AES_BoyarPeralta_20_port_o_1_7;
  wire       [0:0]    sbox_AES_BoyarPeralta_20_port_o_2_0;
  wire       [0:0]    sbox_AES_BoyarPeralta_20_port_o_2_1;
  wire       [0:0]    sbox_AES_BoyarPeralta_20_port_o_2_2;
  wire       [0:0]    sbox_AES_BoyarPeralta_20_port_o_2_3;
  wire       [0:0]    sbox_AES_BoyarPeralta_20_port_o_2_4;
  wire       [0:0]    sbox_AES_BoyarPeralta_20_port_o_2_5;
  wire       [0:0]    sbox_AES_BoyarPeralta_20_port_o_2_6;
  wire       [0:0]    sbox_AES_BoyarPeralta_20_port_o_2_7;
  wire       [0:0]    sbox_AES_BoyarPeralta_20_port_o_3_0;
  wire       [0:0]    sbox_AES_BoyarPeralta_20_port_o_3_1;
  wire       [0:0]    sbox_AES_BoyarPeralta_20_port_o_3_2;
  wire       [0:0]    sbox_AES_BoyarPeralta_20_port_o_3_3;
  wire       [0:0]    sbox_AES_BoyarPeralta_20_port_o_3_4;
  wire       [0:0]    sbox_AES_BoyarPeralta_20_port_o_3_5;
  wire       [0:0]    sbox_AES_BoyarPeralta_20_port_o_3_6;
  wire       [0:0]    sbox_AES_BoyarPeralta_20_port_o_3_7;
  wire       [0:0]    sbox_AES_BoyarPeralta_21_port_o_0_0;
  wire       [0:0]    sbox_AES_BoyarPeralta_21_port_o_0_1;
  wire       [0:0]    sbox_AES_BoyarPeralta_21_port_o_0_2;
  wire       [0:0]    sbox_AES_BoyarPeralta_21_port_o_0_3;
  wire       [0:0]    sbox_AES_BoyarPeralta_21_port_o_0_4;
  wire       [0:0]    sbox_AES_BoyarPeralta_21_port_o_0_5;
  wire       [0:0]    sbox_AES_BoyarPeralta_21_port_o_0_6;
  wire       [0:0]    sbox_AES_BoyarPeralta_21_port_o_0_7;
  wire       [0:0]    sbox_AES_BoyarPeralta_21_port_o_1_0;
  wire       [0:0]    sbox_AES_BoyarPeralta_21_port_o_1_1;
  wire       [0:0]    sbox_AES_BoyarPeralta_21_port_o_1_2;
  wire       [0:0]    sbox_AES_BoyarPeralta_21_port_o_1_3;
  wire       [0:0]    sbox_AES_BoyarPeralta_21_port_o_1_4;
  wire       [0:0]    sbox_AES_BoyarPeralta_21_port_o_1_5;
  wire       [0:0]    sbox_AES_BoyarPeralta_21_port_o_1_6;
  wire       [0:0]    sbox_AES_BoyarPeralta_21_port_o_1_7;
  wire       [0:0]    sbox_AES_BoyarPeralta_21_port_o_2_0;
  wire       [0:0]    sbox_AES_BoyarPeralta_21_port_o_2_1;
  wire       [0:0]    sbox_AES_BoyarPeralta_21_port_o_2_2;
  wire       [0:0]    sbox_AES_BoyarPeralta_21_port_o_2_3;
  wire       [0:0]    sbox_AES_BoyarPeralta_21_port_o_2_4;
  wire       [0:0]    sbox_AES_BoyarPeralta_21_port_o_2_5;
  wire       [0:0]    sbox_AES_BoyarPeralta_21_port_o_2_6;
  wire       [0:0]    sbox_AES_BoyarPeralta_21_port_o_2_7;
  wire       [0:0]    sbox_AES_BoyarPeralta_21_port_o_3_0;
  wire       [0:0]    sbox_AES_BoyarPeralta_21_port_o_3_1;
  wire       [0:0]    sbox_AES_BoyarPeralta_21_port_o_3_2;
  wire       [0:0]    sbox_AES_BoyarPeralta_21_port_o_3_3;
  wire       [0:0]    sbox_AES_BoyarPeralta_21_port_o_3_4;
  wire       [0:0]    sbox_AES_BoyarPeralta_21_port_o_3_5;
  wire       [0:0]    sbox_AES_BoyarPeralta_21_port_o_3_6;
  wire       [0:0]    sbox_AES_BoyarPeralta_21_port_o_3_7;
  wire       [0:0]    sbox_AES_BoyarPeralta_22_port_o_0_0;
  wire       [0:0]    sbox_AES_BoyarPeralta_22_port_o_0_1;
  wire       [0:0]    sbox_AES_BoyarPeralta_22_port_o_0_2;
  wire       [0:0]    sbox_AES_BoyarPeralta_22_port_o_0_3;
  wire       [0:0]    sbox_AES_BoyarPeralta_22_port_o_0_4;
  wire       [0:0]    sbox_AES_BoyarPeralta_22_port_o_0_5;
  wire       [0:0]    sbox_AES_BoyarPeralta_22_port_o_0_6;
  wire       [0:0]    sbox_AES_BoyarPeralta_22_port_o_0_7;
  wire       [0:0]    sbox_AES_BoyarPeralta_22_port_o_1_0;
  wire       [0:0]    sbox_AES_BoyarPeralta_22_port_o_1_1;
  wire       [0:0]    sbox_AES_BoyarPeralta_22_port_o_1_2;
  wire       [0:0]    sbox_AES_BoyarPeralta_22_port_o_1_3;
  wire       [0:0]    sbox_AES_BoyarPeralta_22_port_o_1_4;
  wire       [0:0]    sbox_AES_BoyarPeralta_22_port_o_1_5;
  wire       [0:0]    sbox_AES_BoyarPeralta_22_port_o_1_6;
  wire       [0:0]    sbox_AES_BoyarPeralta_22_port_o_1_7;
  wire       [0:0]    sbox_AES_BoyarPeralta_22_port_o_2_0;
  wire       [0:0]    sbox_AES_BoyarPeralta_22_port_o_2_1;
  wire       [0:0]    sbox_AES_BoyarPeralta_22_port_o_2_2;
  wire       [0:0]    sbox_AES_BoyarPeralta_22_port_o_2_3;
  wire       [0:0]    sbox_AES_BoyarPeralta_22_port_o_2_4;
  wire       [0:0]    sbox_AES_BoyarPeralta_22_port_o_2_5;
  wire       [0:0]    sbox_AES_BoyarPeralta_22_port_o_2_6;
  wire       [0:0]    sbox_AES_BoyarPeralta_22_port_o_2_7;
  wire       [0:0]    sbox_AES_BoyarPeralta_22_port_o_3_0;
  wire       [0:0]    sbox_AES_BoyarPeralta_22_port_o_3_1;
  wire       [0:0]    sbox_AES_BoyarPeralta_22_port_o_3_2;
  wire       [0:0]    sbox_AES_BoyarPeralta_22_port_o_3_3;
  wire       [0:0]    sbox_AES_BoyarPeralta_22_port_o_3_4;
  wire       [0:0]    sbox_AES_BoyarPeralta_22_port_o_3_5;
  wire       [0:0]    sbox_AES_BoyarPeralta_22_port_o_3_6;
  wire       [0:0]    sbox_AES_BoyarPeralta_22_port_o_3_7;
  wire       [0:0]    sbox_AES_BoyarPeralta_23_port_o_0_0;
  wire       [0:0]    sbox_AES_BoyarPeralta_23_port_o_0_1;
  wire       [0:0]    sbox_AES_BoyarPeralta_23_port_o_0_2;
  wire       [0:0]    sbox_AES_BoyarPeralta_23_port_o_0_3;
  wire       [0:0]    sbox_AES_BoyarPeralta_23_port_o_0_4;
  wire       [0:0]    sbox_AES_BoyarPeralta_23_port_o_0_5;
  wire       [0:0]    sbox_AES_BoyarPeralta_23_port_o_0_6;
  wire       [0:0]    sbox_AES_BoyarPeralta_23_port_o_0_7;
  wire       [0:0]    sbox_AES_BoyarPeralta_23_port_o_1_0;
  wire       [0:0]    sbox_AES_BoyarPeralta_23_port_o_1_1;
  wire       [0:0]    sbox_AES_BoyarPeralta_23_port_o_1_2;
  wire       [0:0]    sbox_AES_BoyarPeralta_23_port_o_1_3;
  wire       [0:0]    sbox_AES_BoyarPeralta_23_port_o_1_4;
  wire       [0:0]    sbox_AES_BoyarPeralta_23_port_o_1_5;
  wire       [0:0]    sbox_AES_BoyarPeralta_23_port_o_1_6;
  wire       [0:0]    sbox_AES_BoyarPeralta_23_port_o_1_7;
  wire       [0:0]    sbox_AES_BoyarPeralta_23_port_o_2_0;
  wire       [0:0]    sbox_AES_BoyarPeralta_23_port_o_2_1;
  wire       [0:0]    sbox_AES_BoyarPeralta_23_port_o_2_2;
  wire       [0:0]    sbox_AES_BoyarPeralta_23_port_o_2_3;
  wire       [0:0]    sbox_AES_BoyarPeralta_23_port_o_2_4;
  wire       [0:0]    sbox_AES_BoyarPeralta_23_port_o_2_5;
  wire       [0:0]    sbox_AES_BoyarPeralta_23_port_o_2_6;
  wire       [0:0]    sbox_AES_BoyarPeralta_23_port_o_2_7;
  wire       [0:0]    sbox_AES_BoyarPeralta_23_port_o_3_0;
  wire       [0:0]    sbox_AES_BoyarPeralta_23_port_o_3_1;
  wire       [0:0]    sbox_AES_BoyarPeralta_23_port_o_3_2;
  wire       [0:0]    sbox_AES_BoyarPeralta_23_port_o_3_3;
  wire       [0:0]    sbox_AES_BoyarPeralta_23_port_o_3_4;
  wire       [0:0]    sbox_AES_BoyarPeralta_23_port_o_3_5;
  wire       [0:0]    sbox_AES_BoyarPeralta_23_port_o_3_6;
  wire       [0:0]    sbox_AES_BoyarPeralta_23_port_o_3_7;
  wire       [0:0]    sbox_AES_BoyarPeralta_24_port_o_0_0;
  wire       [0:0]    sbox_AES_BoyarPeralta_24_port_o_0_1;
  wire       [0:0]    sbox_AES_BoyarPeralta_24_port_o_0_2;
  wire       [0:0]    sbox_AES_BoyarPeralta_24_port_o_0_3;
  wire       [0:0]    sbox_AES_BoyarPeralta_24_port_o_0_4;
  wire       [0:0]    sbox_AES_BoyarPeralta_24_port_o_0_5;
  wire       [0:0]    sbox_AES_BoyarPeralta_24_port_o_0_6;
  wire       [0:0]    sbox_AES_BoyarPeralta_24_port_o_0_7;
  wire       [0:0]    sbox_AES_BoyarPeralta_24_port_o_1_0;
  wire       [0:0]    sbox_AES_BoyarPeralta_24_port_o_1_1;
  wire       [0:0]    sbox_AES_BoyarPeralta_24_port_o_1_2;
  wire       [0:0]    sbox_AES_BoyarPeralta_24_port_o_1_3;
  wire       [0:0]    sbox_AES_BoyarPeralta_24_port_o_1_4;
  wire       [0:0]    sbox_AES_BoyarPeralta_24_port_o_1_5;
  wire       [0:0]    sbox_AES_BoyarPeralta_24_port_o_1_6;
  wire       [0:0]    sbox_AES_BoyarPeralta_24_port_o_1_7;
  wire       [0:0]    sbox_AES_BoyarPeralta_24_port_o_2_0;
  wire       [0:0]    sbox_AES_BoyarPeralta_24_port_o_2_1;
  wire       [0:0]    sbox_AES_BoyarPeralta_24_port_o_2_2;
  wire       [0:0]    sbox_AES_BoyarPeralta_24_port_o_2_3;
  wire       [0:0]    sbox_AES_BoyarPeralta_24_port_o_2_4;
  wire       [0:0]    sbox_AES_BoyarPeralta_24_port_o_2_5;
  wire       [0:0]    sbox_AES_BoyarPeralta_24_port_o_2_6;
  wire       [0:0]    sbox_AES_BoyarPeralta_24_port_o_2_7;
  wire       [0:0]    sbox_AES_BoyarPeralta_24_port_o_3_0;
  wire       [0:0]    sbox_AES_BoyarPeralta_24_port_o_3_1;
  wire       [0:0]    sbox_AES_BoyarPeralta_24_port_o_3_2;
  wire       [0:0]    sbox_AES_BoyarPeralta_24_port_o_3_3;
  wire       [0:0]    sbox_AES_BoyarPeralta_24_port_o_3_4;
  wire       [0:0]    sbox_AES_BoyarPeralta_24_port_o_3_5;
  wire       [0:0]    sbox_AES_BoyarPeralta_24_port_o_3_6;
  wire       [0:0]    sbox_AES_BoyarPeralta_24_port_o_3_7;
  wire       [0:0]    sbox_AES_BoyarPeralta_25_port_o_0_0;
  wire       [0:0]    sbox_AES_BoyarPeralta_25_port_o_0_1;
  wire       [0:0]    sbox_AES_BoyarPeralta_25_port_o_0_2;
  wire       [0:0]    sbox_AES_BoyarPeralta_25_port_o_0_3;
  wire       [0:0]    sbox_AES_BoyarPeralta_25_port_o_0_4;
  wire       [0:0]    sbox_AES_BoyarPeralta_25_port_o_0_5;
  wire       [0:0]    sbox_AES_BoyarPeralta_25_port_o_0_6;
  wire       [0:0]    sbox_AES_BoyarPeralta_25_port_o_0_7;
  wire       [0:0]    sbox_AES_BoyarPeralta_25_port_o_1_0;
  wire       [0:0]    sbox_AES_BoyarPeralta_25_port_o_1_1;
  wire       [0:0]    sbox_AES_BoyarPeralta_25_port_o_1_2;
  wire       [0:0]    sbox_AES_BoyarPeralta_25_port_o_1_3;
  wire       [0:0]    sbox_AES_BoyarPeralta_25_port_o_1_4;
  wire       [0:0]    sbox_AES_BoyarPeralta_25_port_o_1_5;
  wire       [0:0]    sbox_AES_BoyarPeralta_25_port_o_1_6;
  wire       [0:0]    sbox_AES_BoyarPeralta_25_port_o_1_7;
  wire       [0:0]    sbox_AES_BoyarPeralta_25_port_o_2_0;
  wire       [0:0]    sbox_AES_BoyarPeralta_25_port_o_2_1;
  wire       [0:0]    sbox_AES_BoyarPeralta_25_port_o_2_2;
  wire       [0:0]    sbox_AES_BoyarPeralta_25_port_o_2_3;
  wire       [0:0]    sbox_AES_BoyarPeralta_25_port_o_2_4;
  wire       [0:0]    sbox_AES_BoyarPeralta_25_port_o_2_5;
  wire       [0:0]    sbox_AES_BoyarPeralta_25_port_o_2_6;
  wire       [0:0]    sbox_AES_BoyarPeralta_25_port_o_2_7;
  wire       [0:0]    sbox_AES_BoyarPeralta_25_port_o_3_0;
  wire       [0:0]    sbox_AES_BoyarPeralta_25_port_o_3_1;
  wire       [0:0]    sbox_AES_BoyarPeralta_25_port_o_3_2;
  wire       [0:0]    sbox_AES_BoyarPeralta_25_port_o_3_3;
  wire       [0:0]    sbox_AES_BoyarPeralta_25_port_o_3_4;
  wire       [0:0]    sbox_AES_BoyarPeralta_25_port_o_3_5;
  wire       [0:0]    sbox_AES_BoyarPeralta_25_port_o_3_6;
  wire       [0:0]    sbox_AES_BoyarPeralta_25_port_o_3_7;
  wire       [0:0]    sbox_AES_BoyarPeralta_26_port_o_0_0;
  wire       [0:0]    sbox_AES_BoyarPeralta_26_port_o_0_1;
  wire       [0:0]    sbox_AES_BoyarPeralta_26_port_o_0_2;
  wire       [0:0]    sbox_AES_BoyarPeralta_26_port_o_0_3;
  wire       [0:0]    sbox_AES_BoyarPeralta_26_port_o_0_4;
  wire       [0:0]    sbox_AES_BoyarPeralta_26_port_o_0_5;
  wire       [0:0]    sbox_AES_BoyarPeralta_26_port_o_0_6;
  wire       [0:0]    sbox_AES_BoyarPeralta_26_port_o_0_7;
  wire       [0:0]    sbox_AES_BoyarPeralta_26_port_o_1_0;
  wire       [0:0]    sbox_AES_BoyarPeralta_26_port_o_1_1;
  wire       [0:0]    sbox_AES_BoyarPeralta_26_port_o_1_2;
  wire       [0:0]    sbox_AES_BoyarPeralta_26_port_o_1_3;
  wire       [0:0]    sbox_AES_BoyarPeralta_26_port_o_1_4;
  wire       [0:0]    sbox_AES_BoyarPeralta_26_port_o_1_5;
  wire       [0:0]    sbox_AES_BoyarPeralta_26_port_o_1_6;
  wire       [0:0]    sbox_AES_BoyarPeralta_26_port_o_1_7;
  wire       [0:0]    sbox_AES_BoyarPeralta_26_port_o_2_0;
  wire       [0:0]    sbox_AES_BoyarPeralta_26_port_o_2_1;
  wire       [0:0]    sbox_AES_BoyarPeralta_26_port_o_2_2;
  wire       [0:0]    sbox_AES_BoyarPeralta_26_port_o_2_3;
  wire       [0:0]    sbox_AES_BoyarPeralta_26_port_o_2_4;
  wire       [0:0]    sbox_AES_BoyarPeralta_26_port_o_2_5;
  wire       [0:0]    sbox_AES_BoyarPeralta_26_port_o_2_6;
  wire       [0:0]    sbox_AES_BoyarPeralta_26_port_o_2_7;
  wire       [0:0]    sbox_AES_BoyarPeralta_26_port_o_3_0;
  wire       [0:0]    sbox_AES_BoyarPeralta_26_port_o_3_1;
  wire       [0:0]    sbox_AES_BoyarPeralta_26_port_o_3_2;
  wire       [0:0]    sbox_AES_BoyarPeralta_26_port_o_3_3;
  wire       [0:0]    sbox_AES_BoyarPeralta_26_port_o_3_4;
  wire       [0:0]    sbox_AES_BoyarPeralta_26_port_o_3_5;
  wire       [0:0]    sbox_AES_BoyarPeralta_26_port_o_3_6;
  wire       [0:0]    sbox_AES_BoyarPeralta_26_port_o_3_7;
  wire       [0:0]    sbox_AES_BoyarPeralta_27_port_o_0_0;
  wire       [0:0]    sbox_AES_BoyarPeralta_27_port_o_0_1;
  wire       [0:0]    sbox_AES_BoyarPeralta_27_port_o_0_2;
  wire       [0:0]    sbox_AES_BoyarPeralta_27_port_o_0_3;
  wire       [0:0]    sbox_AES_BoyarPeralta_27_port_o_0_4;
  wire       [0:0]    sbox_AES_BoyarPeralta_27_port_o_0_5;
  wire       [0:0]    sbox_AES_BoyarPeralta_27_port_o_0_6;
  wire       [0:0]    sbox_AES_BoyarPeralta_27_port_o_0_7;
  wire       [0:0]    sbox_AES_BoyarPeralta_27_port_o_1_0;
  wire       [0:0]    sbox_AES_BoyarPeralta_27_port_o_1_1;
  wire       [0:0]    sbox_AES_BoyarPeralta_27_port_o_1_2;
  wire       [0:0]    sbox_AES_BoyarPeralta_27_port_o_1_3;
  wire       [0:0]    sbox_AES_BoyarPeralta_27_port_o_1_4;
  wire       [0:0]    sbox_AES_BoyarPeralta_27_port_o_1_5;
  wire       [0:0]    sbox_AES_BoyarPeralta_27_port_o_1_6;
  wire       [0:0]    sbox_AES_BoyarPeralta_27_port_o_1_7;
  wire       [0:0]    sbox_AES_BoyarPeralta_27_port_o_2_0;
  wire       [0:0]    sbox_AES_BoyarPeralta_27_port_o_2_1;
  wire       [0:0]    sbox_AES_BoyarPeralta_27_port_o_2_2;
  wire       [0:0]    sbox_AES_BoyarPeralta_27_port_o_2_3;
  wire       [0:0]    sbox_AES_BoyarPeralta_27_port_o_2_4;
  wire       [0:0]    sbox_AES_BoyarPeralta_27_port_o_2_5;
  wire       [0:0]    sbox_AES_BoyarPeralta_27_port_o_2_6;
  wire       [0:0]    sbox_AES_BoyarPeralta_27_port_o_2_7;
  wire       [0:0]    sbox_AES_BoyarPeralta_27_port_o_3_0;
  wire       [0:0]    sbox_AES_BoyarPeralta_27_port_o_3_1;
  wire       [0:0]    sbox_AES_BoyarPeralta_27_port_o_3_2;
  wire       [0:0]    sbox_AES_BoyarPeralta_27_port_o_3_3;
  wire       [0:0]    sbox_AES_BoyarPeralta_27_port_o_3_4;
  wire       [0:0]    sbox_AES_BoyarPeralta_27_port_o_3_5;
  wire       [0:0]    sbox_AES_BoyarPeralta_27_port_o_3_6;
  wire       [0:0]    sbox_AES_BoyarPeralta_27_port_o_3_7;
  wire       [0:0]    sbox_AES_BoyarPeralta_28_port_o_0_0;
  wire       [0:0]    sbox_AES_BoyarPeralta_28_port_o_0_1;
  wire       [0:0]    sbox_AES_BoyarPeralta_28_port_o_0_2;
  wire       [0:0]    sbox_AES_BoyarPeralta_28_port_o_0_3;
  wire       [0:0]    sbox_AES_BoyarPeralta_28_port_o_0_4;
  wire       [0:0]    sbox_AES_BoyarPeralta_28_port_o_0_5;
  wire       [0:0]    sbox_AES_BoyarPeralta_28_port_o_0_6;
  wire       [0:0]    sbox_AES_BoyarPeralta_28_port_o_0_7;
  wire       [0:0]    sbox_AES_BoyarPeralta_28_port_o_1_0;
  wire       [0:0]    sbox_AES_BoyarPeralta_28_port_o_1_1;
  wire       [0:0]    sbox_AES_BoyarPeralta_28_port_o_1_2;
  wire       [0:0]    sbox_AES_BoyarPeralta_28_port_o_1_3;
  wire       [0:0]    sbox_AES_BoyarPeralta_28_port_o_1_4;
  wire       [0:0]    sbox_AES_BoyarPeralta_28_port_o_1_5;
  wire       [0:0]    sbox_AES_BoyarPeralta_28_port_o_1_6;
  wire       [0:0]    sbox_AES_BoyarPeralta_28_port_o_1_7;
  wire       [0:0]    sbox_AES_BoyarPeralta_28_port_o_2_0;
  wire       [0:0]    sbox_AES_BoyarPeralta_28_port_o_2_1;
  wire       [0:0]    sbox_AES_BoyarPeralta_28_port_o_2_2;
  wire       [0:0]    sbox_AES_BoyarPeralta_28_port_o_2_3;
  wire       [0:0]    sbox_AES_BoyarPeralta_28_port_o_2_4;
  wire       [0:0]    sbox_AES_BoyarPeralta_28_port_o_2_5;
  wire       [0:0]    sbox_AES_BoyarPeralta_28_port_o_2_6;
  wire       [0:0]    sbox_AES_BoyarPeralta_28_port_o_2_7;
  wire       [0:0]    sbox_AES_BoyarPeralta_28_port_o_3_0;
  wire       [0:0]    sbox_AES_BoyarPeralta_28_port_o_3_1;
  wire       [0:0]    sbox_AES_BoyarPeralta_28_port_o_3_2;
  wire       [0:0]    sbox_AES_BoyarPeralta_28_port_o_3_3;
  wire       [0:0]    sbox_AES_BoyarPeralta_28_port_o_3_4;
  wire       [0:0]    sbox_AES_BoyarPeralta_28_port_o_3_5;
  wire       [0:0]    sbox_AES_BoyarPeralta_28_port_o_3_6;
  wire       [0:0]    sbox_AES_BoyarPeralta_28_port_o_3_7;
  wire       [0:0]    sbox_AES_BoyarPeralta_29_port_o_0_0;
  wire       [0:0]    sbox_AES_BoyarPeralta_29_port_o_0_1;
  wire       [0:0]    sbox_AES_BoyarPeralta_29_port_o_0_2;
  wire       [0:0]    sbox_AES_BoyarPeralta_29_port_o_0_3;
  wire       [0:0]    sbox_AES_BoyarPeralta_29_port_o_0_4;
  wire       [0:0]    sbox_AES_BoyarPeralta_29_port_o_0_5;
  wire       [0:0]    sbox_AES_BoyarPeralta_29_port_o_0_6;
  wire       [0:0]    sbox_AES_BoyarPeralta_29_port_o_0_7;
  wire       [0:0]    sbox_AES_BoyarPeralta_29_port_o_1_0;
  wire       [0:0]    sbox_AES_BoyarPeralta_29_port_o_1_1;
  wire       [0:0]    sbox_AES_BoyarPeralta_29_port_o_1_2;
  wire       [0:0]    sbox_AES_BoyarPeralta_29_port_o_1_3;
  wire       [0:0]    sbox_AES_BoyarPeralta_29_port_o_1_4;
  wire       [0:0]    sbox_AES_BoyarPeralta_29_port_o_1_5;
  wire       [0:0]    sbox_AES_BoyarPeralta_29_port_o_1_6;
  wire       [0:0]    sbox_AES_BoyarPeralta_29_port_o_1_7;
  wire       [0:0]    sbox_AES_BoyarPeralta_29_port_o_2_0;
  wire       [0:0]    sbox_AES_BoyarPeralta_29_port_o_2_1;
  wire       [0:0]    sbox_AES_BoyarPeralta_29_port_o_2_2;
  wire       [0:0]    sbox_AES_BoyarPeralta_29_port_o_2_3;
  wire       [0:0]    sbox_AES_BoyarPeralta_29_port_o_2_4;
  wire       [0:0]    sbox_AES_BoyarPeralta_29_port_o_2_5;
  wire       [0:0]    sbox_AES_BoyarPeralta_29_port_o_2_6;
  wire       [0:0]    sbox_AES_BoyarPeralta_29_port_o_2_7;
  wire       [0:0]    sbox_AES_BoyarPeralta_29_port_o_3_0;
  wire       [0:0]    sbox_AES_BoyarPeralta_29_port_o_3_1;
  wire       [0:0]    sbox_AES_BoyarPeralta_29_port_o_3_2;
  wire       [0:0]    sbox_AES_BoyarPeralta_29_port_o_3_3;
  wire       [0:0]    sbox_AES_BoyarPeralta_29_port_o_3_4;
  wire       [0:0]    sbox_AES_BoyarPeralta_29_port_o_3_5;
  wire       [0:0]    sbox_AES_BoyarPeralta_29_port_o_3_6;
  wire       [0:0]    sbox_AES_BoyarPeralta_29_port_o_3_7;
  wire       [0:0]    sbox_AES_BoyarPeralta_30_port_o_0_0;
  wire       [0:0]    sbox_AES_BoyarPeralta_30_port_o_0_1;
  wire       [0:0]    sbox_AES_BoyarPeralta_30_port_o_0_2;
  wire       [0:0]    sbox_AES_BoyarPeralta_30_port_o_0_3;
  wire       [0:0]    sbox_AES_BoyarPeralta_30_port_o_0_4;
  wire       [0:0]    sbox_AES_BoyarPeralta_30_port_o_0_5;
  wire       [0:0]    sbox_AES_BoyarPeralta_30_port_o_0_6;
  wire       [0:0]    sbox_AES_BoyarPeralta_30_port_o_0_7;
  wire       [0:0]    sbox_AES_BoyarPeralta_30_port_o_1_0;
  wire       [0:0]    sbox_AES_BoyarPeralta_30_port_o_1_1;
  wire       [0:0]    sbox_AES_BoyarPeralta_30_port_o_1_2;
  wire       [0:0]    sbox_AES_BoyarPeralta_30_port_o_1_3;
  wire       [0:0]    sbox_AES_BoyarPeralta_30_port_o_1_4;
  wire       [0:0]    sbox_AES_BoyarPeralta_30_port_o_1_5;
  wire       [0:0]    sbox_AES_BoyarPeralta_30_port_o_1_6;
  wire       [0:0]    sbox_AES_BoyarPeralta_30_port_o_1_7;
  wire       [0:0]    sbox_AES_BoyarPeralta_30_port_o_2_0;
  wire       [0:0]    sbox_AES_BoyarPeralta_30_port_o_2_1;
  wire       [0:0]    sbox_AES_BoyarPeralta_30_port_o_2_2;
  wire       [0:0]    sbox_AES_BoyarPeralta_30_port_o_2_3;
  wire       [0:0]    sbox_AES_BoyarPeralta_30_port_o_2_4;
  wire       [0:0]    sbox_AES_BoyarPeralta_30_port_o_2_5;
  wire       [0:0]    sbox_AES_BoyarPeralta_30_port_o_2_6;
  wire       [0:0]    sbox_AES_BoyarPeralta_30_port_o_2_7;
  wire       [0:0]    sbox_AES_BoyarPeralta_30_port_o_3_0;
  wire       [0:0]    sbox_AES_BoyarPeralta_30_port_o_3_1;
  wire       [0:0]    sbox_AES_BoyarPeralta_30_port_o_3_2;
  wire       [0:0]    sbox_AES_BoyarPeralta_30_port_o_3_3;
  wire       [0:0]    sbox_AES_BoyarPeralta_30_port_o_3_4;
  wire       [0:0]    sbox_AES_BoyarPeralta_30_port_o_3_5;
  wire       [0:0]    sbox_AES_BoyarPeralta_30_port_o_3_6;
  wire       [0:0]    sbox_AES_BoyarPeralta_30_port_o_3_7;
  wire       [0:0]    sbox_AES_BoyarPeralta_31_port_o_0_0;
  wire       [0:0]    sbox_AES_BoyarPeralta_31_port_o_0_1;
  wire       [0:0]    sbox_AES_BoyarPeralta_31_port_o_0_2;
  wire       [0:0]    sbox_AES_BoyarPeralta_31_port_o_0_3;
  wire       [0:0]    sbox_AES_BoyarPeralta_31_port_o_0_4;
  wire       [0:0]    sbox_AES_BoyarPeralta_31_port_o_0_5;
  wire       [0:0]    sbox_AES_BoyarPeralta_31_port_o_0_6;
  wire       [0:0]    sbox_AES_BoyarPeralta_31_port_o_0_7;
  wire       [0:0]    sbox_AES_BoyarPeralta_31_port_o_1_0;
  wire       [0:0]    sbox_AES_BoyarPeralta_31_port_o_1_1;
  wire       [0:0]    sbox_AES_BoyarPeralta_31_port_o_1_2;
  wire       [0:0]    sbox_AES_BoyarPeralta_31_port_o_1_3;
  wire       [0:0]    sbox_AES_BoyarPeralta_31_port_o_1_4;
  wire       [0:0]    sbox_AES_BoyarPeralta_31_port_o_1_5;
  wire       [0:0]    sbox_AES_BoyarPeralta_31_port_o_1_6;
  wire       [0:0]    sbox_AES_BoyarPeralta_31_port_o_1_7;
  wire       [0:0]    sbox_AES_BoyarPeralta_31_port_o_2_0;
  wire       [0:0]    sbox_AES_BoyarPeralta_31_port_o_2_1;
  wire       [0:0]    sbox_AES_BoyarPeralta_31_port_o_2_2;
  wire       [0:0]    sbox_AES_BoyarPeralta_31_port_o_2_3;
  wire       [0:0]    sbox_AES_BoyarPeralta_31_port_o_2_4;
  wire       [0:0]    sbox_AES_BoyarPeralta_31_port_o_2_5;
  wire       [0:0]    sbox_AES_BoyarPeralta_31_port_o_2_6;
  wire       [0:0]    sbox_AES_BoyarPeralta_31_port_o_2_7;
  wire       [0:0]    sbox_AES_BoyarPeralta_31_port_o_3_0;
  wire       [0:0]    sbox_AES_BoyarPeralta_31_port_o_3_1;
  wire       [0:0]    sbox_AES_BoyarPeralta_31_port_o_3_2;
  wire       [0:0]    sbox_AES_BoyarPeralta_31_port_o_3_3;
  wire       [0:0]    sbox_AES_BoyarPeralta_31_port_o_3_4;
  wire       [0:0]    sbox_AES_BoyarPeralta_31_port_o_3_5;
  wire       [0:0]    sbox_AES_BoyarPeralta_31_port_o_3_6;
  wire       [0:0]    sbox_AES_BoyarPeralta_31_port_o_3_7;
  wire       [0:0]    shiftRows_port_state_out_0_0_0;
  wire       [0:0]    shiftRows_port_state_out_0_0_1;
  wire       [0:0]    shiftRows_port_state_out_0_0_2;
  wire       [0:0]    shiftRows_port_state_out_0_0_3;
  wire       [0:0]    shiftRows_port_state_out_0_0_4;
  wire       [0:0]    shiftRows_port_state_out_0_0_5;
  wire       [0:0]    shiftRows_port_state_out_0_0_6;
  wire       [0:0]    shiftRows_port_state_out_0_0_7;
  wire       [0:0]    shiftRows_port_state_out_0_1_0;
  wire       [0:0]    shiftRows_port_state_out_0_1_1;
  wire       [0:0]    shiftRows_port_state_out_0_1_2;
  wire       [0:0]    shiftRows_port_state_out_0_1_3;
  wire       [0:0]    shiftRows_port_state_out_0_1_4;
  wire       [0:0]    shiftRows_port_state_out_0_1_5;
  wire       [0:0]    shiftRows_port_state_out_0_1_6;
  wire       [0:0]    shiftRows_port_state_out_0_1_7;
  wire       [0:0]    shiftRows_port_state_out_0_2_0;
  wire       [0:0]    shiftRows_port_state_out_0_2_1;
  wire       [0:0]    shiftRows_port_state_out_0_2_2;
  wire       [0:0]    shiftRows_port_state_out_0_2_3;
  wire       [0:0]    shiftRows_port_state_out_0_2_4;
  wire       [0:0]    shiftRows_port_state_out_0_2_5;
  wire       [0:0]    shiftRows_port_state_out_0_2_6;
  wire       [0:0]    shiftRows_port_state_out_0_2_7;
  wire       [0:0]    shiftRows_port_state_out_0_3_0;
  wire       [0:0]    shiftRows_port_state_out_0_3_1;
  wire       [0:0]    shiftRows_port_state_out_0_3_2;
  wire       [0:0]    shiftRows_port_state_out_0_3_3;
  wire       [0:0]    shiftRows_port_state_out_0_3_4;
  wire       [0:0]    shiftRows_port_state_out_0_3_5;
  wire       [0:0]    shiftRows_port_state_out_0_3_6;
  wire       [0:0]    shiftRows_port_state_out_0_3_7;
  wire       [0:0]    shiftRows_port_state_out_1_0_0;
  wire       [0:0]    shiftRows_port_state_out_1_0_1;
  wire       [0:0]    shiftRows_port_state_out_1_0_2;
  wire       [0:0]    shiftRows_port_state_out_1_0_3;
  wire       [0:0]    shiftRows_port_state_out_1_0_4;
  wire       [0:0]    shiftRows_port_state_out_1_0_5;
  wire       [0:0]    shiftRows_port_state_out_1_0_6;
  wire       [0:0]    shiftRows_port_state_out_1_0_7;
  wire       [0:0]    shiftRows_port_state_out_1_1_0;
  wire       [0:0]    shiftRows_port_state_out_1_1_1;
  wire       [0:0]    shiftRows_port_state_out_1_1_2;
  wire       [0:0]    shiftRows_port_state_out_1_1_3;
  wire       [0:0]    shiftRows_port_state_out_1_1_4;
  wire       [0:0]    shiftRows_port_state_out_1_1_5;
  wire       [0:0]    shiftRows_port_state_out_1_1_6;
  wire       [0:0]    shiftRows_port_state_out_1_1_7;
  wire       [0:0]    shiftRows_port_state_out_1_2_0;
  wire       [0:0]    shiftRows_port_state_out_1_2_1;
  wire       [0:0]    shiftRows_port_state_out_1_2_2;
  wire       [0:0]    shiftRows_port_state_out_1_2_3;
  wire       [0:0]    shiftRows_port_state_out_1_2_4;
  wire       [0:0]    shiftRows_port_state_out_1_2_5;
  wire       [0:0]    shiftRows_port_state_out_1_2_6;
  wire       [0:0]    shiftRows_port_state_out_1_2_7;
  wire       [0:0]    shiftRows_port_state_out_1_3_0;
  wire       [0:0]    shiftRows_port_state_out_1_3_1;
  wire       [0:0]    shiftRows_port_state_out_1_3_2;
  wire       [0:0]    shiftRows_port_state_out_1_3_3;
  wire       [0:0]    shiftRows_port_state_out_1_3_4;
  wire       [0:0]    shiftRows_port_state_out_1_3_5;
  wire       [0:0]    shiftRows_port_state_out_1_3_6;
  wire       [0:0]    shiftRows_port_state_out_1_3_7;
  wire       [0:0]    shiftRows_port_state_out_2_0_0;
  wire       [0:0]    shiftRows_port_state_out_2_0_1;
  wire       [0:0]    shiftRows_port_state_out_2_0_2;
  wire       [0:0]    shiftRows_port_state_out_2_0_3;
  wire       [0:0]    shiftRows_port_state_out_2_0_4;
  wire       [0:0]    shiftRows_port_state_out_2_0_5;
  wire       [0:0]    shiftRows_port_state_out_2_0_6;
  wire       [0:0]    shiftRows_port_state_out_2_0_7;
  wire       [0:0]    shiftRows_port_state_out_2_1_0;
  wire       [0:0]    shiftRows_port_state_out_2_1_1;
  wire       [0:0]    shiftRows_port_state_out_2_1_2;
  wire       [0:0]    shiftRows_port_state_out_2_1_3;
  wire       [0:0]    shiftRows_port_state_out_2_1_4;
  wire       [0:0]    shiftRows_port_state_out_2_1_5;
  wire       [0:0]    shiftRows_port_state_out_2_1_6;
  wire       [0:0]    shiftRows_port_state_out_2_1_7;
  wire       [0:0]    shiftRows_port_state_out_2_2_0;
  wire       [0:0]    shiftRows_port_state_out_2_2_1;
  wire       [0:0]    shiftRows_port_state_out_2_2_2;
  wire       [0:0]    shiftRows_port_state_out_2_2_3;
  wire       [0:0]    shiftRows_port_state_out_2_2_4;
  wire       [0:0]    shiftRows_port_state_out_2_2_5;
  wire       [0:0]    shiftRows_port_state_out_2_2_6;
  wire       [0:0]    shiftRows_port_state_out_2_2_7;
  wire       [0:0]    shiftRows_port_state_out_2_3_0;
  wire       [0:0]    shiftRows_port_state_out_2_3_1;
  wire       [0:0]    shiftRows_port_state_out_2_3_2;
  wire       [0:0]    shiftRows_port_state_out_2_3_3;
  wire       [0:0]    shiftRows_port_state_out_2_3_4;
  wire       [0:0]    shiftRows_port_state_out_2_3_5;
  wire       [0:0]    shiftRows_port_state_out_2_3_6;
  wire       [0:0]    shiftRows_port_state_out_2_3_7;
  wire       [0:0]    shiftRows_port_state_out_3_0_0;
  wire       [0:0]    shiftRows_port_state_out_3_0_1;
  wire       [0:0]    shiftRows_port_state_out_3_0_2;
  wire       [0:0]    shiftRows_port_state_out_3_0_3;
  wire       [0:0]    shiftRows_port_state_out_3_0_4;
  wire       [0:0]    shiftRows_port_state_out_3_0_5;
  wire       [0:0]    shiftRows_port_state_out_3_0_6;
  wire       [0:0]    shiftRows_port_state_out_3_0_7;
  wire       [0:0]    shiftRows_port_state_out_3_1_0;
  wire       [0:0]    shiftRows_port_state_out_3_1_1;
  wire       [0:0]    shiftRows_port_state_out_3_1_2;
  wire       [0:0]    shiftRows_port_state_out_3_1_3;
  wire       [0:0]    shiftRows_port_state_out_3_1_4;
  wire       [0:0]    shiftRows_port_state_out_3_1_5;
  wire       [0:0]    shiftRows_port_state_out_3_1_6;
  wire       [0:0]    shiftRows_port_state_out_3_1_7;
  wire       [0:0]    shiftRows_port_state_out_3_2_0;
  wire       [0:0]    shiftRows_port_state_out_3_2_1;
  wire       [0:0]    shiftRows_port_state_out_3_2_2;
  wire       [0:0]    shiftRows_port_state_out_3_2_3;
  wire       [0:0]    shiftRows_port_state_out_3_2_4;
  wire       [0:0]    shiftRows_port_state_out_3_2_5;
  wire       [0:0]    shiftRows_port_state_out_3_2_6;
  wire       [0:0]    shiftRows_port_state_out_3_2_7;
  wire       [0:0]    shiftRows_port_state_out_3_3_0;
  wire       [0:0]    shiftRows_port_state_out_3_3_1;
  wire       [0:0]    shiftRows_port_state_out_3_3_2;
  wire       [0:0]    shiftRows_port_state_out_3_3_3;
  wire       [0:0]    shiftRows_port_state_out_3_3_4;
  wire       [0:0]    shiftRows_port_state_out_3_3_5;
  wire       [0:0]    shiftRows_port_state_out_3_3_6;
  wire       [0:0]    shiftRows_port_state_out_3_3_7;
  wire       [0:0]    shiftRows_port_state_out_4_0_0;
  wire       [0:0]    shiftRows_port_state_out_4_0_1;
  wire       [0:0]    shiftRows_port_state_out_4_0_2;
  wire       [0:0]    shiftRows_port_state_out_4_0_3;
  wire       [0:0]    shiftRows_port_state_out_4_0_4;
  wire       [0:0]    shiftRows_port_state_out_4_0_5;
  wire       [0:0]    shiftRows_port_state_out_4_0_6;
  wire       [0:0]    shiftRows_port_state_out_4_0_7;
  wire       [0:0]    shiftRows_port_state_out_4_1_0;
  wire       [0:0]    shiftRows_port_state_out_4_1_1;
  wire       [0:0]    shiftRows_port_state_out_4_1_2;
  wire       [0:0]    shiftRows_port_state_out_4_1_3;
  wire       [0:0]    shiftRows_port_state_out_4_1_4;
  wire       [0:0]    shiftRows_port_state_out_4_1_5;
  wire       [0:0]    shiftRows_port_state_out_4_1_6;
  wire       [0:0]    shiftRows_port_state_out_4_1_7;
  wire       [0:0]    shiftRows_port_state_out_4_2_0;
  wire       [0:0]    shiftRows_port_state_out_4_2_1;
  wire       [0:0]    shiftRows_port_state_out_4_2_2;
  wire       [0:0]    shiftRows_port_state_out_4_2_3;
  wire       [0:0]    shiftRows_port_state_out_4_2_4;
  wire       [0:0]    shiftRows_port_state_out_4_2_5;
  wire       [0:0]    shiftRows_port_state_out_4_2_6;
  wire       [0:0]    shiftRows_port_state_out_4_2_7;
  wire       [0:0]    shiftRows_port_state_out_4_3_0;
  wire       [0:0]    shiftRows_port_state_out_4_3_1;
  wire       [0:0]    shiftRows_port_state_out_4_3_2;
  wire       [0:0]    shiftRows_port_state_out_4_3_3;
  wire       [0:0]    shiftRows_port_state_out_4_3_4;
  wire       [0:0]    shiftRows_port_state_out_4_3_5;
  wire       [0:0]    shiftRows_port_state_out_4_3_6;
  wire       [0:0]    shiftRows_port_state_out_4_3_7;
  wire       [0:0]    shiftRows_port_state_out_5_0_0;
  wire       [0:0]    shiftRows_port_state_out_5_0_1;
  wire       [0:0]    shiftRows_port_state_out_5_0_2;
  wire       [0:0]    shiftRows_port_state_out_5_0_3;
  wire       [0:0]    shiftRows_port_state_out_5_0_4;
  wire       [0:0]    shiftRows_port_state_out_5_0_5;
  wire       [0:0]    shiftRows_port_state_out_5_0_6;
  wire       [0:0]    shiftRows_port_state_out_5_0_7;
  wire       [0:0]    shiftRows_port_state_out_5_1_0;
  wire       [0:0]    shiftRows_port_state_out_5_1_1;
  wire       [0:0]    shiftRows_port_state_out_5_1_2;
  wire       [0:0]    shiftRows_port_state_out_5_1_3;
  wire       [0:0]    shiftRows_port_state_out_5_1_4;
  wire       [0:0]    shiftRows_port_state_out_5_1_5;
  wire       [0:0]    shiftRows_port_state_out_5_1_6;
  wire       [0:0]    shiftRows_port_state_out_5_1_7;
  wire       [0:0]    shiftRows_port_state_out_5_2_0;
  wire       [0:0]    shiftRows_port_state_out_5_2_1;
  wire       [0:0]    shiftRows_port_state_out_5_2_2;
  wire       [0:0]    shiftRows_port_state_out_5_2_3;
  wire       [0:0]    shiftRows_port_state_out_5_2_4;
  wire       [0:0]    shiftRows_port_state_out_5_2_5;
  wire       [0:0]    shiftRows_port_state_out_5_2_6;
  wire       [0:0]    shiftRows_port_state_out_5_2_7;
  wire       [0:0]    shiftRows_port_state_out_5_3_0;
  wire       [0:0]    shiftRows_port_state_out_5_3_1;
  wire       [0:0]    shiftRows_port_state_out_5_3_2;
  wire       [0:0]    shiftRows_port_state_out_5_3_3;
  wire       [0:0]    shiftRows_port_state_out_5_3_4;
  wire       [0:0]    shiftRows_port_state_out_5_3_5;
  wire       [0:0]    shiftRows_port_state_out_5_3_6;
  wire       [0:0]    shiftRows_port_state_out_5_3_7;
  wire       [0:0]    shiftRows_port_state_out_6_0_0;
  wire       [0:0]    shiftRows_port_state_out_6_0_1;
  wire       [0:0]    shiftRows_port_state_out_6_0_2;
  wire       [0:0]    shiftRows_port_state_out_6_0_3;
  wire       [0:0]    shiftRows_port_state_out_6_0_4;
  wire       [0:0]    shiftRows_port_state_out_6_0_5;
  wire       [0:0]    shiftRows_port_state_out_6_0_6;
  wire       [0:0]    shiftRows_port_state_out_6_0_7;
  wire       [0:0]    shiftRows_port_state_out_6_1_0;
  wire       [0:0]    shiftRows_port_state_out_6_1_1;
  wire       [0:0]    shiftRows_port_state_out_6_1_2;
  wire       [0:0]    shiftRows_port_state_out_6_1_3;
  wire       [0:0]    shiftRows_port_state_out_6_1_4;
  wire       [0:0]    shiftRows_port_state_out_6_1_5;
  wire       [0:0]    shiftRows_port_state_out_6_1_6;
  wire       [0:0]    shiftRows_port_state_out_6_1_7;
  wire       [0:0]    shiftRows_port_state_out_6_2_0;
  wire       [0:0]    shiftRows_port_state_out_6_2_1;
  wire       [0:0]    shiftRows_port_state_out_6_2_2;
  wire       [0:0]    shiftRows_port_state_out_6_2_3;
  wire       [0:0]    shiftRows_port_state_out_6_2_4;
  wire       [0:0]    shiftRows_port_state_out_6_2_5;
  wire       [0:0]    shiftRows_port_state_out_6_2_6;
  wire       [0:0]    shiftRows_port_state_out_6_2_7;
  wire       [0:0]    shiftRows_port_state_out_6_3_0;
  wire       [0:0]    shiftRows_port_state_out_6_3_1;
  wire       [0:0]    shiftRows_port_state_out_6_3_2;
  wire       [0:0]    shiftRows_port_state_out_6_3_3;
  wire       [0:0]    shiftRows_port_state_out_6_3_4;
  wire       [0:0]    shiftRows_port_state_out_6_3_5;
  wire       [0:0]    shiftRows_port_state_out_6_3_6;
  wire       [0:0]    shiftRows_port_state_out_6_3_7;
  wire       [0:0]    shiftRows_port_state_out_7_0_0;
  wire       [0:0]    shiftRows_port_state_out_7_0_1;
  wire       [0:0]    shiftRows_port_state_out_7_0_2;
  wire       [0:0]    shiftRows_port_state_out_7_0_3;
  wire       [0:0]    shiftRows_port_state_out_7_0_4;
  wire       [0:0]    shiftRows_port_state_out_7_0_5;
  wire       [0:0]    shiftRows_port_state_out_7_0_6;
  wire       [0:0]    shiftRows_port_state_out_7_0_7;
  wire       [0:0]    shiftRows_port_state_out_7_1_0;
  wire       [0:0]    shiftRows_port_state_out_7_1_1;
  wire       [0:0]    shiftRows_port_state_out_7_1_2;
  wire       [0:0]    shiftRows_port_state_out_7_1_3;
  wire       [0:0]    shiftRows_port_state_out_7_1_4;
  wire       [0:0]    shiftRows_port_state_out_7_1_5;
  wire       [0:0]    shiftRows_port_state_out_7_1_6;
  wire       [0:0]    shiftRows_port_state_out_7_1_7;
  wire       [0:0]    shiftRows_port_state_out_7_2_0;
  wire       [0:0]    shiftRows_port_state_out_7_2_1;
  wire       [0:0]    shiftRows_port_state_out_7_2_2;
  wire       [0:0]    shiftRows_port_state_out_7_2_3;
  wire       [0:0]    shiftRows_port_state_out_7_2_4;
  wire       [0:0]    shiftRows_port_state_out_7_2_5;
  wire       [0:0]    shiftRows_port_state_out_7_2_6;
  wire       [0:0]    shiftRows_port_state_out_7_2_7;
  wire       [0:0]    shiftRows_port_state_out_7_3_0;
  wire       [0:0]    shiftRows_port_state_out_7_3_1;
  wire       [0:0]    shiftRows_port_state_out_7_3_2;
  wire       [0:0]    shiftRows_port_state_out_7_3_3;
  wire       [0:0]    shiftRows_port_state_out_7_3_4;
  wire       [0:0]    shiftRows_port_state_out_7_3_5;
  wire       [0:0]    shiftRows_port_state_out_7_3_6;
  wire       [0:0]    shiftRows_port_state_out_7_3_7;
  wire       [0:0]    shiftRows_port_state_out_8_0_0;
  wire       [0:0]    shiftRows_port_state_out_8_0_1;
  wire       [0:0]    shiftRows_port_state_out_8_0_2;
  wire       [0:0]    shiftRows_port_state_out_8_0_3;
  wire       [0:0]    shiftRows_port_state_out_8_0_4;
  wire       [0:0]    shiftRows_port_state_out_8_0_5;
  wire       [0:0]    shiftRows_port_state_out_8_0_6;
  wire       [0:0]    shiftRows_port_state_out_8_0_7;
  wire       [0:0]    shiftRows_port_state_out_8_1_0;
  wire       [0:0]    shiftRows_port_state_out_8_1_1;
  wire       [0:0]    shiftRows_port_state_out_8_1_2;
  wire       [0:0]    shiftRows_port_state_out_8_1_3;
  wire       [0:0]    shiftRows_port_state_out_8_1_4;
  wire       [0:0]    shiftRows_port_state_out_8_1_5;
  wire       [0:0]    shiftRows_port_state_out_8_1_6;
  wire       [0:0]    shiftRows_port_state_out_8_1_7;
  wire       [0:0]    shiftRows_port_state_out_8_2_0;
  wire       [0:0]    shiftRows_port_state_out_8_2_1;
  wire       [0:0]    shiftRows_port_state_out_8_2_2;
  wire       [0:0]    shiftRows_port_state_out_8_2_3;
  wire       [0:0]    shiftRows_port_state_out_8_2_4;
  wire       [0:0]    shiftRows_port_state_out_8_2_5;
  wire       [0:0]    shiftRows_port_state_out_8_2_6;
  wire       [0:0]    shiftRows_port_state_out_8_2_7;
  wire       [0:0]    shiftRows_port_state_out_8_3_0;
  wire       [0:0]    shiftRows_port_state_out_8_3_1;
  wire       [0:0]    shiftRows_port_state_out_8_3_2;
  wire       [0:0]    shiftRows_port_state_out_8_3_3;
  wire       [0:0]    shiftRows_port_state_out_8_3_4;
  wire       [0:0]    shiftRows_port_state_out_8_3_5;
  wire       [0:0]    shiftRows_port_state_out_8_3_6;
  wire       [0:0]    shiftRows_port_state_out_8_3_7;
  wire       [0:0]    shiftRows_port_state_out_9_0_0;
  wire       [0:0]    shiftRows_port_state_out_9_0_1;
  wire       [0:0]    shiftRows_port_state_out_9_0_2;
  wire       [0:0]    shiftRows_port_state_out_9_0_3;
  wire       [0:0]    shiftRows_port_state_out_9_0_4;
  wire       [0:0]    shiftRows_port_state_out_9_0_5;
  wire       [0:0]    shiftRows_port_state_out_9_0_6;
  wire       [0:0]    shiftRows_port_state_out_9_0_7;
  wire       [0:0]    shiftRows_port_state_out_9_1_0;
  wire       [0:0]    shiftRows_port_state_out_9_1_1;
  wire       [0:0]    shiftRows_port_state_out_9_1_2;
  wire       [0:0]    shiftRows_port_state_out_9_1_3;
  wire       [0:0]    shiftRows_port_state_out_9_1_4;
  wire       [0:0]    shiftRows_port_state_out_9_1_5;
  wire       [0:0]    shiftRows_port_state_out_9_1_6;
  wire       [0:0]    shiftRows_port_state_out_9_1_7;
  wire       [0:0]    shiftRows_port_state_out_9_2_0;
  wire       [0:0]    shiftRows_port_state_out_9_2_1;
  wire       [0:0]    shiftRows_port_state_out_9_2_2;
  wire       [0:0]    shiftRows_port_state_out_9_2_3;
  wire       [0:0]    shiftRows_port_state_out_9_2_4;
  wire       [0:0]    shiftRows_port_state_out_9_2_5;
  wire       [0:0]    shiftRows_port_state_out_9_2_6;
  wire       [0:0]    shiftRows_port_state_out_9_2_7;
  wire       [0:0]    shiftRows_port_state_out_9_3_0;
  wire       [0:0]    shiftRows_port_state_out_9_3_1;
  wire       [0:0]    shiftRows_port_state_out_9_3_2;
  wire       [0:0]    shiftRows_port_state_out_9_3_3;
  wire       [0:0]    shiftRows_port_state_out_9_3_4;
  wire       [0:0]    shiftRows_port_state_out_9_3_5;
  wire       [0:0]    shiftRows_port_state_out_9_3_6;
  wire       [0:0]    shiftRows_port_state_out_9_3_7;
  wire       [0:0]    shiftRows_port_state_out_10_0_0;
  wire       [0:0]    shiftRows_port_state_out_10_0_1;
  wire       [0:0]    shiftRows_port_state_out_10_0_2;
  wire       [0:0]    shiftRows_port_state_out_10_0_3;
  wire       [0:0]    shiftRows_port_state_out_10_0_4;
  wire       [0:0]    shiftRows_port_state_out_10_0_5;
  wire       [0:0]    shiftRows_port_state_out_10_0_6;
  wire       [0:0]    shiftRows_port_state_out_10_0_7;
  wire       [0:0]    shiftRows_port_state_out_10_1_0;
  wire       [0:0]    shiftRows_port_state_out_10_1_1;
  wire       [0:0]    shiftRows_port_state_out_10_1_2;
  wire       [0:0]    shiftRows_port_state_out_10_1_3;
  wire       [0:0]    shiftRows_port_state_out_10_1_4;
  wire       [0:0]    shiftRows_port_state_out_10_1_5;
  wire       [0:0]    shiftRows_port_state_out_10_1_6;
  wire       [0:0]    shiftRows_port_state_out_10_1_7;
  wire       [0:0]    shiftRows_port_state_out_10_2_0;
  wire       [0:0]    shiftRows_port_state_out_10_2_1;
  wire       [0:0]    shiftRows_port_state_out_10_2_2;
  wire       [0:0]    shiftRows_port_state_out_10_2_3;
  wire       [0:0]    shiftRows_port_state_out_10_2_4;
  wire       [0:0]    shiftRows_port_state_out_10_2_5;
  wire       [0:0]    shiftRows_port_state_out_10_2_6;
  wire       [0:0]    shiftRows_port_state_out_10_2_7;
  wire       [0:0]    shiftRows_port_state_out_10_3_0;
  wire       [0:0]    shiftRows_port_state_out_10_3_1;
  wire       [0:0]    shiftRows_port_state_out_10_3_2;
  wire       [0:0]    shiftRows_port_state_out_10_3_3;
  wire       [0:0]    shiftRows_port_state_out_10_3_4;
  wire       [0:0]    shiftRows_port_state_out_10_3_5;
  wire       [0:0]    shiftRows_port_state_out_10_3_6;
  wire       [0:0]    shiftRows_port_state_out_10_3_7;
  wire       [0:0]    shiftRows_port_state_out_11_0_0;
  wire       [0:0]    shiftRows_port_state_out_11_0_1;
  wire       [0:0]    shiftRows_port_state_out_11_0_2;
  wire       [0:0]    shiftRows_port_state_out_11_0_3;
  wire       [0:0]    shiftRows_port_state_out_11_0_4;
  wire       [0:0]    shiftRows_port_state_out_11_0_5;
  wire       [0:0]    shiftRows_port_state_out_11_0_6;
  wire       [0:0]    shiftRows_port_state_out_11_0_7;
  wire       [0:0]    shiftRows_port_state_out_11_1_0;
  wire       [0:0]    shiftRows_port_state_out_11_1_1;
  wire       [0:0]    shiftRows_port_state_out_11_1_2;
  wire       [0:0]    shiftRows_port_state_out_11_1_3;
  wire       [0:0]    shiftRows_port_state_out_11_1_4;
  wire       [0:0]    shiftRows_port_state_out_11_1_5;
  wire       [0:0]    shiftRows_port_state_out_11_1_6;
  wire       [0:0]    shiftRows_port_state_out_11_1_7;
  wire       [0:0]    shiftRows_port_state_out_11_2_0;
  wire       [0:0]    shiftRows_port_state_out_11_2_1;
  wire       [0:0]    shiftRows_port_state_out_11_2_2;
  wire       [0:0]    shiftRows_port_state_out_11_2_3;
  wire       [0:0]    shiftRows_port_state_out_11_2_4;
  wire       [0:0]    shiftRows_port_state_out_11_2_5;
  wire       [0:0]    shiftRows_port_state_out_11_2_6;
  wire       [0:0]    shiftRows_port_state_out_11_2_7;
  wire       [0:0]    shiftRows_port_state_out_11_3_0;
  wire       [0:0]    shiftRows_port_state_out_11_3_1;
  wire       [0:0]    shiftRows_port_state_out_11_3_2;
  wire       [0:0]    shiftRows_port_state_out_11_3_3;
  wire       [0:0]    shiftRows_port_state_out_11_3_4;
  wire       [0:0]    shiftRows_port_state_out_11_3_5;
  wire       [0:0]    shiftRows_port_state_out_11_3_6;
  wire       [0:0]    shiftRows_port_state_out_11_3_7;
  wire       [0:0]    shiftRows_port_state_out_12_0_0;
  wire       [0:0]    shiftRows_port_state_out_12_0_1;
  wire       [0:0]    shiftRows_port_state_out_12_0_2;
  wire       [0:0]    shiftRows_port_state_out_12_0_3;
  wire       [0:0]    shiftRows_port_state_out_12_0_4;
  wire       [0:0]    shiftRows_port_state_out_12_0_5;
  wire       [0:0]    shiftRows_port_state_out_12_0_6;
  wire       [0:0]    shiftRows_port_state_out_12_0_7;
  wire       [0:0]    shiftRows_port_state_out_12_1_0;
  wire       [0:0]    shiftRows_port_state_out_12_1_1;
  wire       [0:0]    shiftRows_port_state_out_12_1_2;
  wire       [0:0]    shiftRows_port_state_out_12_1_3;
  wire       [0:0]    shiftRows_port_state_out_12_1_4;
  wire       [0:0]    shiftRows_port_state_out_12_1_5;
  wire       [0:0]    shiftRows_port_state_out_12_1_6;
  wire       [0:0]    shiftRows_port_state_out_12_1_7;
  wire       [0:0]    shiftRows_port_state_out_12_2_0;
  wire       [0:0]    shiftRows_port_state_out_12_2_1;
  wire       [0:0]    shiftRows_port_state_out_12_2_2;
  wire       [0:0]    shiftRows_port_state_out_12_2_3;
  wire       [0:0]    shiftRows_port_state_out_12_2_4;
  wire       [0:0]    shiftRows_port_state_out_12_2_5;
  wire       [0:0]    shiftRows_port_state_out_12_2_6;
  wire       [0:0]    shiftRows_port_state_out_12_2_7;
  wire       [0:0]    shiftRows_port_state_out_12_3_0;
  wire       [0:0]    shiftRows_port_state_out_12_3_1;
  wire       [0:0]    shiftRows_port_state_out_12_3_2;
  wire       [0:0]    shiftRows_port_state_out_12_3_3;
  wire       [0:0]    shiftRows_port_state_out_12_3_4;
  wire       [0:0]    shiftRows_port_state_out_12_3_5;
  wire       [0:0]    shiftRows_port_state_out_12_3_6;
  wire       [0:0]    shiftRows_port_state_out_12_3_7;
  wire       [0:0]    shiftRows_port_state_out_13_0_0;
  wire       [0:0]    shiftRows_port_state_out_13_0_1;
  wire       [0:0]    shiftRows_port_state_out_13_0_2;
  wire       [0:0]    shiftRows_port_state_out_13_0_3;
  wire       [0:0]    shiftRows_port_state_out_13_0_4;
  wire       [0:0]    shiftRows_port_state_out_13_0_5;
  wire       [0:0]    shiftRows_port_state_out_13_0_6;
  wire       [0:0]    shiftRows_port_state_out_13_0_7;
  wire       [0:0]    shiftRows_port_state_out_13_1_0;
  wire       [0:0]    shiftRows_port_state_out_13_1_1;
  wire       [0:0]    shiftRows_port_state_out_13_1_2;
  wire       [0:0]    shiftRows_port_state_out_13_1_3;
  wire       [0:0]    shiftRows_port_state_out_13_1_4;
  wire       [0:0]    shiftRows_port_state_out_13_1_5;
  wire       [0:0]    shiftRows_port_state_out_13_1_6;
  wire       [0:0]    shiftRows_port_state_out_13_1_7;
  wire       [0:0]    shiftRows_port_state_out_13_2_0;
  wire       [0:0]    shiftRows_port_state_out_13_2_1;
  wire       [0:0]    shiftRows_port_state_out_13_2_2;
  wire       [0:0]    shiftRows_port_state_out_13_2_3;
  wire       [0:0]    shiftRows_port_state_out_13_2_4;
  wire       [0:0]    shiftRows_port_state_out_13_2_5;
  wire       [0:0]    shiftRows_port_state_out_13_2_6;
  wire       [0:0]    shiftRows_port_state_out_13_2_7;
  wire       [0:0]    shiftRows_port_state_out_13_3_0;
  wire       [0:0]    shiftRows_port_state_out_13_3_1;
  wire       [0:0]    shiftRows_port_state_out_13_3_2;
  wire       [0:0]    shiftRows_port_state_out_13_3_3;
  wire       [0:0]    shiftRows_port_state_out_13_3_4;
  wire       [0:0]    shiftRows_port_state_out_13_3_5;
  wire       [0:0]    shiftRows_port_state_out_13_3_6;
  wire       [0:0]    shiftRows_port_state_out_13_3_7;
  wire       [0:0]    shiftRows_port_state_out_14_0_0;
  wire       [0:0]    shiftRows_port_state_out_14_0_1;
  wire       [0:0]    shiftRows_port_state_out_14_0_2;
  wire       [0:0]    shiftRows_port_state_out_14_0_3;
  wire       [0:0]    shiftRows_port_state_out_14_0_4;
  wire       [0:0]    shiftRows_port_state_out_14_0_5;
  wire       [0:0]    shiftRows_port_state_out_14_0_6;
  wire       [0:0]    shiftRows_port_state_out_14_0_7;
  wire       [0:0]    shiftRows_port_state_out_14_1_0;
  wire       [0:0]    shiftRows_port_state_out_14_1_1;
  wire       [0:0]    shiftRows_port_state_out_14_1_2;
  wire       [0:0]    shiftRows_port_state_out_14_1_3;
  wire       [0:0]    shiftRows_port_state_out_14_1_4;
  wire       [0:0]    shiftRows_port_state_out_14_1_5;
  wire       [0:0]    shiftRows_port_state_out_14_1_6;
  wire       [0:0]    shiftRows_port_state_out_14_1_7;
  wire       [0:0]    shiftRows_port_state_out_14_2_0;
  wire       [0:0]    shiftRows_port_state_out_14_2_1;
  wire       [0:0]    shiftRows_port_state_out_14_2_2;
  wire       [0:0]    shiftRows_port_state_out_14_2_3;
  wire       [0:0]    shiftRows_port_state_out_14_2_4;
  wire       [0:0]    shiftRows_port_state_out_14_2_5;
  wire       [0:0]    shiftRows_port_state_out_14_2_6;
  wire       [0:0]    shiftRows_port_state_out_14_2_7;
  wire       [0:0]    shiftRows_port_state_out_14_3_0;
  wire       [0:0]    shiftRows_port_state_out_14_3_1;
  wire       [0:0]    shiftRows_port_state_out_14_3_2;
  wire       [0:0]    shiftRows_port_state_out_14_3_3;
  wire       [0:0]    shiftRows_port_state_out_14_3_4;
  wire       [0:0]    shiftRows_port_state_out_14_3_5;
  wire       [0:0]    shiftRows_port_state_out_14_3_6;
  wire       [0:0]    shiftRows_port_state_out_14_3_7;
  wire       [0:0]    shiftRows_port_state_out_15_0_0;
  wire       [0:0]    shiftRows_port_state_out_15_0_1;
  wire       [0:0]    shiftRows_port_state_out_15_0_2;
  wire       [0:0]    shiftRows_port_state_out_15_0_3;
  wire       [0:0]    shiftRows_port_state_out_15_0_4;
  wire       [0:0]    shiftRows_port_state_out_15_0_5;
  wire       [0:0]    shiftRows_port_state_out_15_0_6;
  wire       [0:0]    shiftRows_port_state_out_15_0_7;
  wire       [0:0]    shiftRows_port_state_out_15_1_0;
  wire       [0:0]    shiftRows_port_state_out_15_1_1;
  wire       [0:0]    shiftRows_port_state_out_15_1_2;
  wire       [0:0]    shiftRows_port_state_out_15_1_3;
  wire       [0:0]    shiftRows_port_state_out_15_1_4;
  wire       [0:0]    shiftRows_port_state_out_15_1_5;
  wire       [0:0]    shiftRows_port_state_out_15_1_6;
  wire       [0:0]    shiftRows_port_state_out_15_1_7;
  wire       [0:0]    shiftRows_port_state_out_15_2_0;
  wire       [0:0]    shiftRows_port_state_out_15_2_1;
  wire       [0:0]    shiftRows_port_state_out_15_2_2;
  wire       [0:0]    shiftRows_port_state_out_15_2_3;
  wire       [0:0]    shiftRows_port_state_out_15_2_4;
  wire       [0:0]    shiftRows_port_state_out_15_2_5;
  wire       [0:0]    shiftRows_port_state_out_15_2_6;
  wire       [0:0]    shiftRows_port_state_out_15_2_7;
  wire       [0:0]    shiftRows_port_state_out_15_3_0;
  wire       [0:0]    shiftRows_port_state_out_15_3_1;
  wire       [0:0]    shiftRows_port_state_out_15_3_2;
  wire       [0:0]    shiftRows_port_state_out_15_3_3;
  wire       [0:0]    shiftRows_port_state_out_15_3_4;
  wire       [0:0]    shiftRows_port_state_out_15_3_5;
  wire       [0:0]    shiftRows_port_state_out_15_3_6;
  wire       [0:0]    shiftRows_port_state_out_15_3_7;
  wire       [0:0]    mixColumns_port_state_out_0_0_0;
  wire       [0:0]    mixColumns_port_state_out_0_0_1;
  wire       [0:0]    mixColumns_port_state_out_0_0_2;
  wire       [0:0]    mixColumns_port_state_out_0_0_3;
  wire       [0:0]    mixColumns_port_state_out_0_0_4;
  wire       [0:0]    mixColumns_port_state_out_0_0_5;
  wire       [0:0]    mixColumns_port_state_out_0_0_6;
  wire       [0:0]    mixColumns_port_state_out_0_0_7;
  wire       [0:0]    mixColumns_port_state_out_0_1_0;
  wire       [0:0]    mixColumns_port_state_out_0_1_1;
  wire       [0:0]    mixColumns_port_state_out_0_1_2;
  wire       [0:0]    mixColumns_port_state_out_0_1_3;
  wire       [0:0]    mixColumns_port_state_out_0_1_4;
  wire       [0:0]    mixColumns_port_state_out_0_1_5;
  wire       [0:0]    mixColumns_port_state_out_0_1_6;
  wire       [0:0]    mixColumns_port_state_out_0_1_7;
  wire       [0:0]    mixColumns_port_state_out_0_2_0;
  wire       [0:0]    mixColumns_port_state_out_0_2_1;
  wire       [0:0]    mixColumns_port_state_out_0_2_2;
  wire       [0:0]    mixColumns_port_state_out_0_2_3;
  wire       [0:0]    mixColumns_port_state_out_0_2_4;
  wire       [0:0]    mixColumns_port_state_out_0_2_5;
  wire       [0:0]    mixColumns_port_state_out_0_2_6;
  wire       [0:0]    mixColumns_port_state_out_0_2_7;
  wire       [0:0]    mixColumns_port_state_out_0_3_0;
  wire       [0:0]    mixColumns_port_state_out_0_3_1;
  wire       [0:0]    mixColumns_port_state_out_0_3_2;
  wire       [0:0]    mixColumns_port_state_out_0_3_3;
  wire       [0:0]    mixColumns_port_state_out_0_3_4;
  wire       [0:0]    mixColumns_port_state_out_0_3_5;
  wire       [0:0]    mixColumns_port_state_out_0_3_6;
  wire       [0:0]    mixColumns_port_state_out_0_3_7;
  wire       [0:0]    mixColumns_port_state_out_1_0_0;
  wire       [0:0]    mixColumns_port_state_out_1_0_1;
  wire       [0:0]    mixColumns_port_state_out_1_0_2;
  wire       [0:0]    mixColumns_port_state_out_1_0_3;
  wire       [0:0]    mixColumns_port_state_out_1_0_4;
  wire       [0:0]    mixColumns_port_state_out_1_0_5;
  wire       [0:0]    mixColumns_port_state_out_1_0_6;
  wire       [0:0]    mixColumns_port_state_out_1_0_7;
  wire       [0:0]    mixColumns_port_state_out_1_1_0;
  wire       [0:0]    mixColumns_port_state_out_1_1_1;
  wire       [0:0]    mixColumns_port_state_out_1_1_2;
  wire       [0:0]    mixColumns_port_state_out_1_1_3;
  wire       [0:0]    mixColumns_port_state_out_1_1_4;
  wire       [0:0]    mixColumns_port_state_out_1_1_5;
  wire       [0:0]    mixColumns_port_state_out_1_1_6;
  wire       [0:0]    mixColumns_port_state_out_1_1_7;
  wire       [0:0]    mixColumns_port_state_out_1_2_0;
  wire       [0:0]    mixColumns_port_state_out_1_2_1;
  wire       [0:0]    mixColumns_port_state_out_1_2_2;
  wire       [0:0]    mixColumns_port_state_out_1_2_3;
  wire       [0:0]    mixColumns_port_state_out_1_2_4;
  wire       [0:0]    mixColumns_port_state_out_1_2_5;
  wire       [0:0]    mixColumns_port_state_out_1_2_6;
  wire       [0:0]    mixColumns_port_state_out_1_2_7;
  wire       [0:0]    mixColumns_port_state_out_1_3_0;
  wire       [0:0]    mixColumns_port_state_out_1_3_1;
  wire       [0:0]    mixColumns_port_state_out_1_3_2;
  wire       [0:0]    mixColumns_port_state_out_1_3_3;
  wire       [0:0]    mixColumns_port_state_out_1_3_4;
  wire       [0:0]    mixColumns_port_state_out_1_3_5;
  wire       [0:0]    mixColumns_port_state_out_1_3_6;
  wire       [0:0]    mixColumns_port_state_out_1_3_7;
  wire       [0:0]    mixColumns_port_state_out_2_0_0;
  wire       [0:0]    mixColumns_port_state_out_2_0_1;
  wire       [0:0]    mixColumns_port_state_out_2_0_2;
  wire       [0:0]    mixColumns_port_state_out_2_0_3;
  wire       [0:0]    mixColumns_port_state_out_2_0_4;
  wire       [0:0]    mixColumns_port_state_out_2_0_5;
  wire       [0:0]    mixColumns_port_state_out_2_0_6;
  wire       [0:0]    mixColumns_port_state_out_2_0_7;
  wire       [0:0]    mixColumns_port_state_out_2_1_0;
  wire       [0:0]    mixColumns_port_state_out_2_1_1;
  wire       [0:0]    mixColumns_port_state_out_2_1_2;
  wire       [0:0]    mixColumns_port_state_out_2_1_3;
  wire       [0:0]    mixColumns_port_state_out_2_1_4;
  wire       [0:0]    mixColumns_port_state_out_2_1_5;
  wire       [0:0]    mixColumns_port_state_out_2_1_6;
  wire       [0:0]    mixColumns_port_state_out_2_1_7;
  wire       [0:0]    mixColumns_port_state_out_2_2_0;
  wire       [0:0]    mixColumns_port_state_out_2_2_1;
  wire       [0:0]    mixColumns_port_state_out_2_2_2;
  wire       [0:0]    mixColumns_port_state_out_2_2_3;
  wire       [0:0]    mixColumns_port_state_out_2_2_4;
  wire       [0:0]    mixColumns_port_state_out_2_2_5;
  wire       [0:0]    mixColumns_port_state_out_2_2_6;
  wire       [0:0]    mixColumns_port_state_out_2_2_7;
  wire       [0:0]    mixColumns_port_state_out_2_3_0;
  wire       [0:0]    mixColumns_port_state_out_2_3_1;
  wire       [0:0]    mixColumns_port_state_out_2_3_2;
  wire       [0:0]    mixColumns_port_state_out_2_3_3;
  wire       [0:0]    mixColumns_port_state_out_2_3_4;
  wire       [0:0]    mixColumns_port_state_out_2_3_5;
  wire       [0:0]    mixColumns_port_state_out_2_3_6;
  wire       [0:0]    mixColumns_port_state_out_2_3_7;
  wire       [0:0]    mixColumns_port_state_out_3_0_0;
  wire       [0:0]    mixColumns_port_state_out_3_0_1;
  wire       [0:0]    mixColumns_port_state_out_3_0_2;
  wire       [0:0]    mixColumns_port_state_out_3_0_3;
  wire       [0:0]    mixColumns_port_state_out_3_0_4;
  wire       [0:0]    mixColumns_port_state_out_3_0_5;
  wire       [0:0]    mixColumns_port_state_out_3_0_6;
  wire       [0:0]    mixColumns_port_state_out_3_0_7;
  wire       [0:0]    mixColumns_port_state_out_3_1_0;
  wire       [0:0]    mixColumns_port_state_out_3_1_1;
  wire       [0:0]    mixColumns_port_state_out_3_1_2;
  wire       [0:0]    mixColumns_port_state_out_3_1_3;
  wire       [0:0]    mixColumns_port_state_out_3_1_4;
  wire       [0:0]    mixColumns_port_state_out_3_1_5;
  wire       [0:0]    mixColumns_port_state_out_3_1_6;
  wire       [0:0]    mixColumns_port_state_out_3_1_7;
  wire       [0:0]    mixColumns_port_state_out_3_2_0;
  wire       [0:0]    mixColumns_port_state_out_3_2_1;
  wire       [0:0]    mixColumns_port_state_out_3_2_2;
  wire       [0:0]    mixColumns_port_state_out_3_2_3;
  wire       [0:0]    mixColumns_port_state_out_3_2_4;
  wire       [0:0]    mixColumns_port_state_out_3_2_5;
  wire       [0:0]    mixColumns_port_state_out_3_2_6;
  wire       [0:0]    mixColumns_port_state_out_3_2_7;
  wire       [0:0]    mixColumns_port_state_out_3_3_0;
  wire       [0:0]    mixColumns_port_state_out_3_3_1;
  wire       [0:0]    mixColumns_port_state_out_3_3_2;
  wire       [0:0]    mixColumns_port_state_out_3_3_3;
  wire       [0:0]    mixColumns_port_state_out_3_3_4;
  wire       [0:0]    mixColumns_port_state_out_3_3_5;
  wire       [0:0]    mixColumns_port_state_out_3_3_6;
  wire       [0:0]    mixColumns_port_state_out_3_3_7;
  wire       [0:0]    mixColumns_port_state_out_4_0_0;
  wire       [0:0]    mixColumns_port_state_out_4_0_1;
  wire       [0:0]    mixColumns_port_state_out_4_0_2;
  wire       [0:0]    mixColumns_port_state_out_4_0_3;
  wire       [0:0]    mixColumns_port_state_out_4_0_4;
  wire       [0:0]    mixColumns_port_state_out_4_0_5;
  wire       [0:0]    mixColumns_port_state_out_4_0_6;
  wire       [0:0]    mixColumns_port_state_out_4_0_7;
  wire       [0:0]    mixColumns_port_state_out_4_1_0;
  wire       [0:0]    mixColumns_port_state_out_4_1_1;
  wire       [0:0]    mixColumns_port_state_out_4_1_2;
  wire       [0:0]    mixColumns_port_state_out_4_1_3;
  wire       [0:0]    mixColumns_port_state_out_4_1_4;
  wire       [0:0]    mixColumns_port_state_out_4_1_5;
  wire       [0:0]    mixColumns_port_state_out_4_1_6;
  wire       [0:0]    mixColumns_port_state_out_4_1_7;
  wire       [0:0]    mixColumns_port_state_out_4_2_0;
  wire       [0:0]    mixColumns_port_state_out_4_2_1;
  wire       [0:0]    mixColumns_port_state_out_4_2_2;
  wire       [0:0]    mixColumns_port_state_out_4_2_3;
  wire       [0:0]    mixColumns_port_state_out_4_2_4;
  wire       [0:0]    mixColumns_port_state_out_4_2_5;
  wire       [0:0]    mixColumns_port_state_out_4_2_6;
  wire       [0:0]    mixColumns_port_state_out_4_2_7;
  wire       [0:0]    mixColumns_port_state_out_4_3_0;
  wire       [0:0]    mixColumns_port_state_out_4_3_1;
  wire       [0:0]    mixColumns_port_state_out_4_3_2;
  wire       [0:0]    mixColumns_port_state_out_4_3_3;
  wire       [0:0]    mixColumns_port_state_out_4_3_4;
  wire       [0:0]    mixColumns_port_state_out_4_3_5;
  wire       [0:0]    mixColumns_port_state_out_4_3_6;
  wire       [0:0]    mixColumns_port_state_out_4_3_7;
  wire       [0:0]    mixColumns_port_state_out_5_0_0;
  wire       [0:0]    mixColumns_port_state_out_5_0_1;
  wire       [0:0]    mixColumns_port_state_out_5_0_2;
  wire       [0:0]    mixColumns_port_state_out_5_0_3;
  wire       [0:0]    mixColumns_port_state_out_5_0_4;
  wire       [0:0]    mixColumns_port_state_out_5_0_5;
  wire       [0:0]    mixColumns_port_state_out_5_0_6;
  wire       [0:0]    mixColumns_port_state_out_5_0_7;
  wire       [0:0]    mixColumns_port_state_out_5_1_0;
  wire       [0:0]    mixColumns_port_state_out_5_1_1;
  wire       [0:0]    mixColumns_port_state_out_5_1_2;
  wire       [0:0]    mixColumns_port_state_out_5_1_3;
  wire       [0:0]    mixColumns_port_state_out_5_1_4;
  wire       [0:0]    mixColumns_port_state_out_5_1_5;
  wire       [0:0]    mixColumns_port_state_out_5_1_6;
  wire       [0:0]    mixColumns_port_state_out_5_1_7;
  wire       [0:0]    mixColumns_port_state_out_5_2_0;
  wire       [0:0]    mixColumns_port_state_out_5_2_1;
  wire       [0:0]    mixColumns_port_state_out_5_2_2;
  wire       [0:0]    mixColumns_port_state_out_5_2_3;
  wire       [0:0]    mixColumns_port_state_out_5_2_4;
  wire       [0:0]    mixColumns_port_state_out_5_2_5;
  wire       [0:0]    mixColumns_port_state_out_5_2_6;
  wire       [0:0]    mixColumns_port_state_out_5_2_7;
  wire       [0:0]    mixColumns_port_state_out_5_3_0;
  wire       [0:0]    mixColumns_port_state_out_5_3_1;
  wire       [0:0]    mixColumns_port_state_out_5_3_2;
  wire       [0:0]    mixColumns_port_state_out_5_3_3;
  wire       [0:0]    mixColumns_port_state_out_5_3_4;
  wire       [0:0]    mixColumns_port_state_out_5_3_5;
  wire       [0:0]    mixColumns_port_state_out_5_3_6;
  wire       [0:0]    mixColumns_port_state_out_5_3_7;
  wire       [0:0]    mixColumns_port_state_out_6_0_0;
  wire       [0:0]    mixColumns_port_state_out_6_0_1;
  wire       [0:0]    mixColumns_port_state_out_6_0_2;
  wire       [0:0]    mixColumns_port_state_out_6_0_3;
  wire       [0:0]    mixColumns_port_state_out_6_0_4;
  wire       [0:0]    mixColumns_port_state_out_6_0_5;
  wire       [0:0]    mixColumns_port_state_out_6_0_6;
  wire       [0:0]    mixColumns_port_state_out_6_0_7;
  wire       [0:0]    mixColumns_port_state_out_6_1_0;
  wire       [0:0]    mixColumns_port_state_out_6_1_1;
  wire       [0:0]    mixColumns_port_state_out_6_1_2;
  wire       [0:0]    mixColumns_port_state_out_6_1_3;
  wire       [0:0]    mixColumns_port_state_out_6_1_4;
  wire       [0:0]    mixColumns_port_state_out_6_1_5;
  wire       [0:0]    mixColumns_port_state_out_6_1_6;
  wire       [0:0]    mixColumns_port_state_out_6_1_7;
  wire       [0:0]    mixColumns_port_state_out_6_2_0;
  wire       [0:0]    mixColumns_port_state_out_6_2_1;
  wire       [0:0]    mixColumns_port_state_out_6_2_2;
  wire       [0:0]    mixColumns_port_state_out_6_2_3;
  wire       [0:0]    mixColumns_port_state_out_6_2_4;
  wire       [0:0]    mixColumns_port_state_out_6_2_5;
  wire       [0:0]    mixColumns_port_state_out_6_2_6;
  wire       [0:0]    mixColumns_port_state_out_6_2_7;
  wire       [0:0]    mixColumns_port_state_out_6_3_0;
  wire       [0:0]    mixColumns_port_state_out_6_3_1;
  wire       [0:0]    mixColumns_port_state_out_6_3_2;
  wire       [0:0]    mixColumns_port_state_out_6_3_3;
  wire       [0:0]    mixColumns_port_state_out_6_3_4;
  wire       [0:0]    mixColumns_port_state_out_6_3_5;
  wire       [0:0]    mixColumns_port_state_out_6_3_6;
  wire       [0:0]    mixColumns_port_state_out_6_3_7;
  wire       [0:0]    mixColumns_port_state_out_7_0_0;
  wire       [0:0]    mixColumns_port_state_out_7_0_1;
  wire       [0:0]    mixColumns_port_state_out_7_0_2;
  wire       [0:0]    mixColumns_port_state_out_7_0_3;
  wire       [0:0]    mixColumns_port_state_out_7_0_4;
  wire       [0:0]    mixColumns_port_state_out_7_0_5;
  wire       [0:0]    mixColumns_port_state_out_7_0_6;
  wire       [0:0]    mixColumns_port_state_out_7_0_7;
  wire       [0:0]    mixColumns_port_state_out_7_1_0;
  wire       [0:0]    mixColumns_port_state_out_7_1_1;
  wire       [0:0]    mixColumns_port_state_out_7_1_2;
  wire       [0:0]    mixColumns_port_state_out_7_1_3;
  wire       [0:0]    mixColumns_port_state_out_7_1_4;
  wire       [0:0]    mixColumns_port_state_out_7_1_5;
  wire       [0:0]    mixColumns_port_state_out_7_1_6;
  wire       [0:0]    mixColumns_port_state_out_7_1_7;
  wire       [0:0]    mixColumns_port_state_out_7_2_0;
  wire       [0:0]    mixColumns_port_state_out_7_2_1;
  wire       [0:0]    mixColumns_port_state_out_7_2_2;
  wire       [0:0]    mixColumns_port_state_out_7_2_3;
  wire       [0:0]    mixColumns_port_state_out_7_2_4;
  wire       [0:0]    mixColumns_port_state_out_7_2_5;
  wire       [0:0]    mixColumns_port_state_out_7_2_6;
  wire       [0:0]    mixColumns_port_state_out_7_2_7;
  wire       [0:0]    mixColumns_port_state_out_7_3_0;
  wire       [0:0]    mixColumns_port_state_out_7_3_1;
  wire       [0:0]    mixColumns_port_state_out_7_3_2;
  wire       [0:0]    mixColumns_port_state_out_7_3_3;
  wire       [0:0]    mixColumns_port_state_out_7_3_4;
  wire       [0:0]    mixColumns_port_state_out_7_3_5;
  wire       [0:0]    mixColumns_port_state_out_7_3_6;
  wire       [0:0]    mixColumns_port_state_out_7_3_7;
  wire       [0:0]    mixColumns_port_state_out_8_0_0;
  wire       [0:0]    mixColumns_port_state_out_8_0_1;
  wire       [0:0]    mixColumns_port_state_out_8_0_2;
  wire       [0:0]    mixColumns_port_state_out_8_0_3;
  wire       [0:0]    mixColumns_port_state_out_8_0_4;
  wire       [0:0]    mixColumns_port_state_out_8_0_5;
  wire       [0:0]    mixColumns_port_state_out_8_0_6;
  wire       [0:0]    mixColumns_port_state_out_8_0_7;
  wire       [0:0]    mixColumns_port_state_out_8_1_0;
  wire       [0:0]    mixColumns_port_state_out_8_1_1;
  wire       [0:0]    mixColumns_port_state_out_8_1_2;
  wire       [0:0]    mixColumns_port_state_out_8_1_3;
  wire       [0:0]    mixColumns_port_state_out_8_1_4;
  wire       [0:0]    mixColumns_port_state_out_8_1_5;
  wire       [0:0]    mixColumns_port_state_out_8_1_6;
  wire       [0:0]    mixColumns_port_state_out_8_1_7;
  wire       [0:0]    mixColumns_port_state_out_8_2_0;
  wire       [0:0]    mixColumns_port_state_out_8_2_1;
  wire       [0:0]    mixColumns_port_state_out_8_2_2;
  wire       [0:0]    mixColumns_port_state_out_8_2_3;
  wire       [0:0]    mixColumns_port_state_out_8_2_4;
  wire       [0:0]    mixColumns_port_state_out_8_2_5;
  wire       [0:0]    mixColumns_port_state_out_8_2_6;
  wire       [0:0]    mixColumns_port_state_out_8_2_7;
  wire       [0:0]    mixColumns_port_state_out_8_3_0;
  wire       [0:0]    mixColumns_port_state_out_8_3_1;
  wire       [0:0]    mixColumns_port_state_out_8_3_2;
  wire       [0:0]    mixColumns_port_state_out_8_3_3;
  wire       [0:0]    mixColumns_port_state_out_8_3_4;
  wire       [0:0]    mixColumns_port_state_out_8_3_5;
  wire       [0:0]    mixColumns_port_state_out_8_3_6;
  wire       [0:0]    mixColumns_port_state_out_8_3_7;
  wire       [0:0]    mixColumns_port_state_out_9_0_0;
  wire       [0:0]    mixColumns_port_state_out_9_0_1;
  wire       [0:0]    mixColumns_port_state_out_9_0_2;
  wire       [0:0]    mixColumns_port_state_out_9_0_3;
  wire       [0:0]    mixColumns_port_state_out_9_0_4;
  wire       [0:0]    mixColumns_port_state_out_9_0_5;
  wire       [0:0]    mixColumns_port_state_out_9_0_6;
  wire       [0:0]    mixColumns_port_state_out_9_0_7;
  wire       [0:0]    mixColumns_port_state_out_9_1_0;
  wire       [0:0]    mixColumns_port_state_out_9_1_1;
  wire       [0:0]    mixColumns_port_state_out_9_1_2;
  wire       [0:0]    mixColumns_port_state_out_9_1_3;
  wire       [0:0]    mixColumns_port_state_out_9_1_4;
  wire       [0:0]    mixColumns_port_state_out_9_1_5;
  wire       [0:0]    mixColumns_port_state_out_9_1_6;
  wire       [0:0]    mixColumns_port_state_out_9_1_7;
  wire       [0:0]    mixColumns_port_state_out_9_2_0;
  wire       [0:0]    mixColumns_port_state_out_9_2_1;
  wire       [0:0]    mixColumns_port_state_out_9_2_2;
  wire       [0:0]    mixColumns_port_state_out_9_2_3;
  wire       [0:0]    mixColumns_port_state_out_9_2_4;
  wire       [0:0]    mixColumns_port_state_out_9_2_5;
  wire       [0:0]    mixColumns_port_state_out_9_2_6;
  wire       [0:0]    mixColumns_port_state_out_9_2_7;
  wire       [0:0]    mixColumns_port_state_out_9_3_0;
  wire       [0:0]    mixColumns_port_state_out_9_3_1;
  wire       [0:0]    mixColumns_port_state_out_9_3_2;
  wire       [0:0]    mixColumns_port_state_out_9_3_3;
  wire       [0:0]    mixColumns_port_state_out_9_3_4;
  wire       [0:0]    mixColumns_port_state_out_9_3_5;
  wire       [0:0]    mixColumns_port_state_out_9_3_6;
  wire       [0:0]    mixColumns_port_state_out_9_3_7;
  wire       [0:0]    mixColumns_port_state_out_10_0_0;
  wire       [0:0]    mixColumns_port_state_out_10_0_1;
  wire       [0:0]    mixColumns_port_state_out_10_0_2;
  wire       [0:0]    mixColumns_port_state_out_10_0_3;
  wire       [0:0]    mixColumns_port_state_out_10_0_4;
  wire       [0:0]    mixColumns_port_state_out_10_0_5;
  wire       [0:0]    mixColumns_port_state_out_10_0_6;
  wire       [0:0]    mixColumns_port_state_out_10_0_7;
  wire       [0:0]    mixColumns_port_state_out_10_1_0;
  wire       [0:0]    mixColumns_port_state_out_10_1_1;
  wire       [0:0]    mixColumns_port_state_out_10_1_2;
  wire       [0:0]    mixColumns_port_state_out_10_1_3;
  wire       [0:0]    mixColumns_port_state_out_10_1_4;
  wire       [0:0]    mixColumns_port_state_out_10_1_5;
  wire       [0:0]    mixColumns_port_state_out_10_1_6;
  wire       [0:0]    mixColumns_port_state_out_10_1_7;
  wire       [0:0]    mixColumns_port_state_out_10_2_0;
  wire       [0:0]    mixColumns_port_state_out_10_2_1;
  wire       [0:0]    mixColumns_port_state_out_10_2_2;
  wire       [0:0]    mixColumns_port_state_out_10_2_3;
  wire       [0:0]    mixColumns_port_state_out_10_2_4;
  wire       [0:0]    mixColumns_port_state_out_10_2_5;
  wire       [0:0]    mixColumns_port_state_out_10_2_6;
  wire       [0:0]    mixColumns_port_state_out_10_2_7;
  wire       [0:0]    mixColumns_port_state_out_10_3_0;
  wire       [0:0]    mixColumns_port_state_out_10_3_1;
  wire       [0:0]    mixColumns_port_state_out_10_3_2;
  wire       [0:0]    mixColumns_port_state_out_10_3_3;
  wire       [0:0]    mixColumns_port_state_out_10_3_4;
  wire       [0:0]    mixColumns_port_state_out_10_3_5;
  wire       [0:0]    mixColumns_port_state_out_10_3_6;
  wire       [0:0]    mixColumns_port_state_out_10_3_7;
  wire       [0:0]    mixColumns_port_state_out_11_0_0;
  wire       [0:0]    mixColumns_port_state_out_11_0_1;
  wire       [0:0]    mixColumns_port_state_out_11_0_2;
  wire       [0:0]    mixColumns_port_state_out_11_0_3;
  wire       [0:0]    mixColumns_port_state_out_11_0_4;
  wire       [0:0]    mixColumns_port_state_out_11_0_5;
  wire       [0:0]    mixColumns_port_state_out_11_0_6;
  wire       [0:0]    mixColumns_port_state_out_11_0_7;
  wire       [0:0]    mixColumns_port_state_out_11_1_0;
  wire       [0:0]    mixColumns_port_state_out_11_1_1;
  wire       [0:0]    mixColumns_port_state_out_11_1_2;
  wire       [0:0]    mixColumns_port_state_out_11_1_3;
  wire       [0:0]    mixColumns_port_state_out_11_1_4;
  wire       [0:0]    mixColumns_port_state_out_11_1_5;
  wire       [0:0]    mixColumns_port_state_out_11_1_6;
  wire       [0:0]    mixColumns_port_state_out_11_1_7;
  wire       [0:0]    mixColumns_port_state_out_11_2_0;
  wire       [0:0]    mixColumns_port_state_out_11_2_1;
  wire       [0:0]    mixColumns_port_state_out_11_2_2;
  wire       [0:0]    mixColumns_port_state_out_11_2_3;
  wire       [0:0]    mixColumns_port_state_out_11_2_4;
  wire       [0:0]    mixColumns_port_state_out_11_2_5;
  wire       [0:0]    mixColumns_port_state_out_11_2_6;
  wire       [0:0]    mixColumns_port_state_out_11_2_7;
  wire       [0:0]    mixColumns_port_state_out_11_3_0;
  wire       [0:0]    mixColumns_port_state_out_11_3_1;
  wire       [0:0]    mixColumns_port_state_out_11_3_2;
  wire       [0:0]    mixColumns_port_state_out_11_3_3;
  wire       [0:0]    mixColumns_port_state_out_11_3_4;
  wire       [0:0]    mixColumns_port_state_out_11_3_5;
  wire       [0:0]    mixColumns_port_state_out_11_3_6;
  wire       [0:0]    mixColumns_port_state_out_11_3_7;
  wire       [0:0]    mixColumns_port_state_out_12_0_0;
  wire       [0:0]    mixColumns_port_state_out_12_0_1;
  wire       [0:0]    mixColumns_port_state_out_12_0_2;
  wire       [0:0]    mixColumns_port_state_out_12_0_3;
  wire       [0:0]    mixColumns_port_state_out_12_0_4;
  wire       [0:0]    mixColumns_port_state_out_12_0_5;
  wire       [0:0]    mixColumns_port_state_out_12_0_6;
  wire       [0:0]    mixColumns_port_state_out_12_0_7;
  wire       [0:0]    mixColumns_port_state_out_12_1_0;
  wire       [0:0]    mixColumns_port_state_out_12_1_1;
  wire       [0:0]    mixColumns_port_state_out_12_1_2;
  wire       [0:0]    mixColumns_port_state_out_12_1_3;
  wire       [0:0]    mixColumns_port_state_out_12_1_4;
  wire       [0:0]    mixColumns_port_state_out_12_1_5;
  wire       [0:0]    mixColumns_port_state_out_12_1_6;
  wire       [0:0]    mixColumns_port_state_out_12_1_7;
  wire       [0:0]    mixColumns_port_state_out_12_2_0;
  wire       [0:0]    mixColumns_port_state_out_12_2_1;
  wire       [0:0]    mixColumns_port_state_out_12_2_2;
  wire       [0:0]    mixColumns_port_state_out_12_2_3;
  wire       [0:0]    mixColumns_port_state_out_12_2_4;
  wire       [0:0]    mixColumns_port_state_out_12_2_5;
  wire       [0:0]    mixColumns_port_state_out_12_2_6;
  wire       [0:0]    mixColumns_port_state_out_12_2_7;
  wire       [0:0]    mixColumns_port_state_out_12_3_0;
  wire       [0:0]    mixColumns_port_state_out_12_3_1;
  wire       [0:0]    mixColumns_port_state_out_12_3_2;
  wire       [0:0]    mixColumns_port_state_out_12_3_3;
  wire       [0:0]    mixColumns_port_state_out_12_3_4;
  wire       [0:0]    mixColumns_port_state_out_12_3_5;
  wire       [0:0]    mixColumns_port_state_out_12_3_6;
  wire       [0:0]    mixColumns_port_state_out_12_3_7;
  wire       [0:0]    mixColumns_port_state_out_13_0_0;
  wire       [0:0]    mixColumns_port_state_out_13_0_1;
  wire       [0:0]    mixColumns_port_state_out_13_0_2;
  wire       [0:0]    mixColumns_port_state_out_13_0_3;
  wire       [0:0]    mixColumns_port_state_out_13_0_4;
  wire       [0:0]    mixColumns_port_state_out_13_0_5;
  wire       [0:0]    mixColumns_port_state_out_13_0_6;
  wire       [0:0]    mixColumns_port_state_out_13_0_7;
  wire       [0:0]    mixColumns_port_state_out_13_1_0;
  wire       [0:0]    mixColumns_port_state_out_13_1_1;
  wire       [0:0]    mixColumns_port_state_out_13_1_2;
  wire       [0:0]    mixColumns_port_state_out_13_1_3;
  wire       [0:0]    mixColumns_port_state_out_13_1_4;
  wire       [0:0]    mixColumns_port_state_out_13_1_5;
  wire       [0:0]    mixColumns_port_state_out_13_1_6;
  wire       [0:0]    mixColumns_port_state_out_13_1_7;
  wire       [0:0]    mixColumns_port_state_out_13_2_0;
  wire       [0:0]    mixColumns_port_state_out_13_2_1;
  wire       [0:0]    mixColumns_port_state_out_13_2_2;
  wire       [0:0]    mixColumns_port_state_out_13_2_3;
  wire       [0:0]    mixColumns_port_state_out_13_2_4;
  wire       [0:0]    mixColumns_port_state_out_13_2_5;
  wire       [0:0]    mixColumns_port_state_out_13_2_6;
  wire       [0:0]    mixColumns_port_state_out_13_2_7;
  wire       [0:0]    mixColumns_port_state_out_13_3_0;
  wire       [0:0]    mixColumns_port_state_out_13_3_1;
  wire       [0:0]    mixColumns_port_state_out_13_3_2;
  wire       [0:0]    mixColumns_port_state_out_13_3_3;
  wire       [0:0]    mixColumns_port_state_out_13_3_4;
  wire       [0:0]    mixColumns_port_state_out_13_3_5;
  wire       [0:0]    mixColumns_port_state_out_13_3_6;
  wire       [0:0]    mixColumns_port_state_out_13_3_7;
  wire       [0:0]    mixColumns_port_state_out_14_0_0;
  wire       [0:0]    mixColumns_port_state_out_14_0_1;
  wire       [0:0]    mixColumns_port_state_out_14_0_2;
  wire       [0:0]    mixColumns_port_state_out_14_0_3;
  wire       [0:0]    mixColumns_port_state_out_14_0_4;
  wire       [0:0]    mixColumns_port_state_out_14_0_5;
  wire       [0:0]    mixColumns_port_state_out_14_0_6;
  wire       [0:0]    mixColumns_port_state_out_14_0_7;
  wire       [0:0]    mixColumns_port_state_out_14_1_0;
  wire       [0:0]    mixColumns_port_state_out_14_1_1;
  wire       [0:0]    mixColumns_port_state_out_14_1_2;
  wire       [0:0]    mixColumns_port_state_out_14_1_3;
  wire       [0:0]    mixColumns_port_state_out_14_1_4;
  wire       [0:0]    mixColumns_port_state_out_14_1_5;
  wire       [0:0]    mixColumns_port_state_out_14_1_6;
  wire       [0:0]    mixColumns_port_state_out_14_1_7;
  wire       [0:0]    mixColumns_port_state_out_14_2_0;
  wire       [0:0]    mixColumns_port_state_out_14_2_1;
  wire       [0:0]    mixColumns_port_state_out_14_2_2;
  wire       [0:0]    mixColumns_port_state_out_14_2_3;
  wire       [0:0]    mixColumns_port_state_out_14_2_4;
  wire       [0:0]    mixColumns_port_state_out_14_2_5;
  wire       [0:0]    mixColumns_port_state_out_14_2_6;
  wire       [0:0]    mixColumns_port_state_out_14_2_7;
  wire       [0:0]    mixColumns_port_state_out_14_3_0;
  wire       [0:0]    mixColumns_port_state_out_14_3_1;
  wire       [0:0]    mixColumns_port_state_out_14_3_2;
  wire       [0:0]    mixColumns_port_state_out_14_3_3;
  wire       [0:0]    mixColumns_port_state_out_14_3_4;
  wire       [0:0]    mixColumns_port_state_out_14_3_5;
  wire       [0:0]    mixColumns_port_state_out_14_3_6;
  wire       [0:0]    mixColumns_port_state_out_14_3_7;
  wire       [0:0]    mixColumns_port_state_out_15_0_0;
  wire       [0:0]    mixColumns_port_state_out_15_0_1;
  wire       [0:0]    mixColumns_port_state_out_15_0_2;
  wire       [0:0]    mixColumns_port_state_out_15_0_3;
  wire       [0:0]    mixColumns_port_state_out_15_0_4;
  wire       [0:0]    mixColumns_port_state_out_15_0_5;
  wire       [0:0]    mixColumns_port_state_out_15_0_6;
  wire       [0:0]    mixColumns_port_state_out_15_0_7;
  wire       [0:0]    mixColumns_port_state_out_15_1_0;
  wire       [0:0]    mixColumns_port_state_out_15_1_1;
  wire       [0:0]    mixColumns_port_state_out_15_1_2;
  wire       [0:0]    mixColumns_port_state_out_15_1_3;
  wire       [0:0]    mixColumns_port_state_out_15_1_4;
  wire       [0:0]    mixColumns_port_state_out_15_1_5;
  wire       [0:0]    mixColumns_port_state_out_15_1_6;
  wire       [0:0]    mixColumns_port_state_out_15_1_7;
  wire       [0:0]    mixColumns_port_state_out_15_2_0;
  wire       [0:0]    mixColumns_port_state_out_15_2_1;
  wire       [0:0]    mixColumns_port_state_out_15_2_2;
  wire       [0:0]    mixColumns_port_state_out_15_2_3;
  wire       [0:0]    mixColumns_port_state_out_15_2_4;
  wire       [0:0]    mixColumns_port_state_out_15_2_5;
  wire       [0:0]    mixColumns_port_state_out_15_2_6;
  wire       [0:0]    mixColumns_port_state_out_15_2_7;
  wire       [0:0]    mixColumns_port_state_out_15_3_0;
  wire       [0:0]    mixColumns_port_state_out_15_3_1;
  wire       [0:0]    mixColumns_port_state_out_15_3_2;
  wire       [0:0]    mixColumns_port_state_out_15_3_3;
  wire       [0:0]    mixColumns_port_state_out_15_3_4;
  wire       [0:0]    mixColumns_port_state_out_15_3_5;
  wire       [0:0]    mixColumns_port_state_out_15_3_6;
  wire       [0:0]    mixColumns_port_state_out_15_3_7;
  wire       [0:0]    subBytes_out_0_0_0;
  wire       [0:0]    subBytes_out_0_0_1;
  wire       [0:0]    subBytes_out_0_0_2;
  wire       [0:0]    subBytes_out_0_0_3;
  wire       [0:0]    subBytes_out_0_0_4;
  wire       [0:0]    subBytes_out_0_0_5;
  wire       [0:0]    subBytes_out_0_0_6;
  wire       [0:0]    subBytes_out_0_0_7;
  wire       [0:0]    subBytes_out_0_1_0;
  wire       [0:0]    subBytes_out_0_1_1;
  wire       [0:0]    subBytes_out_0_1_2;
  wire       [0:0]    subBytes_out_0_1_3;
  wire       [0:0]    subBytes_out_0_1_4;
  wire       [0:0]    subBytes_out_0_1_5;
  wire       [0:0]    subBytes_out_0_1_6;
  wire       [0:0]    subBytes_out_0_1_7;
  wire       [0:0]    subBytes_out_0_2_0;
  wire       [0:0]    subBytes_out_0_2_1;
  wire       [0:0]    subBytes_out_0_2_2;
  wire       [0:0]    subBytes_out_0_2_3;
  wire       [0:0]    subBytes_out_0_2_4;
  wire       [0:0]    subBytes_out_0_2_5;
  wire       [0:0]    subBytes_out_0_2_6;
  wire       [0:0]    subBytes_out_0_2_7;
  wire       [0:0]    subBytes_out_0_3_0;
  wire       [0:0]    subBytes_out_0_3_1;
  wire       [0:0]    subBytes_out_0_3_2;
  wire       [0:0]    subBytes_out_0_3_3;
  wire       [0:0]    subBytes_out_0_3_4;
  wire       [0:0]    subBytes_out_0_3_5;
  wire       [0:0]    subBytes_out_0_3_6;
  wire       [0:0]    subBytes_out_0_3_7;
  wire       [0:0]    subBytes_out_1_0_0;
  wire       [0:0]    subBytes_out_1_0_1;
  wire       [0:0]    subBytes_out_1_0_2;
  wire       [0:0]    subBytes_out_1_0_3;
  wire       [0:0]    subBytes_out_1_0_4;
  wire       [0:0]    subBytes_out_1_0_5;
  wire       [0:0]    subBytes_out_1_0_6;
  wire       [0:0]    subBytes_out_1_0_7;
  wire       [0:0]    subBytes_out_1_1_0;
  wire       [0:0]    subBytes_out_1_1_1;
  wire       [0:0]    subBytes_out_1_1_2;
  wire       [0:0]    subBytes_out_1_1_3;
  wire       [0:0]    subBytes_out_1_1_4;
  wire       [0:0]    subBytes_out_1_1_5;
  wire       [0:0]    subBytes_out_1_1_6;
  wire       [0:0]    subBytes_out_1_1_7;
  wire       [0:0]    subBytes_out_1_2_0;
  wire       [0:0]    subBytes_out_1_2_1;
  wire       [0:0]    subBytes_out_1_2_2;
  wire       [0:0]    subBytes_out_1_2_3;
  wire       [0:0]    subBytes_out_1_2_4;
  wire       [0:0]    subBytes_out_1_2_5;
  wire       [0:0]    subBytes_out_1_2_6;
  wire       [0:0]    subBytes_out_1_2_7;
  wire       [0:0]    subBytes_out_1_3_0;
  wire       [0:0]    subBytes_out_1_3_1;
  wire       [0:0]    subBytes_out_1_3_2;
  wire       [0:0]    subBytes_out_1_3_3;
  wire       [0:0]    subBytes_out_1_3_4;
  wire       [0:0]    subBytes_out_1_3_5;
  wire       [0:0]    subBytes_out_1_3_6;
  wire       [0:0]    subBytes_out_1_3_7;
  wire       [0:0]    subBytes_out_2_0_0;
  wire       [0:0]    subBytes_out_2_0_1;
  wire       [0:0]    subBytes_out_2_0_2;
  wire       [0:0]    subBytes_out_2_0_3;
  wire       [0:0]    subBytes_out_2_0_4;
  wire       [0:0]    subBytes_out_2_0_5;
  wire       [0:0]    subBytes_out_2_0_6;
  wire       [0:0]    subBytes_out_2_0_7;
  wire       [0:0]    subBytes_out_2_1_0;
  wire       [0:0]    subBytes_out_2_1_1;
  wire       [0:0]    subBytes_out_2_1_2;
  wire       [0:0]    subBytes_out_2_1_3;
  wire       [0:0]    subBytes_out_2_1_4;
  wire       [0:0]    subBytes_out_2_1_5;
  wire       [0:0]    subBytes_out_2_1_6;
  wire       [0:0]    subBytes_out_2_1_7;
  wire       [0:0]    subBytes_out_2_2_0;
  wire       [0:0]    subBytes_out_2_2_1;
  wire       [0:0]    subBytes_out_2_2_2;
  wire       [0:0]    subBytes_out_2_2_3;
  wire       [0:0]    subBytes_out_2_2_4;
  wire       [0:0]    subBytes_out_2_2_5;
  wire       [0:0]    subBytes_out_2_2_6;
  wire       [0:0]    subBytes_out_2_2_7;
  wire       [0:0]    subBytes_out_2_3_0;
  wire       [0:0]    subBytes_out_2_3_1;
  wire       [0:0]    subBytes_out_2_3_2;
  wire       [0:0]    subBytes_out_2_3_3;
  wire       [0:0]    subBytes_out_2_3_4;
  wire       [0:0]    subBytes_out_2_3_5;
  wire       [0:0]    subBytes_out_2_3_6;
  wire       [0:0]    subBytes_out_2_3_7;
  wire       [0:0]    subBytes_out_3_0_0;
  wire       [0:0]    subBytes_out_3_0_1;
  wire       [0:0]    subBytes_out_3_0_2;
  wire       [0:0]    subBytes_out_3_0_3;
  wire       [0:0]    subBytes_out_3_0_4;
  wire       [0:0]    subBytes_out_3_0_5;
  wire       [0:0]    subBytes_out_3_0_6;
  wire       [0:0]    subBytes_out_3_0_7;
  wire       [0:0]    subBytes_out_3_1_0;
  wire       [0:0]    subBytes_out_3_1_1;
  wire       [0:0]    subBytes_out_3_1_2;
  wire       [0:0]    subBytes_out_3_1_3;
  wire       [0:0]    subBytes_out_3_1_4;
  wire       [0:0]    subBytes_out_3_1_5;
  wire       [0:0]    subBytes_out_3_1_6;
  wire       [0:0]    subBytes_out_3_1_7;
  wire       [0:0]    subBytes_out_3_2_0;
  wire       [0:0]    subBytes_out_3_2_1;
  wire       [0:0]    subBytes_out_3_2_2;
  wire       [0:0]    subBytes_out_3_2_3;
  wire       [0:0]    subBytes_out_3_2_4;
  wire       [0:0]    subBytes_out_3_2_5;
  wire       [0:0]    subBytes_out_3_2_6;
  wire       [0:0]    subBytes_out_3_2_7;
  wire       [0:0]    subBytes_out_3_3_0;
  wire       [0:0]    subBytes_out_3_3_1;
  wire       [0:0]    subBytes_out_3_3_2;
  wire       [0:0]    subBytes_out_3_3_3;
  wire       [0:0]    subBytes_out_3_3_4;
  wire       [0:0]    subBytes_out_3_3_5;
  wire       [0:0]    subBytes_out_3_3_6;
  wire       [0:0]    subBytes_out_3_3_7;
  wire       [0:0]    subBytes_out_4_0_0;
  wire       [0:0]    subBytes_out_4_0_1;
  wire       [0:0]    subBytes_out_4_0_2;
  wire       [0:0]    subBytes_out_4_0_3;
  wire       [0:0]    subBytes_out_4_0_4;
  wire       [0:0]    subBytes_out_4_0_5;
  wire       [0:0]    subBytes_out_4_0_6;
  wire       [0:0]    subBytes_out_4_0_7;
  wire       [0:0]    subBytes_out_4_1_0;
  wire       [0:0]    subBytes_out_4_1_1;
  wire       [0:0]    subBytes_out_4_1_2;
  wire       [0:0]    subBytes_out_4_1_3;
  wire       [0:0]    subBytes_out_4_1_4;
  wire       [0:0]    subBytes_out_4_1_5;
  wire       [0:0]    subBytes_out_4_1_6;
  wire       [0:0]    subBytes_out_4_1_7;
  wire       [0:0]    subBytes_out_4_2_0;
  wire       [0:0]    subBytes_out_4_2_1;
  wire       [0:0]    subBytes_out_4_2_2;
  wire       [0:0]    subBytes_out_4_2_3;
  wire       [0:0]    subBytes_out_4_2_4;
  wire       [0:0]    subBytes_out_4_2_5;
  wire       [0:0]    subBytes_out_4_2_6;
  wire       [0:0]    subBytes_out_4_2_7;
  wire       [0:0]    subBytes_out_4_3_0;
  wire       [0:0]    subBytes_out_4_3_1;
  wire       [0:0]    subBytes_out_4_3_2;
  wire       [0:0]    subBytes_out_4_3_3;
  wire       [0:0]    subBytes_out_4_3_4;
  wire       [0:0]    subBytes_out_4_3_5;
  wire       [0:0]    subBytes_out_4_3_6;
  wire       [0:0]    subBytes_out_4_3_7;
  wire       [0:0]    subBytes_out_5_0_0;
  wire       [0:0]    subBytes_out_5_0_1;
  wire       [0:0]    subBytes_out_5_0_2;
  wire       [0:0]    subBytes_out_5_0_3;
  wire       [0:0]    subBytes_out_5_0_4;
  wire       [0:0]    subBytes_out_5_0_5;
  wire       [0:0]    subBytes_out_5_0_6;
  wire       [0:0]    subBytes_out_5_0_7;
  wire       [0:0]    subBytes_out_5_1_0;
  wire       [0:0]    subBytes_out_5_1_1;
  wire       [0:0]    subBytes_out_5_1_2;
  wire       [0:0]    subBytes_out_5_1_3;
  wire       [0:0]    subBytes_out_5_1_4;
  wire       [0:0]    subBytes_out_5_1_5;
  wire       [0:0]    subBytes_out_5_1_6;
  wire       [0:0]    subBytes_out_5_1_7;
  wire       [0:0]    subBytes_out_5_2_0;
  wire       [0:0]    subBytes_out_5_2_1;
  wire       [0:0]    subBytes_out_5_2_2;
  wire       [0:0]    subBytes_out_5_2_3;
  wire       [0:0]    subBytes_out_5_2_4;
  wire       [0:0]    subBytes_out_5_2_5;
  wire       [0:0]    subBytes_out_5_2_6;
  wire       [0:0]    subBytes_out_5_2_7;
  wire       [0:0]    subBytes_out_5_3_0;
  wire       [0:0]    subBytes_out_5_3_1;
  wire       [0:0]    subBytes_out_5_3_2;
  wire       [0:0]    subBytes_out_5_3_3;
  wire       [0:0]    subBytes_out_5_3_4;
  wire       [0:0]    subBytes_out_5_3_5;
  wire       [0:0]    subBytes_out_5_3_6;
  wire       [0:0]    subBytes_out_5_3_7;
  wire       [0:0]    subBytes_out_6_0_0;
  wire       [0:0]    subBytes_out_6_0_1;
  wire       [0:0]    subBytes_out_6_0_2;
  wire       [0:0]    subBytes_out_6_0_3;
  wire       [0:0]    subBytes_out_6_0_4;
  wire       [0:0]    subBytes_out_6_0_5;
  wire       [0:0]    subBytes_out_6_0_6;
  wire       [0:0]    subBytes_out_6_0_7;
  wire       [0:0]    subBytes_out_6_1_0;
  wire       [0:0]    subBytes_out_6_1_1;
  wire       [0:0]    subBytes_out_6_1_2;
  wire       [0:0]    subBytes_out_6_1_3;
  wire       [0:0]    subBytes_out_6_1_4;
  wire       [0:0]    subBytes_out_6_1_5;
  wire       [0:0]    subBytes_out_6_1_6;
  wire       [0:0]    subBytes_out_6_1_7;
  wire       [0:0]    subBytes_out_6_2_0;
  wire       [0:0]    subBytes_out_6_2_1;
  wire       [0:0]    subBytes_out_6_2_2;
  wire       [0:0]    subBytes_out_6_2_3;
  wire       [0:0]    subBytes_out_6_2_4;
  wire       [0:0]    subBytes_out_6_2_5;
  wire       [0:0]    subBytes_out_6_2_6;
  wire       [0:0]    subBytes_out_6_2_7;
  wire       [0:0]    subBytes_out_6_3_0;
  wire       [0:0]    subBytes_out_6_3_1;
  wire       [0:0]    subBytes_out_6_3_2;
  wire       [0:0]    subBytes_out_6_3_3;
  wire       [0:0]    subBytes_out_6_3_4;
  wire       [0:0]    subBytes_out_6_3_5;
  wire       [0:0]    subBytes_out_6_3_6;
  wire       [0:0]    subBytes_out_6_3_7;
  wire       [0:0]    subBytes_out_7_0_0;
  wire       [0:0]    subBytes_out_7_0_1;
  wire       [0:0]    subBytes_out_7_0_2;
  wire       [0:0]    subBytes_out_7_0_3;
  wire       [0:0]    subBytes_out_7_0_4;
  wire       [0:0]    subBytes_out_7_0_5;
  wire       [0:0]    subBytes_out_7_0_6;
  wire       [0:0]    subBytes_out_7_0_7;
  wire       [0:0]    subBytes_out_7_1_0;
  wire       [0:0]    subBytes_out_7_1_1;
  wire       [0:0]    subBytes_out_7_1_2;
  wire       [0:0]    subBytes_out_7_1_3;
  wire       [0:0]    subBytes_out_7_1_4;
  wire       [0:0]    subBytes_out_7_1_5;
  wire       [0:0]    subBytes_out_7_1_6;
  wire       [0:0]    subBytes_out_7_1_7;
  wire       [0:0]    subBytes_out_7_2_0;
  wire       [0:0]    subBytes_out_7_2_1;
  wire       [0:0]    subBytes_out_7_2_2;
  wire       [0:0]    subBytes_out_7_2_3;
  wire       [0:0]    subBytes_out_7_2_4;
  wire       [0:0]    subBytes_out_7_2_5;
  wire       [0:0]    subBytes_out_7_2_6;
  wire       [0:0]    subBytes_out_7_2_7;
  wire       [0:0]    subBytes_out_7_3_0;
  wire       [0:0]    subBytes_out_7_3_1;
  wire       [0:0]    subBytes_out_7_3_2;
  wire       [0:0]    subBytes_out_7_3_3;
  wire       [0:0]    subBytes_out_7_3_4;
  wire       [0:0]    subBytes_out_7_3_5;
  wire       [0:0]    subBytes_out_7_3_6;
  wire       [0:0]    subBytes_out_7_3_7;
  wire       [0:0]    subBytes_out_8_0_0;
  wire       [0:0]    subBytes_out_8_0_1;
  wire       [0:0]    subBytes_out_8_0_2;
  wire       [0:0]    subBytes_out_8_0_3;
  wire       [0:0]    subBytes_out_8_0_4;
  wire       [0:0]    subBytes_out_8_0_5;
  wire       [0:0]    subBytes_out_8_0_6;
  wire       [0:0]    subBytes_out_8_0_7;
  wire       [0:0]    subBytes_out_8_1_0;
  wire       [0:0]    subBytes_out_8_1_1;
  wire       [0:0]    subBytes_out_8_1_2;
  wire       [0:0]    subBytes_out_8_1_3;
  wire       [0:0]    subBytes_out_8_1_4;
  wire       [0:0]    subBytes_out_8_1_5;
  wire       [0:0]    subBytes_out_8_1_6;
  wire       [0:0]    subBytes_out_8_1_7;
  wire       [0:0]    subBytes_out_8_2_0;
  wire       [0:0]    subBytes_out_8_2_1;
  wire       [0:0]    subBytes_out_8_2_2;
  wire       [0:0]    subBytes_out_8_2_3;
  wire       [0:0]    subBytes_out_8_2_4;
  wire       [0:0]    subBytes_out_8_2_5;
  wire       [0:0]    subBytes_out_8_2_6;
  wire       [0:0]    subBytes_out_8_2_7;
  wire       [0:0]    subBytes_out_8_3_0;
  wire       [0:0]    subBytes_out_8_3_1;
  wire       [0:0]    subBytes_out_8_3_2;
  wire       [0:0]    subBytes_out_8_3_3;
  wire       [0:0]    subBytes_out_8_3_4;
  wire       [0:0]    subBytes_out_8_3_5;
  wire       [0:0]    subBytes_out_8_3_6;
  wire       [0:0]    subBytes_out_8_3_7;
  wire       [0:0]    subBytes_out_9_0_0;
  wire       [0:0]    subBytes_out_9_0_1;
  wire       [0:0]    subBytes_out_9_0_2;
  wire       [0:0]    subBytes_out_9_0_3;
  wire       [0:0]    subBytes_out_9_0_4;
  wire       [0:0]    subBytes_out_9_0_5;
  wire       [0:0]    subBytes_out_9_0_6;
  wire       [0:0]    subBytes_out_9_0_7;
  wire       [0:0]    subBytes_out_9_1_0;
  wire       [0:0]    subBytes_out_9_1_1;
  wire       [0:0]    subBytes_out_9_1_2;
  wire       [0:0]    subBytes_out_9_1_3;
  wire       [0:0]    subBytes_out_9_1_4;
  wire       [0:0]    subBytes_out_9_1_5;
  wire       [0:0]    subBytes_out_9_1_6;
  wire       [0:0]    subBytes_out_9_1_7;
  wire       [0:0]    subBytes_out_9_2_0;
  wire       [0:0]    subBytes_out_9_2_1;
  wire       [0:0]    subBytes_out_9_2_2;
  wire       [0:0]    subBytes_out_9_2_3;
  wire       [0:0]    subBytes_out_9_2_4;
  wire       [0:0]    subBytes_out_9_2_5;
  wire       [0:0]    subBytes_out_9_2_6;
  wire       [0:0]    subBytes_out_9_2_7;
  wire       [0:0]    subBytes_out_9_3_0;
  wire       [0:0]    subBytes_out_9_3_1;
  wire       [0:0]    subBytes_out_9_3_2;
  wire       [0:0]    subBytes_out_9_3_3;
  wire       [0:0]    subBytes_out_9_3_4;
  wire       [0:0]    subBytes_out_9_3_5;
  wire       [0:0]    subBytes_out_9_3_6;
  wire       [0:0]    subBytes_out_9_3_7;
  wire       [0:0]    subBytes_out_10_0_0;
  wire       [0:0]    subBytes_out_10_0_1;
  wire       [0:0]    subBytes_out_10_0_2;
  wire       [0:0]    subBytes_out_10_0_3;
  wire       [0:0]    subBytes_out_10_0_4;
  wire       [0:0]    subBytes_out_10_0_5;
  wire       [0:0]    subBytes_out_10_0_6;
  wire       [0:0]    subBytes_out_10_0_7;
  wire       [0:0]    subBytes_out_10_1_0;
  wire       [0:0]    subBytes_out_10_1_1;
  wire       [0:0]    subBytes_out_10_1_2;
  wire       [0:0]    subBytes_out_10_1_3;
  wire       [0:0]    subBytes_out_10_1_4;
  wire       [0:0]    subBytes_out_10_1_5;
  wire       [0:0]    subBytes_out_10_1_6;
  wire       [0:0]    subBytes_out_10_1_7;
  wire       [0:0]    subBytes_out_10_2_0;
  wire       [0:0]    subBytes_out_10_2_1;
  wire       [0:0]    subBytes_out_10_2_2;
  wire       [0:0]    subBytes_out_10_2_3;
  wire       [0:0]    subBytes_out_10_2_4;
  wire       [0:0]    subBytes_out_10_2_5;
  wire       [0:0]    subBytes_out_10_2_6;
  wire       [0:0]    subBytes_out_10_2_7;
  wire       [0:0]    subBytes_out_10_3_0;
  wire       [0:0]    subBytes_out_10_3_1;
  wire       [0:0]    subBytes_out_10_3_2;
  wire       [0:0]    subBytes_out_10_3_3;
  wire       [0:0]    subBytes_out_10_3_4;
  wire       [0:0]    subBytes_out_10_3_5;
  wire       [0:0]    subBytes_out_10_3_6;
  wire       [0:0]    subBytes_out_10_3_7;
  wire       [0:0]    subBytes_out_11_0_0;
  wire       [0:0]    subBytes_out_11_0_1;
  wire       [0:0]    subBytes_out_11_0_2;
  wire       [0:0]    subBytes_out_11_0_3;
  wire       [0:0]    subBytes_out_11_0_4;
  wire       [0:0]    subBytes_out_11_0_5;
  wire       [0:0]    subBytes_out_11_0_6;
  wire       [0:0]    subBytes_out_11_0_7;
  wire       [0:0]    subBytes_out_11_1_0;
  wire       [0:0]    subBytes_out_11_1_1;
  wire       [0:0]    subBytes_out_11_1_2;
  wire       [0:0]    subBytes_out_11_1_3;
  wire       [0:0]    subBytes_out_11_1_4;
  wire       [0:0]    subBytes_out_11_1_5;
  wire       [0:0]    subBytes_out_11_1_6;
  wire       [0:0]    subBytes_out_11_1_7;
  wire       [0:0]    subBytes_out_11_2_0;
  wire       [0:0]    subBytes_out_11_2_1;
  wire       [0:0]    subBytes_out_11_2_2;
  wire       [0:0]    subBytes_out_11_2_3;
  wire       [0:0]    subBytes_out_11_2_4;
  wire       [0:0]    subBytes_out_11_2_5;
  wire       [0:0]    subBytes_out_11_2_6;
  wire       [0:0]    subBytes_out_11_2_7;
  wire       [0:0]    subBytes_out_11_3_0;
  wire       [0:0]    subBytes_out_11_3_1;
  wire       [0:0]    subBytes_out_11_3_2;
  wire       [0:0]    subBytes_out_11_3_3;
  wire       [0:0]    subBytes_out_11_3_4;
  wire       [0:0]    subBytes_out_11_3_5;
  wire       [0:0]    subBytes_out_11_3_6;
  wire       [0:0]    subBytes_out_11_3_7;
  wire       [0:0]    subBytes_out_12_0_0;
  wire       [0:0]    subBytes_out_12_0_1;
  wire       [0:0]    subBytes_out_12_0_2;
  wire       [0:0]    subBytes_out_12_0_3;
  wire       [0:0]    subBytes_out_12_0_4;
  wire       [0:0]    subBytes_out_12_0_5;
  wire       [0:0]    subBytes_out_12_0_6;
  wire       [0:0]    subBytes_out_12_0_7;
  wire       [0:0]    subBytes_out_12_1_0;
  wire       [0:0]    subBytes_out_12_1_1;
  wire       [0:0]    subBytes_out_12_1_2;
  wire       [0:0]    subBytes_out_12_1_3;
  wire       [0:0]    subBytes_out_12_1_4;
  wire       [0:0]    subBytes_out_12_1_5;
  wire       [0:0]    subBytes_out_12_1_6;
  wire       [0:0]    subBytes_out_12_1_7;
  wire       [0:0]    subBytes_out_12_2_0;
  wire       [0:0]    subBytes_out_12_2_1;
  wire       [0:0]    subBytes_out_12_2_2;
  wire       [0:0]    subBytes_out_12_2_3;
  wire       [0:0]    subBytes_out_12_2_4;
  wire       [0:0]    subBytes_out_12_2_5;
  wire       [0:0]    subBytes_out_12_2_6;
  wire       [0:0]    subBytes_out_12_2_7;
  wire       [0:0]    subBytes_out_12_3_0;
  wire       [0:0]    subBytes_out_12_3_1;
  wire       [0:0]    subBytes_out_12_3_2;
  wire       [0:0]    subBytes_out_12_3_3;
  wire       [0:0]    subBytes_out_12_3_4;
  wire       [0:0]    subBytes_out_12_3_5;
  wire       [0:0]    subBytes_out_12_3_6;
  wire       [0:0]    subBytes_out_12_3_7;
  wire       [0:0]    subBytes_out_13_0_0;
  wire       [0:0]    subBytes_out_13_0_1;
  wire       [0:0]    subBytes_out_13_0_2;
  wire       [0:0]    subBytes_out_13_0_3;
  wire       [0:0]    subBytes_out_13_0_4;
  wire       [0:0]    subBytes_out_13_0_5;
  wire       [0:0]    subBytes_out_13_0_6;
  wire       [0:0]    subBytes_out_13_0_7;
  wire       [0:0]    subBytes_out_13_1_0;
  wire       [0:0]    subBytes_out_13_1_1;
  wire       [0:0]    subBytes_out_13_1_2;
  wire       [0:0]    subBytes_out_13_1_3;
  wire       [0:0]    subBytes_out_13_1_4;
  wire       [0:0]    subBytes_out_13_1_5;
  wire       [0:0]    subBytes_out_13_1_6;
  wire       [0:0]    subBytes_out_13_1_7;
  wire       [0:0]    subBytes_out_13_2_0;
  wire       [0:0]    subBytes_out_13_2_1;
  wire       [0:0]    subBytes_out_13_2_2;
  wire       [0:0]    subBytes_out_13_2_3;
  wire       [0:0]    subBytes_out_13_2_4;
  wire       [0:0]    subBytes_out_13_2_5;
  wire       [0:0]    subBytes_out_13_2_6;
  wire       [0:0]    subBytes_out_13_2_7;
  wire       [0:0]    subBytes_out_13_3_0;
  wire       [0:0]    subBytes_out_13_3_1;
  wire       [0:0]    subBytes_out_13_3_2;
  wire       [0:0]    subBytes_out_13_3_3;
  wire       [0:0]    subBytes_out_13_3_4;
  wire       [0:0]    subBytes_out_13_3_5;
  wire       [0:0]    subBytes_out_13_3_6;
  wire       [0:0]    subBytes_out_13_3_7;
  wire       [0:0]    subBytes_out_14_0_0;
  wire       [0:0]    subBytes_out_14_0_1;
  wire       [0:0]    subBytes_out_14_0_2;
  wire       [0:0]    subBytes_out_14_0_3;
  wire       [0:0]    subBytes_out_14_0_4;
  wire       [0:0]    subBytes_out_14_0_5;
  wire       [0:0]    subBytes_out_14_0_6;
  wire       [0:0]    subBytes_out_14_0_7;
  wire       [0:0]    subBytes_out_14_1_0;
  wire       [0:0]    subBytes_out_14_1_1;
  wire       [0:0]    subBytes_out_14_1_2;
  wire       [0:0]    subBytes_out_14_1_3;
  wire       [0:0]    subBytes_out_14_1_4;
  wire       [0:0]    subBytes_out_14_1_5;
  wire       [0:0]    subBytes_out_14_1_6;
  wire       [0:0]    subBytes_out_14_1_7;
  wire       [0:0]    subBytes_out_14_2_0;
  wire       [0:0]    subBytes_out_14_2_1;
  wire       [0:0]    subBytes_out_14_2_2;
  wire       [0:0]    subBytes_out_14_2_3;
  wire       [0:0]    subBytes_out_14_2_4;
  wire       [0:0]    subBytes_out_14_2_5;
  wire       [0:0]    subBytes_out_14_2_6;
  wire       [0:0]    subBytes_out_14_2_7;
  wire       [0:0]    subBytes_out_14_3_0;
  wire       [0:0]    subBytes_out_14_3_1;
  wire       [0:0]    subBytes_out_14_3_2;
  wire       [0:0]    subBytes_out_14_3_3;
  wire       [0:0]    subBytes_out_14_3_4;
  wire       [0:0]    subBytes_out_14_3_5;
  wire       [0:0]    subBytes_out_14_3_6;
  wire       [0:0]    subBytes_out_14_3_7;
  wire       [0:0]    subBytes_out_15_0_0;
  wire       [0:0]    subBytes_out_15_0_1;
  wire       [0:0]    subBytes_out_15_0_2;
  wire       [0:0]    subBytes_out_15_0_3;
  wire       [0:0]    subBytes_out_15_0_4;
  wire       [0:0]    subBytes_out_15_0_5;
  wire       [0:0]    subBytes_out_15_0_6;
  wire       [0:0]    subBytes_out_15_0_7;
  wire       [0:0]    subBytes_out_15_1_0;
  wire       [0:0]    subBytes_out_15_1_1;
  wire       [0:0]    subBytes_out_15_1_2;
  wire       [0:0]    subBytes_out_15_1_3;
  wire       [0:0]    subBytes_out_15_1_4;
  wire       [0:0]    subBytes_out_15_1_5;
  wire       [0:0]    subBytes_out_15_1_6;
  wire       [0:0]    subBytes_out_15_1_7;
  wire       [0:0]    subBytes_out_15_2_0;
  wire       [0:0]    subBytes_out_15_2_1;
  wire       [0:0]    subBytes_out_15_2_2;
  wire       [0:0]    subBytes_out_15_2_3;
  wire       [0:0]    subBytes_out_15_2_4;
  wire       [0:0]    subBytes_out_15_2_5;
  wire       [0:0]    subBytes_out_15_2_6;
  wire       [0:0]    subBytes_out_15_2_7;
  wire       [0:0]    subBytes_out_15_3_0;
  wire       [0:0]    subBytes_out_15_3_1;
  wire       [0:0]    subBytes_out_15_3_2;
  wire       [0:0]    subBytes_out_15_3_3;
  wire       [0:0]    subBytes_out_15_3_4;
  wire       [0:0]    subBytes_out_15_3_5;
  wire       [0:0]    subBytes_out_15_3_6;
  wire       [0:0]    subBytes_out_15_3_7;
  reg        [0:0]    roundReg_0_0_0;
  reg        [0:0]    roundReg_0_0_1;
  reg        [0:0]    roundReg_0_0_2;
  reg        [0:0]    roundReg_0_0_3;
  reg        [0:0]    roundReg_0_0_4;
  reg        [0:0]    roundReg_0_0_5;
  reg        [0:0]    roundReg_0_0_6;
  reg        [0:0]    roundReg_0_0_7;
  reg        [0:0]    roundReg_0_1_0;
  reg        [0:0]    roundReg_0_1_1;
  reg        [0:0]    roundReg_0_1_2;
  reg        [0:0]    roundReg_0_1_3;
  reg        [0:0]    roundReg_0_1_4;
  reg        [0:0]    roundReg_0_1_5;
  reg        [0:0]    roundReg_0_1_6;
  reg        [0:0]    roundReg_0_1_7;
  reg        [0:0]    roundReg_0_2_0;
  reg        [0:0]    roundReg_0_2_1;
  reg        [0:0]    roundReg_0_2_2;
  reg        [0:0]    roundReg_0_2_3;
  reg        [0:0]    roundReg_0_2_4;
  reg        [0:0]    roundReg_0_2_5;
  reg        [0:0]    roundReg_0_2_6;
  reg        [0:0]    roundReg_0_2_7;
  reg        [0:0]    roundReg_0_3_0;
  reg        [0:0]    roundReg_0_3_1;
  reg        [0:0]    roundReg_0_3_2;
  reg        [0:0]    roundReg_0_3_3;
  reg        [0:0]    roundReg_0_3_4;
  reg        [0:0]    roundReg_0_3_5;
  reg        [0:0]    roundReg_0_3_6;
  reg        [0:0]    roundReg_0_3_7;
  reg        [0:0]    roundReg_1_0_0;
  reg        [0:0]    roundReg_1_0_1;
  reg        [0:0]    roundReg_1_0_2;
  reg        [0:0]    roundReg_1_0_3;
  reg        [0:0]    roundReg_1_0_4;
  reg        [0:0]    roundReg_1_0_5;
  reg        [0:0]    roundReg_1_0_6;
  reg        [0:0]    roundReg_1_0_7;
  reg        [0:0]    roundReg_1_1_0;
  reg        [0:0]    roundReg_1_1_1;
  reg        [0:0]    roundReg_1_1_2;
  reg        [0:0]    roundReg_1_1_3;
  reg        [0:0]    roundReg_1_1_4;
  reg        [0:0]    roundReg_1_1_5;
  reg        [0:0]    roundReg_1_1_6;
  reg        [0:0]    roundReg_1_1_7;
  reg        [0:0]    roundReg_1_2_0;
  reg        [0:0]    roundReg_1_2_1;
  reg        [0:0]    roundReg_1_2_2;
  reg        [0:0]    roundReg_1_2_3;
  reg        [0:0]    roundReg_1_2_4;
  reg        [0:0]    roundReg_1_2_5;
  reg        [0:0]    roundReg_1_2_6;
  reg        [0:0]    roundReg_1_2_7;
  reg        [0:0]    roundReg_1_3_0;
  reg        [0:0]    roundReg_1_3_1;
  reg        [0:0]    roundReg_1_3_2;
  reg        [0:0]    roundReg_1_3_3;
  reg        [0:0]    roundReg_1_3_4;
  reg        [0:0]    roundReg_1_3_5;
  reg        [0:0]    roundReg_1_3_6;
  reg        [0:0]    roundReg_1_3_7;
  reg        [0:0]    roundReg_2_0_0;
  reg        [0:0]    roundReg_2_0_1;
  reg        [0:0]    roundReg_2_0_2;
  reg        [0:0]    roundReg_2_0_3;
  reg        [0:0]    roundReg_2_0_4;
  reg        [0:0]    roundReg_2_0_5;
  reg        [0:0]    roundReg_2_0_6;
  reg        [0:0]    roundReg_2_0_7;
  reg        [0:0]    roundReg_2_1_0;
  reg        [0:0]    roundReg_2_1_1;
  reg        [0:0]    roundReg_2_1_2;
  reg        [0:0]    roundReg_2_1_3;
  reg        [0:0]    roundReg_2_1_4;
  reg        [0:0]    roundReg_2_1_5;
  reg        [0:0]    roundReg_2_1_6;
  reg        [0:0]    roundReg_2_1_7;
  reg        [0:0]    roundReg_2_2_0;
  reg        [0:0]    roundReg_2_2_1;
  reg        [0:0]    roundReg_2_2_2;
  reg        [0:0]    roundReg_2_2_3;
  reg        [0:0]    roundReg_2_2_4;
  reg        [0:0]    roundReg_2_2_5;
  reg        [0:0]    roundReg_2_2_6;
  reg        [0:0]    roundReg_2_2_7;
  reg        [0:0]    roundReg_2_3_0;
  reg        [0:0]    roundReg_2_3_1;
  reg        [0:0]    roundReg_2_3_2;
  reg        [0:0]    roundReg_2_3_3;
  reg        [0:0]    roundReg_2_3_4;
  reg        [0:0]    roundReg_2_3_5;
  reg        [0:0]    roundReg_2_3_6;
  reg        [0:0]    roundReg_2_3_7;
  reg        [0:0]    roundReg_3_0_0;
  reg        [0:0]    roundReg_3_0_1;
  reg        [0:0]    roundReg_3_0_2;
  reg        [0:0]    roundReg_3_0_3;
  reg        [0:0]    roundReg_3_0_4;
  reg        [0:0]    roundReg_3_0_5;
  reg        [0:0]    roundReg_3_0_6;
  reg        [0:0]    roundReg_3_0_7;
  reg        [0:0]    roundReg_3_1_0;
  reg        [0:0]    roundReg_3_1_1;
  reg        [0:0]    roundReg_3_1_2;
  reg        [0:0]    roundReg_3_1_3;
  reg        [0:0]    roundReg_3_1_4;
  reg        [0:0]    roundReg_3_1_5;
  reg        [0:0]    roundReg_3_1_6;
  reg        [0:0]    roundReg_3_1_7;
  reg        [0:0]    roundReg_3_2_0;
  reg        [0:0]    roundReg_3_2_1;
  reg        [0:0]    roundReg_3_2_2;
  reg        [0:0]    roundReg_3_2_3;
  reg        [0:0]    roundReg_3_2_4;
  reg        [0:0]    roundReg_3_2_5;
  reg        [0:0]    roundReg_3_2_6;
  reg        [0:0]    roundReg_3_2_7;
  reg        [0:0]    roundReg_3_3_0;
  reg        [0:0]    roundReg_3_3_1;
  reg        [0:0]    roundReg_3_3_2;
  reg        [0:0]    roundReg_3_3_3;
  reg        [0:0]    roundReg_3_3_4;
  reg        [0:0]    roundReg_3_3_5;
  reg        [0:0]    roundReg_3_3_6;
  reg        [0:0]    roundReg_3_3_7;
  reg        [0:0]    roundReg_4_0_0;
  reg        [0:0]    roundReg_4_0_1;
  reg        [0:0]    roundReg_4_0_2;
  reg        [0:0]    roundReg_4_0_3;
  reg        [0:0]    roundReg_4_0_4;
  reg        [0:0]    roundReg_4_0_5;
  reg        [0:0]    roundReg_4_0_6;
  reg        [0:0]    roundReg_4_0_7;
  reg        [0:0]    roundReg_4_1_0;
  reg        [0:0]    roundReg_4_1_1;
  reg        [0:0]    roundReg_4_1_2;
  reg        [0:0]    roundReg_4_1_3;
  reg        [0:0]    roundReg_4_1_4;
  reg        [0:0]    roundReg_4_1_5;
  reg        [0:0]    roundReg_4_1_6;
  reg        [0:0]    roundReg_4_1_7;
  reg        [0:0]    roundReg_4_2_0;
  reg        [0:0]    roundReg_4_2_1;
  reg        [0:0]    roundReg_4_2_2;
  reg        [0:0]    roundReg_4_2_3;
  reg        [0:0]    roundReg_4_2_4;
  reg        [0:0]    roundReg_4_2_5;
  reg        [0:0]    roundReg_4_2_6;
  reg        [0:0]    roundReg_4_2_7;
  reg        [0:0]    roundReg_4_3_0;
  reg        [0:0]    roundReg_4_3_1;
  reg        [0:0]    roundReg_4_3_2;
  reg        [0:0]    roundReg_4_3_3;
  reg        [0:0]    roundReg_4_3_4;
  reg        [0:0]    roundReg_4_3_5;
  reg        [0:0]    roundReg_4_3_6;
  reg        [0:0]    roundReg_4_3_7;
  reg        [0:0]    roundReg_5_0_0;
  reg        [0:0]    roundReg_5_0_1;
  reg        [0:0]    roundReg_5_0_2;
  reg        [0:0]    roundReg_5_0_3;
  reg        [0:0]    roundReg_5_0_4;
  reg        [0:0]    roundReg_5_0_5;
  reg        [0:0]    roundReg_5_0_6;
  reg        [0:0]    roundReg_5_0_7;
  reg        [0:0]    roundReg_5_1_0;
  reg        [0:0]    roundReg_5_1_1;
  reg        [0:0]    roundReg_5_1_2;
  reg        [0:0]    roundReg_5_1_3;
  reg        [0:0]    roundReg_5_1_4;
  reg        [0:0]    roundReg_5_1_5;
  reg        [0:0]    roundReg_5_1_6;
  reg        [0:0]    roundReg_5_1_7;
  reg        [0:0]    roundReg_5_2_0;
  reg        [0:0]    roundReg_5_2_1;
  reg        [0:0]    roundReg_5_2_2;
  reg        [0:0]    roundReg_5_2_3;
  reg        [0:0]    roundReg_5_2_4;
  reg        [0:0]    roundReg_5_2_5;
  reg        [0:0]    roundReg_5_2_6;
  reg        [0:0]    roundReg_5_2_7;
  reg        [0:0]    roundReg_5_3_0;
  reg        [0:0]    roundReg_5_3_1;
  reg        [0:0]    roundReg_5_3_2;
  reg        [0:0]    roundReg_5_3_3;
  reg        [0:0]    roundReg_5_3_4;
  reg        [0:0]    roundReg_5_3_5;
  reg        [0:0]    roundReg_5_3_6;
  reg        [0:0]    roundReg_5_3_7;
  reg        [0:0]    roundReg_6_0_0;
  reg        [0:0]    roundReg_6_0_1;
  reg        [0:0]    roundReg_6_0_2;
  reg        [0:0]    roundReg_6_0_3;
  reg        [0:0]    roundReg_6_0_4;
  reg        [0:0]    roundReg_6_0_5;
  reg        [0:0]    roundReg_6_0_6;
  reg        [0:0]    roundReg_6_0_7;
  reg        [0:0]    roundReg_6_1_0;
  reg        [0:0]    roundReg_6_1_1;
  reg        [0:0]    roundReg_6_1_2;
  reg        [0:0]    roundReg_6_1_3;
  reg        [0:0]    roundReg_6_1_4;
  reg        [0:0]    roundReg_6_1_5;
  reg        [0:0]    roundReg_6_1_6;
  reg        [0:0]    roundReg_6_1_7;
  reg        [0:0]    roundReg_6_2_0;
  reg        [0:0]    roundReg_6_2_1;
  reg        [0:0]    roundReg_6_2_2;
  reg        [0:0]    roundReg_6_2_3;
  reg        [0:0]    roundReg_6_2_4;
  reg        [0:0]    roundReg_6_2_5;
  reg        [0:0]    roundReg_6_2_6;
  reg        [0:0]    roundReg_6_2_7;
  reg        [0:0]    roundReg_6_3_0;
  reg        [0:0]    roundReg_6_3_1;
  reg        [0:0]    roundReg_6_3_2;
  reg        [0:0]    roundReg_6_3_3;
  reg        [0:0]    roundReg_6_3_4;
  reg        [0:0]    roundReg_6_3_5;
  reg        [0:0]    roundReg_6_3_6;
  reg        [0:0]    roundReg_6_3_7;
  reg        [0:0]    roundReg_7_0_0;
  reg        [0:0]    roundReg_7_0_1;
  reg        [0:0]    roundReg_7_0_2;
  reg        [0:0]    roundReg_7_0_3;
  reg        [0:0]    roundReg_7_0_4;
  reg        [0:0]    roundReg_7_0_5;
  reg        [0:0]    roundReg_7_0_6;
  reg        [0:0]    roundReg_7_0_7;
  reg        [0:0]    roundReg_7_1_0;
  reg        [0:0]    roundReg_7_1_1;
  reg        [0:0]    roundReg_7_1_2;
  reg        [0:0]    roundReg_7_1_3;
  reg        [0:0]    roundReg_7_1_4;
  reg        [0:0]    roundReg_7_1_5;
  reg        [0:0]    roundReg_7_1_6;
  reg        [0:0]    roundReg_7_1_7;
  reg        [0:0]    roundReg_7_2_0;
  reg        [0:0]    roundReg_7_2_1;
  reg        [0:0]    roundReg_7_2_2;
  reg        [0:0]    roundReg_7_2_3;
  reg        [0:0]    roundReg_7_2_4;
  reg        [0:0]    roundReg_7_2_5;
  reg        [0:0]    roundReg_7_2_6;
  reg        [0:0]    roundReg_7_2_7;
  reg        [0:0]    roundReg_7_3_0;
  reg        [0:0]    roundReg_7_3_1;
  reg        [0:0]    roundReg_7_3_2;
  reg        [0:0]    roundReg_7_3_3;
  reg        [0:0]    roundReg_7_3_4;
  reg        [0:0]    roundReg_7_3_5;
  reg        [0:0]    roundReg_7_3_6;
  reg        [0:0]    roundReg_7_3_7;
  reg        [0:0]    roundReg_8_0_0;
  reg        [0:0]    roundReg_8_0_1;
  reg        [0:0]    roundReg_8_0_2;
  reg        [0:0]    roundReg_8_0_3;
  reg        [0:0]    roundReg_8_0_4;
  reg        [0:0]    roundReg_8_0_5;
  reg        [0:0]    roundReg_8_0_6;
  reg        [0:0]    roundReg_8_0_7;
  reg        [0:0]    roundReg_8_1_0;
  reg        [0:0]    roundReg_8_1_1;
  reg        [0:0]    roundReg_8_1_2;
  reg        [0:0]    roundReg_8_1_3;
  reg        [0:0]    roundReg_8_1_4;
  reg        [0:0]    roundReg_8_1_5;
  reg        [0:0]    roundReg_8_1_6;
  reg        [0:0]    roundReg_8_1_7;
  reg        [0:0]    roundReg_8_2_0;
  reg        [0:0]    roundReg_8_2_1;
  reg        [0:0]    roundReg_8_2_2;
  reg        [0:0]    roundReg_8_2_3;
  reg        [0:0]    roundReg_8_2_4;
  reg        [0:0]    roundReg_8_2_5;
  reg        [0:0]    roundReg_8_2_6;
  reg        [0:0]    roundReg_8_2_7;
  reg        [0:0]    roundReg_8_3_0;
  reg        [0:0]    roundReg_8_3_1;
  reg        [0:0]    roundReg_8_3_2;
  reg        [0:0]    roundReg_8_3_3;
  reg        [0:0]    roundReg_8_3_4;
  reg        [0:0]    roundReg_8_3_5;
  reg        [0:0]    roundReg_8_3_6;
  reg        [0:0]    roundReg_8_3_7;
  reg        [0:0]    roundReg_9_0_0;
  reg        [0:0]    roundReg_9_0_1;
  reg        [0:0]    roundReg_9_0_2;
  reg        [0:0]    roundReg_9_0_3;
  reg        [0:0]    roundReg_9_0_4;
  reg        [0:0]    roundReg_9_0_5;
  reg        [0:0]    roundReg_9_0_6;
  reg        [0:0]    roundReg_9_0_7;
  reg        [0:0]    roundReg_9_1_0;
  reg        [0:0]    roundReg_9_1_1;
  reg        [0:0]    roundReg_9_1_2;
  reg        [0:0]    roundReg_9_1_3;
  reg        [0:0]    roundReg_9_1_4;
  reg        [0:0]    roundReg_9_1_5;
  reg        [0:0]    roundReg_9_1_6;
  reg        [0:0]    roundReg_9_1_7;
  reg        [0:0]    roundReg_9_2_0;
  reg        [0:0]    roundReg_9_2_1;
  reg        [0:0]    roundReg_9_2_2;
  reg        [0:0]    roundReg_9_2_3;
  reg        [0:0]    roundReg_9_2_4;
  reg        [0:0]    roundReg_9_2_5;
  reg        [0:0]    roundReg_9_2_6;
  reg        [0:0]    roundReg_9_2_7;
  reg        [0:0]    roundReg_9_3_0;
  reg        [0:0]    roundReg_9_3_1;
  reg        [0:0]    roundReg_9_3_2;
  reg        [0:0]    roundReg_9_3_3;
  reg        [0:0]    roundReg_9_3_4;
  reg        [0:0]    roundReg_9_3_5;
  reg        [0:0]    roundReg_9_3_6;
  reg        [0:0]    roundReg_9_3_7;
  reg        [0:0]    roundReg_10_0_0;
  reg        [0:0]    roundReg_10_0_1;
  reg        [0:0]    roundReg_10_0_2;
  reg        [0:0]    roundReg_10_0_3;
  reg        [0:0]    roundReg_10_0_4;
  reg        [0:0]    roundReg_10_0_5;
  reg        [0:0]    roundReg_10_0_6;
  reg        [0:0]    roundReg_10_0_7;
  reg        [0:0]    roundReg_10_1_0;
  reg        [0:0]    roundReg_10_1_1;
  reg        [0:0]    roundReg_10_1_2;
  reg        [0:0]    roundReg_10_1_3;
  reg        [0:0]    roundReg_10_1_4;
  reg        [0:0]    roundReg_10_1_5;
  reg        [0:0]    roundReg_10_1_6;
  reg        [0:0]    roundReg_10_1_7;
  reg        [0:0]    roundReg_10_2_0;
  reg        [0:0]    roundReg_10_2_1;
  reg        [0:0]    roundReg_10_2_2;
  reg        [0:0]    roundReg_10_2_3;
  reg        [0:0]    roundReg_10_2_4;
  reg        [0:0]    roundReg_10_2_5;
  reg        [0:0]    roundReg_10_2_6;
  reg        [0:0]    roundReg_10_2_7;
  reg        [0:0]    roundReg_10_3_0;
  reg        [0:0]    roundReg_10_3_1;
  reg        [0:0]    roundReg_10_3_2;
  reg        [0:0]    roundReg_10_3_3;
  reg        [0:0]    roundReg_10_3_4;
  reg        [0:0]    roundReg_10_3_5;
  reg        [0:0]    roundReg_10_3_6;
  reg        [0:0]    roundReg_10_3_7;
  reg        [0:0]    roundReg_11_0_0;
  reg        [0:0]    roundReg_11_0_1;
  reg        [0:0]    roundReg_11_0_2;
  reg        [0:0]    roundReg_11_0_3;
  reg        [0:0]    roundReg_11_0_4;
  reg        [0:0]    roundReg_11_0_5;
  reg        [0:0]    roundReg_11_0_6;
  reg        [0:0]    roundReg_11_0_7;
  reg        [0:0]    roundReg_11_1_0;
  reg        [0:0]    roundReg_11_1_1;
  reg        [0:0]    roundReg_11_1_2;
  reg        [0:0]    roundReg_11_1_3;
  reg        [0:0]    roundReg_11_1_4;
  reg        [0:0]    roundReg_11_1_5;
  reg        [0:0]    roundReg_11_1_6;
  reg        [0:0]    roundReg_11_1_7;
  reg        [0:0]    roundReg_11_2_0;
  reg        [0:0]    roundReg_11_2_1;
  reg        [0:0]    roundReg_11_2_2;
  reg        [0:0]    roundReg_11_2_3;
  reg        [0:0]    roundReg_11_2_4;
  reg        [0:0]    roundReg_11_2_5;
  reg        [0:0]    roundReg_11_2_6;
  reg        [0:0]    roundReg_11_2_7;
  reg        [0:0]    roundReg_11_3_0;
  reg        [0:0]    roundReg_11_3_1;
  reg        [0:0]    roundReg_11_3_2;
  reg        [0:0]    roundReg_11_3_3;
  reg        [0:0]    roundReg_11_3_4;
  reg        [0:0]    roundReg_11_3_5;
  reg        [0:0]    roundReg_11_3_6;
  reg        [0:0]    roundReg_11_3_7;
  reg        [0:0]    roundReg_12_0_0;
  reg        [0:0]    roundReg_12_0_1;
  reg        [0:0]    roundReg_12_0_2;
  reg        [0:0]    roundReg_12_0_3;
  reg        [0:0]    roundReg_12_0_4;
  reg        [0:0]    roundReg_12_0_5;
  reg        [0:0]    roundReg_12_0_6;
  reg        [0:0]    roundReg_12_0_7;
  reg        [0:0]    roundReg_12_1_0;
  reg        [0:0]    roundReg_12_1_1;
  reg        [0:0]    roundReg_12_1_2;
  reg        [0:0]    roundReg_12_1_3;
  reg        [0:0]    roundReg_12_1_4;
  reg        [0:0]    roundReg_12_1_5;
  reg        [0:0]    roundReg_12_1_6;
  reg        [0:0]    roundReg_12_1_7;
  reg        [0:0]    roundReg_12_2_0;
  reg        [0:0]    roundReg_12_2_1;
  reg        [0:0]    roundReg_12_2_2;
  reg        [0:0]    roundReg_12_2_3;
  reg        [0:0]    roundReg_12_2_4;
  reg        [0:0]    roundReg_12_2_5;
  reg        [0:0]    roundReg_12_2_6;
  reg        [0:0]    roundReg_12_2_7;
  reg        [0:0]    roundReg_12_3_0;
  reg        [0:0]    roundReg_12_3_1;
  reg        [0:0]    roundReg_12_3_2;
  reg        [0:0]    roundReg_12_3_3;
  reg        [0:0]    roundReg_12_3_4;
  reg        [0:0]    roundReg_12_3_5;
  reg        [0:0]    roundReg_12_3_6;
  reg        [0:0]    roundReg_12_3_7;
  reg        [0:0]    roundReg_13_0_0;
  reg        [0:0]    roundReg_13_0_1;
  reg        [0:0]    roundReg_13_0_2;
  reg        [0:0]    roundReg_13_0_3;
  reg        [0:0]    roundReg_13_0_4;
  reg        [0:0]    roundReg_13_0_5;
  reg        [0:0]    roundReg_13_0_6;
  reg        [0:0]    roundReg_13_0_7;
  reg        [0:0]    roundReg_13_1_0;
  reg        [0:0]    roundReg_13_1_1;
  reg        [0:0]    roundReg_13_1_2;
  reg        [0:0]    roundReg_13_1_3;
  reg        [0:0]    roundReg_13_1_4;
  reg        [0:0]    roundReg_13_1_5;
  reg        [0:0]    roundReg_13_1_6;
  reg        [0:0]    roundReg_13_1_7;
  reg        [0:0]    roundReg_13_2_0;
  reg        [0:0]    roundReg_13_2_1;
  reg        [0:0]    roundReg_13_2_2;
  reg        [0:0]    roundReg_13_2_3;
  reg        [0:0]    roundReg_13_2_4;
  reg        [0:0]    roundReg_13_2_5;
  reg        [0:0]    roundReg_13_2_6;
  reg        [0:0]    roundReg_13_2_7;
  reg        [0:0]    roundReg_13_3_0;
  reg        [0:0]    roundReg_13_3_1;
  reg        [0:0]    roundReg_13_3_2;
  reg        [0:0]    roundReg_13_3_3;
  reg        [0:0]    roundReg_13_3_4;
  reg        [0:0]    roundReg_13_3_5;
  reg        [0:0]    roundReg_13_3_6;
  reg        [0:0]    roundReg_13_3_7;
  reg        [0:0]    roundReg_14_0_0;
  reg        [0:0]    roundReg_14_0_1;
  reg        [0:0]    roundReg_14_0_2;
  reg        [0:0]    roundReg_14_0_3;
  reg        [0:0]    roundReg_14_0_4;
  reg        [0:0]    roundReg_14_0_5;
  reg        [0:0]    roundReg_14_0_6;
  reg        [0:0]    roundReg_14_0_7;
  reg        [0:0]    roundReg_14_1_0;
  reg        [0:0]    roundReg_14_1_1;
  reg        [0:0]    roundReg_14_1_2;
  reg        [0:0]    roundReg_14_1_3;
  reg        [0:0]    roundReg_14_1_4;
  reg        [0:0]    roundReg_14_1_5;
  reg        [0:0]    roundReg_14_1_6;
  reg        [0:0]    roundReg_14_1_7;
  reg        [0:0]    roundReg_14_2_0;
  reg        [0:0]    roundReg_14_2_1;
  reg        [0:0]    roundReg_14_2_2;
  reg        [0:0]    roundReg_14_2_3;
  reg        [0:0]    roundReg_14_2_4;
  reg        [0:0]    roundReg_14_2_5;
  reg        [0:0]    roundReg_14_2_6;
  reg        [0:0]    roundReg_14_2_7;
  reg        [0:0]    roundReg_14_3_0;
  reg        [0:0]    roundReg_14_3_1;
  reg        [0:0]    roundReg_14_3_2;
  reg        [0:0]    roundReg_14_3_3;
  reg        [0:0]    roundReg_14_3_4;
  reg        [0:0]    roundReg_14_3_5;
  reg        [0:0]    roundReg_14_3_6;
  reg        [0:0]    roundReg_14_3_7;
  reg        [0:0]    roundReg_15_0_0;
  reg        [0:0]    roundReg_15_0_1;
  reg        [0:0]    roundReg_15_0_2;
  reg        [0:0]    roundReg_15_0_3;
  reg        [0:0]    roundReg_15_0_4;
  reg        [0:0]    roundReg_15_0_5;
  reg        [0:0]    roundReg_15_0_6;
  reg        [0:0]    roundReg_15_0_7;
  reg        [0:0]    roundReg_15_1_0;
  reg        [0:0]    roundReg_15_1_1;
  reg        [0:0]    roundReg_15_1_2;
  reg        [0:0]    roundReg_15_1_3;
  reg        [0:0]    roundReg_15_1_4;
  reg        [0:0]    roundReg_15_1_5;
  reg        [0:0]    roundReg_15_1_6;
  reg        [0:0]    roundReg_15_1_7;
  reg        [0:0]    roundReg_15_2_0;
  reg        [0:0]    roundReg_15_2_1;
  reg        [0:0]    roundReg_15_2_2;
  reg        [0:0]    roundReg_15_2_3;
  reg        [0:0]    roundReg_15_2_4;
  reg        [0:0]    roundReg_15_2_5;
  reg        [0:0]    roundReg_15_2_6;
  reg        [0:0]    roundReg_15_2_7;
  reg        [0:0]    roundReg_15_3_0;
  reg        [0:0]    roundReg_15_3_1;
  reg        [0:0]    roundReg_15_3_2;
  reg        [0:0]    roundReg_15_3_3;
  reg        [0:0]    roundReg_15_3_4;
  reg        [0:0]    roundReg_15_3_5;
  reg        [0:0]    roundReg_15_3_6;
  reg        [0:0]    roundReg_15_3_7;

  AES_KeyAddition keyAdd (
    .port_state_in_0_0_0   (port_state_in_0_0_0         ), //i
    .port_state_in_0_0_1   (port_state_in_0_0_1         ), //i
    .port_state_in_0_0_2   (port_state_in_0_0_2         ), //i
    .port_state_in_0_0_3   (port_state_in_0_0_3         ), //i
    .port_state_in_0_0_4   (port_state_in_0_0_4         ), //i
    .port_state_in_0_0_5   (port_state_in_0_0_5         ), //i
    .port_state_in_0_0_6   (port_state_in_0_0_6         ), //i
    .port_state_in_0_0_7   (port_state_in_0_0_7         ), //i
    .port_state_in_0_1_0   (port_state_in_0_1_0         ), //i
    .port_state_in_0_1_1   (port_state_in_0_1_1         ), //i
    .port_state_in_0_1_2   (port_state_in_0_1_2         ), //i
    .port_state_in_0_1_3   (port_state_in_0_1_3         ), //i
    .port_state_in_0_1_4   (port_state_in_0_1_4         ), //i
    .port_state_in_0_1_5   (port_state_in_0_1_5         ), //i
    .port_state_in_0_1_6   (port_state_in_0_1_6         ), //i
    .port_state_in_0_1_7   (port_state_in_0_1_7         ), //i
    .port_state_in_0_2_0   (port_state_in_0_2_0         ), //i
    .port_state_in_0_2_1   (port_state_in_0_2_1         ), //i
    .port_state_in_0_2_2   (port_state_in_0_2_2         ), //i
    .port_state_in_0_2_3   (port_state_in_0_2_3         ), //i
    .port_state_in_0_2_4   (port_state_in_0_2_4         ), //i
    .port_state_in_0_2_5   (port_state_in_0_2_5         ), //i
    .port_state_in_0_2_6   (port_state_in_0_2_6         ), //i
    .port_state_in_0_2_7   (port_state_in_0_2_7         ), //i
    .port_state_in_0_3_0   (port_state_in_0_3_0         ), //i
    .port_state_in_0_3_1   (port_state_in_0_3_1         ), //i
    .port_state_in_0_3_2   (port_state_in_0_3_2         ), //i
    .port_state_in_0_3_3   (port_state_in_0_3_3         ), //i
    .port_state_in_0_3_4   (port_state_in_0_3_4         ), //i
    .port_state_in_0_3_5   (port_state_in_0_3_5         ), //i
    .port_state_in_0_3_6   (port_state_in_0_3_6         ), //i
    .port_state_in_0_3_7   (port_state_in_0_3_7         ), //i
    .port_state_in_1_0_0   (port_state_in_1_0_0         ), //i
    .port_state_in_1_0_1   (port_state_in_1_0_1         ), //i
    .port_state_in_1_0_2   (port_state_in_1_0_2         ), //i
    .port_state_in_1_0_3   (port_state_in_1_0_3         ), //i
    .port_state_in_1_0_4   (port_state_in_1_0_4         ), //i
    .port_state_in_1_0_5   (port_state_in_1_0_5         ), //i
    .port_state_in_1_0_6   (port_state_in_1_0_6         ), //i
    .port_state_in_1_0_7   (port_state_in_1_0_7         ), //i
    .port_state_in_1_1_0   (port_state_in_1_1_0         ), //i
    .port_state_in_1_1_1   (port_state_in_1_1_1         ), //i
    .port_state_in_1_1_2   (port_state_in_1_1_2         ), //i
    .port_state_in_1_1_3   (port_state_in_1_1_3         ), //i
    .port_state_in_1_1_4   (port_state_in_1_1_4         ), //i
    .port_state_in_1_1_5   (port_state_in_1_1_5         ), //i
    .port_state_in_1_1_6   (port_state_in_1_1_6         ), //i
    .port_state_in_1_1_7   (port_state_in_1_1_7         ), //i
    .port_state_in_1_2_0   (port_state_in_1_2_0         ), //i
    .port_state_in_1_2_1   (port_state_in_1_2_1         ), //i
    .port_state_in_1_2_2   (port_state_in_1_2_2         ), //i
    .port_state_in_1_2_3   (port_state_in_1_2_3         ), //i
    .port_state_in_1_2_4   (port_state_in_1_2_4         ), //i
    .port_state_in_1_2_5   (port_state_in_1_2_5         ), //i
    .port_state_in_1_2_6   (port_state_in_1_2_6         ), //i
    .port_state_in_1_2_7   (port_state_in_1_2_7         ), //i
    .port_state_in_1_3_0   (port_state_in_1_3_0         ), //i
    .port_state_in_1_3_1   (port_state_in_1_3_1         ), //i
    .port_state_in_1_3_2   (port_state_in_1_3_2         ), //i
    .port_state_in_1_3_3   (port_state_in_1_3_3         ), //i
    .port_state_in_1_3_4   (port_state_in_1_3_4         ), //i
    .port_state_in_1_3_5   (port_state_in_1_3_5         ), //i
    .port_state_in_1_3_6   (port_state_in_1_3_6         ), //i
    .port_state_in_1_3_7   (port_state_in_1_3_7         ), //i
    .port_state_in_2_0_0   (port_state_in_2_0_0         ), //i
    .port_state_in_2_0_1   (port_state_in_2_0_1         ), //i
    .port_state_in_2_0_2   (port_state_in_2_0_2         ), //i
    .port_state_in_2_0_3   (port_state_in_2_0_3         ), //i
    .port_state_in_2_0_4   (port_state_in_2_0_4         ), //i
    .port_state_in_2_0_5   (port_state_in_2_0_5         ), //i
    .port_state_in_2_0_6   (port_state_in_2_0_6         ), //i
    .port_state_in_2_0_7   (port_state_in_2_0_7         ), //i
    .port_state_in_2_1_0   (port_state_in_2_1_0         ), //i
    .port_state_in_2_1_1   (port_state_in_2_1_1         ), //i
    .port_state_in_2_1_2   (port_state_in_2_1_2         ), //i
    .port_state_in_2_1_3   (port_state_in_2_1_3         ), //i
    .port_state_in_2_1_4   (port_state_in_2_1_4         ), //i
    .port_state_in_2_1_5   (port_state_in_2_1_5         ), //i
    .port_state_in_2_1_6   (port_state_in_2_1_6         ), //i
    .port_state_in_2_1_7   (port_state_in_2_1_7         ), //i
    .port_state_in_2_2_0   (port_state_in_2_2_0         ), //i
    .port_state_in_2_2_1   (port_state_in_2_2_1         ), //i
    .port_state_in_2_2_2   (port_state_in_2_2_2         ), //i
    .port_state_in_2_2_3   (port_state_in_2_2_3         ), //i
    .port_state_in_2_2_4   (port_state_in_2_2_4         ), //i
    .port_state_in_2_2_5   (port_state_in_2_2_5         ), //i
    .port_state_in_2_2_6   (port_state_in_2_2_6         ), //i
    .port_state_in_2_2_7   (port_state_in_2_2_7         ), //i
    .port_state_in_2_3_0   (port_state_in_2_3_0         ), //i
    .port_state_in_2_3_1   (port_state_in_2_3_1         ), //i
    .port_state_in_2_3_2   (port_state_in_2_3_2         ), //i
    .port_state_in_2_3_3   (port_state_in_2_3_3         ), //i
    .port_state_in_2_3_4   (port_state_in_2_3_4         ), //i
    .port_state_in_2_3_5   (port_state_in_2_3_5         ), //i
    .port_state_in_2_3_6   (port_state_in_2_3_6         ), //i
    .port_state_in_2_3_7   (port_state_in_2_3_7         ), //i
    .port_state_in_3_0_0   (port_state_in_3_0_0         ), //i
    .port_state_in_3_0_1   (port_state_in_3_0_1         ), //i
    .port_state_in_3_0_2   (port_state_in_3_0_2         ), //i
    .port_state_in_3_0_3   (port_state_in_3_0_3         ), //i
    .port_state_in_3_0_4   (port_state_in_3_0_4         ), //i
    .port_state_in_3_0_5   (port_state_in_3_0_5         ), //i
    .port_state_in_3_0_6   (port_state_in_3_0_6         ), //i
    .port_state_in_3_0_7   (port_state_in_3_0_7         ), //i
    .port_state_in_3_1_0   (port_state_in_3_1_0         ), //i
    .port_state_in_3_1_1   (port_state_in_3_1_1         ), //i
    .port_state_in_3_1_2   (port_state_in_3_1_2         ), //i
    .port_state_in_3_1_3   (port_state_in_3_1_3         ), //i
    .port_state_in_3_1_4   (port_state_in_3_1_4         ), //i
    .port_state_in_3_1_5   (port_state_in_3_1_5         ), //i
    .port_state_in_3_1_6   (port_state_in_3_1_6         ), //i
    .port_state_in_3_1_7   (port_state_in_3_1_7         ), //i
    .port_state_in_3_2_0   (port_state_in_3_2_0         ), //i
    .port_state_in_3_2_1   (port_state_in_3_2_1         ), //i
    .port_state_in_3_2_2   (port_state_in_3_2_2         ), //i
    .port_state_in_3_2_3   (port_state_in_3_2_3         ), //i
    .port_state_in_3_2_4   (port_state_in_3_2_4         ), //i
    .port_state_in_3_2_5   (port_state_in_3_2_5         ), //i
    .port_state_in_3_2_6   (port_state_in_3_2_6         ), //i
    .port_state_in_3_2_7   (port_state_in_3_2_7         ), //i
    .port_state_in_3_3_0   (port_state_in_3_3_0         ), //i
    .port_state_in_3_3_1   (port_state_in_3_3_1         ), //i
    .port_state_in_3_3_2   (port_state_in_3_3_2         ), //i
    .port_state_in_3_3_3   (port_state_in_3_3_3         ), //i
    .port_state_in_3_3_4   (port_state_in_3_3_4         ), //i
    .port_state_in_3_3_5   (port_state_in_3_3_5         ), //i
    .port_state_in_3_3_6   (port_state_in_3_3_6         ), //i
    .port_state_in_3_3_7   (port_state_in_3_3_7         ), //i
    .port_state_in_4_0_0   (port_state_in_4_0_0         ), //i
    .port_state_in_4_0_1   (port_state_in_4_0_1         ), //i
    .port_state_in_4_0_2   (port_state_in_4_0_2         ), //i
    .port_state_in_4_0_3   (port_state_in_4_0_3         ), //i
    .port_state_in_4_0_4   (port_state_in_4_0_4         ), //i
    .port_state_in_4_0_5   (port_state_in_4_0_5         ), //i
    .port_state_in_4_0_6   (port_state_in_4_0_6         ), //i
    .port_state_in_4_0_7   (port_state_in_4_0_7         ), //i
    .port_state_in_4_1_0   (port_state_in_4_1_0         ), //i
    .port_state_in_4_1_1   (port_state_in_4_1_1         ), //i
    .port_state_in_4_1_2   (port_state_in_4_1_2         ), //i
    .port_state_in_4_1_3   (port_state_in_4_1_3         ), //i
    .port_state_in_4_1_4   (port_state_in_4_1_4         ), //i
    .port_state_in_4_1_5   (port_state_in_4_1_5         ), //i
    .port_state_in_4_1_6   (port_state_in_4_1_6         ), //i
    .port_state_in_4_1_7   (port_state_in_4_1_7         ), //i
    .port_state_in_4_2_0   (port_state_in_4_2_0         ), //i
    .port_state_in_4_2_1   (port_state_in_4_2_1         ), //i
    .port_state_in_4_2_2   (port_state_in_4_2_2         ), //i
    .port_state_in_4_2_3   (port_state_in_4_2_3         ), //i
    .port_state_in_4_2_4   (port_state_in_4_2_4         ), //i
    .port_state_in_4_2_5   (port_state_in_4_2_5         ), //i
    .port_state_in_4_2_6   (port_state_in_4_2_6         ), //i
    .port_state_in_4_2_7   (port_state_in_4_2_7         ), //i
    .port_state_in_4_3_0   (port_state_in_4_3_0         ), //i
    .port_state_in_4_3_1   (port_state_in_4_3_1         ), //i
    .port_state_in_4_3_2   (port_state_in_4_3_2         ), //i
    .port_state_in_4_3_3   (port_state_in_4_3_3         ), //i
    .port_state_in_4_3_4   (port_state_in_4_3_4         ), //i
    .port_state_in_4_3_5   (port_state_in_4_3_5         ), //i
    .port_state_in_4_3_6   (port_state_in_4_3_6         ), //i
    .port_state_in_4_3_7   (port_state_in_4_3_7         ), //i
    .port_state_in_5_0_0   (port_state_in_5_0_0         ), //i
    .port_state_in_5_0_1   (port_state_in_5_0_1         ), //i
    .port_state_in_5_0_2   (port_state_in_5_0_2         ), //i
    .port_state_in_5_0_3   (port_state_in_5_0_3         ), //i
    .port_state_in_5_0_4   (port_state_in_5_0_4         ), //i
    .port_state_in_5_0_5   (port_state_in_5_0_5         ), //i
    .port_state_in_5_0_6   (port_state_in_5_0_6         ), //i
    .port_state_in_5_0_7   (port_state_in_5_0_7         ), //i
    .port_state_in_5_1_0   (port_state_in_5_1_0         ), //i
    .port_state_in_5_1_1   (port_state_in_5_1_1         ), //i
    .port_state_in_5_1_2   (port_state_in_5_1_2         ), //i
    .port_state_in_5_1_3   (port_state_in_5_1_3         ), //i
    .port_state_in_5_1_4   (port_state_in_5_1_4         ), //i
    .port_state_in_5_1_5   (port_state_in_5_1_5         ), //i
    .port_state_in_5_1_6   (port_state_in_5_1_6         ), //i
    .port_state_in_5_1_7   (port_state_in_5_1_7         ), //i
    .port_state_in_5_2_0   (port_state_in_5_2_0         ), //i
    .port_state_in_5_2_1   (port_state_in_5_2_1         ), //i
    .port_state_in_5_2_2   (port_state_in_5_2_2         ), //i
    .port_state_in_5_2_3   (port_state_in_5_2_3         ), //i
    .port_state_in_5_2_4   (port_state_in_5_2_4         ), //i
    .port_state_in_5_2_5   (port_state_in_5_2_5         ), //i
    .port_state_in_5_2_6   (port_state_in_5_2_6         ), //i
    .port_state_in_5_2_7   (port_state_in_5_2_7         ), //i
    .port_state_in_5_3_0   (port_state_in_5_3_0         ), //i
    .port_state_in_5_3_1   (port_state_in_5_3_1         ), //i
    .port_state_in_5_3_2   (port_state_in_5_3_2         ), //i
    .port_state_in_5_3_3   (port_state_in_5_3_3         ), //i
    .port_state_in_5_3_4   (port_state_in_5_3_4         ), //i
    .port_state_in_5_3_5   (port_state_in_5_3_5         ), //i
    .port_state_in_5_3_6   (port_state_in_5_3_6         ), //i
    .port_state_in_5_3_7   (port_state_in_5_3_7         ), //i
    .port_state_in_6_0_0   (port_state_in_6_0_0         ), //i
    .port_state_in_6_0_1   (port_state_in_6_0_1         ), //i
    .port_state_in_6_0_2   (port_state_in_6_0_2         ), //i
    .port_state_in_6_0_3   (port_state_in_6_0_3         ), //i
    .port_state_in_6_0_4   (port_state_in_6_0_4         ), //i
    .port_state_in_6_0_5   (port_state_in_6_0_5         ), //i
    .port_state_in_6_0_6   (port_state_in_6_0_6         ), //i
    .port_state_in_6_0_7   (port_state_in_6_0_7         ), //i
    .port_state_in_6_1_0   (port_state_in_6_1_0         ), //i
    .port_state_in_6_1_1   (port_state_in_6_1_1         ), //i
    .port_state_in_6_1_2   (port_state_in_6_1_2         ), //i
    .port_state_in_6_1_3   (port_state_in_6_1_3         ), //i
    .port_state_in_6_1_4   (port_state_in_6_1_4         ), //i
    .port_state_in_6_1_5   (port_state_in_6_1_5         ), //i
    .port_state_in_6_1_6   (port_state_in_6_1_6         ), //i
    .port_state_in_6_1_7   (port_state_in_6_1_7         ), //i
    .port_state_in_6_2_0   (port_state_in_6_2_0         ), //i
    .port_state_in_6_2_1   (port_state_in_6_2_1         ), //i
    .port_state_in_6_2_2   (port_state_in_6_2_2         ), //i
    .port_state_in_6_2_3   (port_state_in_6_2_3         ), //i
    .port_state_in_6_2_4   (port_state_in_6_2_4         ), //i
    .port_state_in_6_2_5   (port_state_in_6_2_5         ), //i
    .port_state_in_6_2_6   (port_state_in_6_2_6         ), //i
    .port_state_in_6_2_7   (port_state_in_6_2_7         ), //i
    .port_state_in_6_3_0   (port_state_in_6_3_0         ), //i
    .port_state_in_6_3_1   (port_state_in_6_3_1         ), //i
    .port_state_in_6_3_2   (port_state_in_6_3_2         ), //i
    .port_state_in_6_3_3   (port_state_in_6_3_3         ), //i
    .port_state_in_6_3_4   (port_state_in_6_3_4         ), //i
    .port_state_in_6_3_5   (port_state_in_6_3_5         ), //i
    .port_state_in_6_3_6   (port_state_in_6_3_6         ), //i
    .port_state_in_6_3_7   (port_state_in_6_3_7         ), //i
    .port_state_in_7_0_0   (port_state_in_7_0_0         ), //i
    .port_state_in_7_0_1   (port_state_in_7_0_1         ), //i
    .port_state_in_7_0_2   (port_state_in_7_0_2         ), //i
    .port_state_in_7_0_3   (port_state_in_7_0_3         ), //i
    .port_state_in_7_0_4   (port_state_in_7_0_4         ), //i
    .port_state_in_7_0_5   (port_state_in_7_0_5         ), //i
    .port_state_in_7_0_6   (port_state_in_7_0_6         ), //i
    .port_state_in_7_0_7   (port_state_in_7_0_7         ), //i
    .port_state_in_7_1_0   (port_state_in_7_1_0         ), //i
    .port_state_in_7_1_1   (port_state_in_7_1_1         ), //i
    .port_state_in_7_1_2   (port_state_in_7_1_2         ), //i
    .port_state_in_7_1_3   (port_state_in_7_1_3         ), //i
    .port_state_in_7_1_4   (port_state_in_7_1_4         ), //i
    .port_state_in_7_1_5   (port_state_in_7_1_5         ), //i
    .port_state_in_7_1_6   (port_state_in_7_1_6         ), //i
    .port_state_in_7_1_7   (port_state_in_7_1_7         ), //i
    .port_state_in_7_2_0   (port_state_in_7_2_0         ), //i
    .port_state_in_7_2_1   (port_state_in_7_2_1         ), //i
    .port_state_in_7_2_2   (port_state_in_7_2_2         ), //i
    .port_state_in_7_2_3   (port_state_in_7_2_3         ), //i
    .port_state_in_7_2_4   (port_state_in_7_2_4         ), //i
    .port_state_in_7_2_5   (port_state_in_7_2_5         ), //i
    .port_state_in_7_2_6   (port_state_in_7_2_6         ), //i
    .port_state_in_7_2_7   (port_state_in_7_2_7         ), //i
    .port_state_in_7_3_0   (port_state_in_7_3_0         ), //i
    .port_state_in_7_3_1   (port_state_in_7_3_1         ), //i
    .port_state_in_7_3_2   (port_state_in_7_3_2         ), //i
    .port_state_in_7_3_3   (port_state_in_7_3_3         ), //i
    .port_state_in_7_3_4   (port_state_in_7_3_4         ), //i
    .port_state_in_7_3_5   (port_state_in_7_3_5         ), //i
    .port_state_in_7_3_6   (port_state_in_7_3_6         ), //i
    .port_state_in_7_3_7   (port_state_in_7_3_7         ), //i
    .port_state_in_8_0_0   (port_state_in_8_0_0         ), //i
    .port_state_in_8_0_1   (port_state_in_8_0_1         ), //i
    .port_state_in_8_0_2   (port_state_in_8_0_2         ), //i
    .port_state_in_8_0_3   (port_state_in_8_0_3         ), //i
    .port_state_in_8_0_4   (port_state_in_8_0_4         ), //i
    .port_state_in_8_0_5   (port_state_in_8_0_5         ), //i
    .port_state_in_8_0_6   (port_state_in_8_0_6         ), //i
    .port_state_in_8_0_7   (port_state_in_8_0_7         ), //i
    .port_state_in_8_1_0   (port_state_in_8_1_0         ), //i
    .port_state_in_8_1_1   (port_state_in_8_1_1         ), //i
    .port_state_in_8_1_2   (port_state_in_8_1_2         ), //i
    .port_state_in_8_1_3   (port_state_in_8_1_3         ), //i
    .port_state_in_8_1_4   (port_state_in_8_1_4         ), //i
    .port_state_in_8_1_5   (port_state_in_8_1_5         ), //i
    .port_state_in_8_1_6   (port_state_in_8_1_6         ), //i
    .port_state_in_8_1_7   (port_state_in_8_1_7         ), //i
    .port_state_in_8_2_0   (port_state_in_8_2_0         ), //i
    .port_state_in_8_2_1   (port_state_in_8_2_1         ), //i
    .port_state_in_8_2_2   (port_state_in_8_2_2         ), //i
    .port_state_in_8_2_3   (port_state_in_8_2_3         ), //i
    .port_state_in_8_2_4   (port_state_in_8_2_4         ), //i
    .port_state_in_8_2_5   (port_state_in_8_2_5         ), //i
    .port_state_in_8_2_6   (port_state_in_8_2_6         ), //i
    .port_state_in_8_2_7   (port_state_in_8_2_7         ), //i
    .port_state_in_8_3_0   (port_state_in_8_3_0         ), //i
    .port_state_in_8_3_1   (port_state_in_8_3_1         ), //i
    .port_state_in_8_3_2   (port_state_in_8_3_2         ), //i
    .port_state_in_8_3_3   (port_state_in_8_3_3         ), //i
    .port_state_in_8_3_4   (port_state_in_8_3_4         ), //i
    .port_state_in_8_3_5   (port_state_in_8_3_5         ), //i
    .port_state_in_8_3_6   (port_state_in_8_3_6         ), //i
    .port_state_in_8_3_7   (port_state_in_8_3_7         ), //i
    .port_state_in_9_0_0   (port_state_in_9_0_0         ), //i
    .port_state_in_9_0_1   (port_state_in_9_0_1         ), //i
    .port_state_in_9_0_2   (port_state_in_9_0_2         ), //i
    .port_state_in_9_0_3   (port_state_in_9_0_3         ), //i
    .port_state_in_9_0_4   (port_state_in_9_0_4         ), //i
    .port_state_in_9_0_5   (port_state_in_9_0_5         ), //i
    .port_state_in_9_0_6   (port_state_in_9_0_6         ), //i
    .port_state_in_9_0_7   (port_state_in_9_0_7         ), //i
    .port_state_in_9_1_0   (port_state_in_9_1_0         ), //i
    .port_state_in_9_1_1   (port_state_in_9_1_1         ), //i
    .port_state_in_9_1_2   (port_state_in_9_1_2         ), //i
    .port_state_in_9_1_3   (port_state_in_9_1_3         ), //i
    .port_state_in_9_1_4   (port_state_in_9_1_4         ), //i
    .port_state_in_9_1_5   (port_state_in_9_1_5         ), //i
    .port_state_in_9_1_6   (port_state_in_9_1_6         ), //i
    .port_state_in_9_1_7   (port_state_in_9_1_7         ), //i
    .port_state_in_9_2_0   (port_state_in_9_2_0         ), //i
    .port_state_in_9_2_1   (port_state_in_9_2_1         ), //i
    .port_state_in_9_2_2   (port_state_in_9_2_2         ), //i
    .port_state_in_9_2_3   (port_state_in_9_2_3         ), //i
    .port_state_in_9_2_4   (port_state_in_9_2_4         ), //i
    .port_state_in_9_2_5   (port_state_in_9_2_5         ), //i
    .port_state_in_9_2_6   (port_state_in_9_2_6         ), //i
    .port_state_in_9_2_7   (port_state_in_9_2_7         ), //i
    .port_state_in_9_3_0   (port_state_in_9_3_0         ), //i
    .port_state_in_9_3_1   (port_state_in_9_3_1         ), //i
    .port_state_in_9_3_2   (port_state_in_9_3_2         ), //i
    .port_state_in_9_3_3   (port_state_in_9_3_3         ), //i
    .port_state_in_9_3_4   (port_state_in_9_3_4         ), //i
    .port_state_in_9_3_5   (port_state_in_9_3_5         ), //i
    .port_state_in_9_3_6   (port_state_in_9_3_6         ), //i
    .port_state_in_9_3_7   (port_state_in_9_3_7         ), //i
    .port_state_in_10_0_0  (port_state_in_10_0_0        ), //i
    .port_state_in_10_0_1  (port_state_in_10_0_1        ), //i
    .port_state_in_10_0_2  (port_state_in_10_0_2        ), //i
    .port_state_in_10_0_3  (port_state_in_10_0_3        ), //i
    .port_state_in_10_0_4  (port_state_in_10_0_4        ), //i
    .port_state_in_10_0_5  (port_state_in_10_0_5        ), //i
    .port_state_in_10_0_6  (port_state_in_10_0_6        ), //i
    .port_state_in_10_0_7  (port_state_in_10_0_7        ), //i
    .port_state_in_10_1_0  (port_state_in_10_1_0        ), //i
    .port_state_in_10_1_1  (port_state_in_10_1_1        ), //i
    .port_state_in_10_1_2  (port_state_in_10_1_2        ), //i
    .port_state_in_10_1_3  (port_state_in_10_1_3        ), //i
    .port_state_in_10_1_4  (port_state_in_10_1_4        ), //i
    .port_state_in_10_1_5  (port_state_in_10_1_5        ), //i
    .port_state_in_10_1_6  (port_state_in_10_1_6        ), //i
    .port_state_in_10_1_7  (port_state_in_10_1_7        ), //i
    .port_state_in_10_2_0  (port_state_in_10_2_0        ), //i
    .port_state_in_10_2_1  (port_state_in_10_2_1        ), //i
    .port_state_in_10_2_2  (port_state_in_10_2_2        ), //i
    .port_state_in_10_2_3  (port_state_in_10_2_3        ), //i
    .port_state_in_10_2_4  (port_state_in_10_2_4        ), //i
    .port_state_in_10_2_5  (port_state_in_10_2_5        ), //i
    .port_state_in_10_2_6  (port_state_in_10_2_6        ), //i
    .port_state_in_10_2_7  (port_state_in_10_2_7        ), //i
    .port_state_in_10_3_0  (port_state_in_10_3_0        ), //i
    .port_state_in_10_3_1  (port_state_in_10_3_1        ), //i
    .port_state_in_10_3_2  (port_state_in_10_3_2        ), //i
    .port_state_in_10_3_3  (port_state_in_10_3_3        ), //i
    .port_state_in_10_3_4  (port_state_in_10_3_4        ), //i
    .port_state_in_10_3_5  (port_state_in_10_3_5        ), //i
    .port_state_in_10_3_6  (port_state_in_10_3_6        ), //i
    .port_state_in_10_3_7  (port_state_in_10_3_7        ), //i
    .port_state_in_11_0_0  (port_state_in_11_0_0        ), //i
    .port_state_in_11_0_1  (port_state_in_11_0_1        ), //i
    .port_state_in_11_0_2  (port_state_in_11_0_2        ), //i
    .port_state_in_11_0_3  (port_state_in_11_0_3        ), //i
    .port_state_in_11_0_4  (port_state_in_11_0_4        ), //i
    .port_state_in_11_0_5  (port_state_in_11_0_5        ), //i
    .port_state_in_11_0_6  (port_state_in_11_0_6        ), //i
    .port_state_in_11_0_7  (port_state_in_11_0_7        ), //i
    .port_state_in_11_1_0  (port_state_in_11_1_0        ), //i
    .port_state_in_11_1_1  (port_state_in_11_1_1        ), //i
    .port_state_in_11_1_2  (port_state_in_11_1_2        ), //i
    .port_state_in_11_1_3  (port_state_in_11_1_3        ), //i
    .port_state_in_11_1_4  (port_state_in_11_1_4        ), //i
    .port_state_in_11_1_5  (port_state_in_11_1_5        ), //i
    .port_state_in_11_1_6  (port_state_in_11_1_6        ), //i
    .port_state_in_11_1_7  (port_state_in_11_1_7        ), //i
    .port_state_in_11_2_0  (port_state_in_11_2_0        ), //i
    .port_state_in_11_2_1  (port_state_in_11_2_1        ), //i
    .port_state_in_11_2_2  (port_state_in_11_2_2        ), //i
    .port_state_in_11_2_3  (port_state_in_11_2_3        ), //i
    .port_state_in_11_2_4  (port_state_in_11_2_4        ), //i
    .port_state_in_11_2_5  (port_state_in_11_2_5        ), //i
    .port_state_in_11_2_6  (port_state_in_11_2_6        ), //i
    .port_state_in_11_2_7  (port_state_in_11_2_7        ), //i
    .port_state_in_11_3_0  (port_state_in_11_3_0        ), //i
    .port_state_in_11_3_1  (port_state_in_11_3_1        ), //i
    .port_state_in_11_3_2  (port_state_in_11_3_2        ), //i
    .port_state_in_11_3_3  (port_state_in_11_3_3        ), //i
    .port_state_in_11_3_4  (port_state_in_11_3_4        ), //i
    .port_state_in_11_3_5  (port_state_in_11_3_5        ), //i
    .port_state_in_11_3_6  (port_state_in_11_3_6        ), //i
    .port_state_in_11_3_7  (port_state_in_11_3_7        ), //i
    .port_state_in_12_0_0  (port_state_in_12_0_0        ), //i
    .port_state_in_12_0_1  (port_state_in_12_0_1        ), //i
    .port_state_in_12_0_2  (port_state_in_12_0_2        ), //i
    .port_state_in_12_0_3  (port_state_in_12_0_3        ), //i
    .port_state_in_12_0_4  (port_state_in_12_0_4        ), //i
    .port_state_in_12_0_5  (port_state_in_12_0_5        ), //i
    .port_state_in_12_0_6  (port_state_in_12_0_6        ), //i
    .port_state_in_12_0_7  (port_state_in_12_0_7        ), //i
    .port_state_in_12_1_0  (port_state_in_12_1_0        ), //i
    .port_state_in_12_1_1  (port_state_in_12_1_1        ), //i
    .port_state_in_12_1_2  (port_state_in_12_1_2        ), //i
    .port_state_in_12_1_3  (port_state_in_12_1_3        ), //i
    .port_state_in_12_1_4  (port_state_in_12_1_4        ), //i
    .port_state_in_12_1_5  (port_state_in_12_1_5        ), //i
    .port_state_in_12_1_6  (port_state_in_12_1_6        ), //i
    .port_state_in_12_1_7  (port_state_in_12_1_7        ), //i
    .port_state_in_12_2_0  (port_state_in_12_2_0        ), //i
    .port_state_in_12_2_1  (port_state_in_12_2_1        ), //i
    .port_state_in_12_2_2  (port_state_in_12_2_2        ), //i
    .port_state_in_12_2_3  (port_state_in_12_2_3        ), //i
    .port_state_in_12_2_4  (port_state_in_12_2_4        ), //i
    .port_state_in_12_2_5  (port_state_in_12_2_5        ), //i
    .port_state_in_12_2_6  (port_state_in_12_2_6        ), //i
    .port_state_in_12_2_7  (port_state_in_12_2_7        ), //i
    .port_state_in_12_3_0  (port_state_in_12_3_0        ), //i
    .port_state_in_12_3_1  (port_state_in_12_3_1        ), //i
    .port_state_in_12_3_2  (port_state_in_12_3_2        ), //i
    .port_state_in_12_3_3  (port_state_in_12_3_3        ), //i
    .port_state_in_12_3_4  (port_state_in_12_3_4        ), //i
    .port_state_in_12_3_5  (port_state_in_12_3_5        ), //i
    .port_state_in_12_3_6  (port_state_in_12_3_6        ), //i
    .port_state_in_12_3_7  (port_state_in_12_3_7        ), //i
    .port_state_in_13_0_0  (port_state_in_13_0_0        ), //i
    .port_state_in_13_0_1  (port_state_in_13_0_1        ), //i
    .port_state_in_13_0_2  (port_state_in_13_0_2        ), //i
    .port_state_in_13_0_3  (port_state_in_13_0_3        ), //i
    .port_state_in_13_0_4  (port_state_in_13_0_4        ), //i
    .port_state_in_13_0_5  (port_state_in_13_0_5        ), //i
    .port_state_in_13_0_6  (port_state_in_13_0_6        ), //i
    .port_state_in_13_0_7  (port_state_in_13_0_7        ), //i
    .port_state_in_13_1_0  (port_state_in_13_1_0        ), //i
    .port_state_in_13_1_1  (port_state_in_13_1_1        ), //i
    .port_state_in_13_1_2  (port_state_in_13_1_2        ), //i
    .port_state_in_13_1_3  (port_state_in_13_1_3        ), //i
    .port_state_in_13_1_4  (port_state_in_13_1_4        ), //i
    .port_state_in_13_1_5  (port_state_in_13_1_5        ), //i
    .port_state_in_13_1_6  (port_state_in_13_1_6        ), //i
    .port_state_in_13_1_7  (port_state_in_13_1_7        ), //i
    .port_state_in_13_2_0  (port_state_in_13_2_0        ), //i
    .port_state_in_13_2_1  (port_state_in_13_2_1        ), //i
    .port_state_in_13_2_2  (port_state_in_13_2_2        ), //i
    .port_state_in_13_2_3  (port_state_in_13_2_3        ), //i
    .port_state_in_13_2_4  (port_state_in_13_2_4        ), //i
    .port_state_in_13_2_5  (port_state_in_13_2_5        ), //i
    .port_state_in_13_2_6  (port_state_in_13_2_6        ), //i
    .port_state_in_13_2_7  (port_state_in_13_2_7        ), //i
    .port_state_in_13_3_0  (port_state_in_13_3_0        ), //i
    .port_state_in_13_3_1  (port_state_in_13_3_1        ), //i
    .port_state_in_13_3_2  (port_state_in_13_3_2        ), //i
    .port_state_in_13_3_3  (port_state_in_13_3_3        ), //i
    .port_state_in_13_3_4  (port_state_in_13_3_4        ), //i
    .port_state_in_13_3_5  (port_state_in_13_3_5        ), //i
    .port_state_in_13_3_6  (port_state_in_13_3_6        ), //i
    .port_state_in_13_3_7  (port_state_in_13_3_7        ), //i
    .port_state_in_14_0_0  (port_state_in_14_0_0        ), //i
    .port_state_in_14_0_1  (port_state_in_14_0_1        ), //i
    .port_state_in_14_0_2  (port_state_in_14_0_2        ), //i
    .port_state_in_14_0_3  (port_state_in_14_0_3        ), //i
    .port_state_in_14_0_4  (port_state_in_14_0_4        ), //i
    .port_state_in_14_0_5  (port_state_in_14_0_5        ), //i
    .port_state_in_14_0_6  (port_state_in_14_0_6        ), //i
    .port_state_in_14_0_7  (port_state_in_14_0_7        ), //i
    .port_state_in_14_1_0  (port_state_in_14_1_0        ), //i
    .port_state_in_14_1_1  (port_state_in_14_1_1        ), //i
    .port_state_in_14_1_2  (port_state_in_14_1_2        ), //i
    .port_state_in_14_1_3  (port_state_in_14_1_3        ), //i
    .port_state_in_14_1_4  (port_state_in_14_1_4        ), //i
    .port_state_in_14_1_5  (port_state_in_14_1_5        ), //i
    .port_state_in_14_1_6  (port_state_in_14_1_6        ), //i
    .port_state_in_14_1_7  (port_state_in_14_1_7        ), //i
    .port_state_in_14_2_0  (port_state_in_14_2_0        ), //i
    .port_state_in_14_2_1  (port_state_in_14_2_1        ), //i
    .port_state_in_14_2_2  (port_state_in_14_2_2        ), //i
    .port_state_in_14_2_3  (port_state_in_14_2_3        ), //i
    .port_state_in_14_2_4  (port_state_in_14_2_4        ), //i
    .port_state_in_14_2_5  (port_state_in_14_2_5        ), //i
    .port_state_in_14_2_6  (port_state_in_14_2_6        ), //i
    .port_state_in_14_2_7  (port_state_in_14_2_7        ), //i
    .port_state_in_14_3_0  (port_state_in_14_3_0        ), //i
    .port_state_in_14_3_1  (port_state_in_14_3_1        ), //i
    .port_state_in_14_3_2  (port_state_in_14_3_2        ), //i
    .port_state_in_14_3_3  (port_state_in_14_3_3        ), //i
    .port_state_in_14_3_4  (port_state_in_14_3_4        ), //i
    .port_state_in_14_3_5  (port_state_in_14_3_5        ), //i
    .port_state_in_14_3_6  (port_state_in_14_3_6        ), //i
    .port_state_in_14_3_7  (port_state_in_14_3_7        ), //i
    .port_state_in_15_0_0  (port_state_in_15_0_0        ), //i
    .port_state_in_15_0_1  (port_state_in_15_0_1        ), //i
    .port_state_in_15_0_2  (port_state_in_15_0_2        ), //i
    .port_state_in_15_0_3  (port_state_in_15_0_3        ), //i
    .port_state_in_15_0_4  (port_state_in_15_0_4        ), //i
    .port_state_in_15_0_5  (port_state_in_15_0_5        ), //i
    .port_state_in_15_0_6  (port_state_in_15_0_6        ), //i
    .port_state_in_15_0_7  (port_state_in_15_0_7        ), //i
    .port_state_in_15_1_0  (port_state_in_15_1_0        ), //i
    .port_state_in_15_1_1  (port_state_in_15_1_1        ), //i
    .port_state_in_15_1_2  (port_state_in_15_1_2        ), //i
    .port_state_in_15_1_3  (port_state_in_15_1_3        ), //i
    .port_state_in_15_1_4  (port_state_in_15_1_4        ), //i
    .port_state_in_15_1_5  (port_state_in_15_1_5        ), //i
    .port_state_in_15_1_6  (port_state_in_15_1_6        ), //i
    .port_state_in_15_1_7  (port_state_in_15_1_7        ), //i
    .port_state_in_15_2_0  (port_state_in_15_2_0        ), //i
    .port_state_in_15_2_1  (port_state_in_15_2_1        ), //i
    .port_state_in_15_2_2  (port_state_in_15_2_2        ), //i
    .port_state_in_15_2_3  (port_state_in_15_2_3        ), //i
    .port_state_in_15_2_4  (port_state_in_15_2_4        ), //i
    .port_state_in_15_2_5  (port_state_in_15_2_5        ), //i
    .port_state_in_15_2_6  (port_state_in_15_2_6        ), //i
    .port_state_in_15_2_7  (port_state_in_15_2_7        ), //i
    .port_state_in_15_3_0  (port_state_in_15_3_0        ), //i
    .port_state_in_15_3_1  (port_state_in_15_3_1        ), //i
    .port_state_in_15_3_2  (port_state_in_15_3_2        ), //i
    .port_state_in_15_3_3  (port_state_in_15_3_3        ), //i
    .port_state_in_15_3_4  (port_state_in_15_3_4        ), //i
    .port_state_in_15_3_5  (port_state_in_15_3_5        ), //i
    .port_state_in_15_3_6  (port_state_in_15_3_6        ), //i
    .port_state_in_15_3_7  (port_state_in_15_3_7        ), //i
    .port_key_0_0_0        (port_key_0_0_0              ), //i
    .port_key_0_0_1        (port_key_0_0_1              ), //i
    .port_key_0_0_2        (port_key_0_0_2              ), //i
    .port_key_0_0_3        (port_key_0_0_3              ), //i
    .port_key_0_0_4        (port_key_0_0_4              ), //i
    .port_key_0_0_5        (port_key_0_0_5              ), //i
    .port_key_0_0_6        (port_key_0_0_6              ), //i
    .port_key_0_0_7        (port_key_0_0_7              ), //i
    .port_key_0_1_0        (port_key_0_1_0              ), //i
    .port_key_0_1_1        (port_key_0_1_1              ), //i
    .port_key_0_1_2        (port_key_0_1_2              ), //i
    .port_key_0_1_3        (port_key_0_1_3              ), //i
    .port_key_0_1_4        (port_key_0_1_4              ), //i
    .port_key_0_1_5        (port_key_0_1_5              ), //i
    .port_key_0_1_6        (port_key_0_1_6              ), //i
    .port_key_0_1_7        (port_key_0_1_7              ), //i
    .port_key_0_2_0        (port_key_0_2_0              ), //i
    .port_key_0_2_1        (port_key_0_2_1              ), //i
    .port_key_0_2_2        (port_key_0_2_2              ), //i
    .port_key_0_2_3        (port_key_0_2_3              ), //i
    .port_key_0_2_4        (port_key_0_2_4              ), //i
    .port_key_0_2_5        (port_key_0_2_5              ), //i
    .port_key_0_2_6        (port_key_0_2_6              ), //i
    .port_key_0_2_7        (port_key_0_2_7              ), //i
    .port_key_0_3_0        (port_key_0_3_0              ), //i
    .port_key_0_3_1        (port_key_0_3_1              ), //i
    .port_key_0_3_2        (port_key_0_3_2              ), //i
    .port_key_0_3_3        (port_key_0_3_3              ), //i
    .port_key_0_3_4        (port_key_0_3_4              ), //i
    .port_key_0_3_5        (port_key_0_3_5              ), //i
    .port_key_0_3_6        (port_key_0_3_6              ), //i
    .port_key_0_3_7        (port_key_0_3_7              ), //i
    .port_key_1_0_0        (port_key_1_0_0              ), //i
    .port_key_1_0_1        (port_key_1_0_1              ), //i
    .port_key_1_0_2        (port_key_1_0_2              ), //i
    .port_key_1_0_3        (port_key_1_0_3              ), //i
    .port_key_1_0_4        (port_key_1_0_4              ), //i
    .port_key_1_0_5        (port_key_1_0_5              ), //i
    .port_key_1_0_6        (port_key_1_0_6              ), //i
    .port_key_1_0_7        (port_key_1_0_7              ), //i
    .port_key_1_1_0        (port_key_1_1_0              ), //i
    .port_key_1_1_1        (port_key_1_1_1              ), //i
    .port_key_1_1_2        (port_key_1_1_2              ), //i
    .port_key_1_1_3        (port_key_1_1_3              ), //i
    .port_key_1_1_4        (port_key_1_1_4              ), //i
    .port_key_1_1_5        (port_key_1_1_5              ), //i
    .port_key_1_1_6        (port_key_1_1_6              ), //i
    .port_key_1_1_7        (port_key_1_1_7              ), //i
    .port_key_1_2_0        (port_key_1_2_0              ), //i
    .port_key_1_2_1        (port_key_1_2_1              ), //i
    .port_key_1_2_2        (port_key_1_2_2              ), //i
    .port_key_1_2_3        (port_key_1_2_3              ), //i
    .port_key_1_2_4        (port_key_1_2_4              ), //i
    .port_key_1_2_5        (port_key_1_2_5              ), //i
    .port_key_1_2_6        (port_key_1_2_6              ), //i
    .port_key_1_2_7        (port_key_1_2_7              ), //i
    .port_key_1_3_0        (port_key_1_3_0              ), //i
    .port_key_1_3_1        (port_key_1_3_1              ), //i
    .port_key_1_3_2        (port_key_1_3_2              ), //i
    .port_key_1_3_3        (port_key_1_3_3              ), //i
    .port_key_1_3_4        (port_key_1_3_4              ), //i
    .port_key_1_3_5        (port_key_1_3_5              ), //i
    .port_key_1_3_6        (port_key_1_3_6              ), //i
    .port_key_1_3_7        (port_key_1_3_7              ), //i
    .port_key_2_0_0        (port_key_2_0_0              ), //i
    .port_key_2_0_1        (port_key_2_0_1              ), //i
    .port_key_2_0_2        (port_key_2_0_2              ), //i
    .port_key_2_0_3        (port_key_2_0_3              ), //i
    .port_key_2_0_4        (port_key_2_0_4              ), //i
    .port_key_2_0_5        (port_key_2_0_5              ), //i
    .port_key_2_0_6        (port_key_2_0_6              ), //i
    .port_key_2_0_7        (port_key_2_0_7              ), //i
    .port_key_2_1_0        (port_key_2_1_0              ), //i
    .port_key_2_1_1        (port_key_2_1_1              ), //i
    .port_key_2_1_2        (port_key_2_1_2              ), //i
    .port_key_2_1_3        (port_key_2_1_3              ), //i
    .port_key_2_1_4        (port_key_2_1_4              ), //i
    .port_key_2_1_5        (port_key_2_1_5              ), //i
    .port_key_2_1_6        (port_key_2_1_6              ), //i
    .port_key_2_1_7        (port_key_2_1_7              ), //i
    .port_key_2_2_0        (port_key_2_2_0              ), //i
    .port_key_2_2_1        (port_key_2_2_1              ), //i
    .port_key_2_2_2        (port_key_2_2_2              ), //i
    .port_key_2_2_3        (port_key_2_2_3              ), //i
    .port_key_2_2_4        (port_key_2_2_4              ), //i
    .port_key_2_2_5        (port_key_2_2_5              ), //i
    .port_key_2_2_6        (port_key_2_2_6              ), //i
    .port_key_2_2_7        (port_key_2_2_7              ), //i
    .port_key_2_3_0        (port_key_2_3_0              ), //i
    .port_key_2_3_1        (port_key_2_3_1              ), //i
    .port_key_2_3_2        (port_key_2_3_2              ), //i
    .port_key_2_3_3        (port_key_2_3_3              ), //i
    .port_key_2_3_4        (port_key_2_3_4              ), //i
    .port_key_2_3_5        (port_key_2_3_5              ), //i
    .port_key_2_3_6        (port_key_2_3_6              ), //i
    .port_key_2_3_7        (port_key_2_3_7              ), //i
    .port_key_3_0_0        (port_key_3_0_0              ), //i
    .port_key_3_0_1        (port_key_3_0_1              ), //i
    .port_key_3_0_2        (port_key_3_0_2              ), //i
    .port_key_3_0_3        (port_key_3_0_3              ), //i
    .port_key_3_0_4        (port_key_3_0_4              ), //i
    .port_key_3_0_5        (port_key_3_0_5              ), //i
    .port_key_3_0_6        (port_key_3_0_6              ), //i
    .port_key_3_0_7        (port_key_3_0_7              ), //i
    .port_key_3_1_0        (port_key_3_1_0              ), //i
    .port_key_3_1_1        (port_key_3_1_1              ), //i
    .port_key_3_1_2        (port_key_3_1_2              ), //i
    .port_key_3_1_3        (port_key_3_1_3              ), //i
    .port_key_3_1_4        (port_key_3_1_4              ), //i
    .port_key_3_1_5        (port_key_3_1_5              ), //i
    .port_key_3_1_6        (port_key_3_1_6              ), //i
    .port_key_3_1_7        (port_key_3_1_7              ), //i
    .port_key_3_2_0        (port_key_3_2_0              ), //i
    .port_key_3_2_1        (port_key_3_2_1              ), //i
    .port_key_3_2_2        (port_key_3_2_2              ), //i
    .port_key_3_2_3        (port_key_3_2_3              ), //i
    .port_key_3_2_4        (port_key_3_2_4              ), //i
    .port_key_3_2_5        (port_key_3_2_5              ), //i
    .port_key_3_2_6        (port_key_3_2_6              ), //i
    .port_key_3_2_7        (port_key_3_2_7              ), //i
    .port_key_3_3_0        (port_key_3_3_0              ), //i
    .port_key_3_3_1        (port_key_3_3_1              ), //i
    .port_key_3_3_2        (port_key_3_3_2              ), //i
    .port_key_3_3_3        (port_key_3_3_3              ), //i
    .port_key_3_3_4        (port_key_3_3_4              ), //i
    .port_key_3_3_5        (port_key_3_3_5              ), //i
    .port_key_3_3_6        (port_key_3_3_6              ), //i
    .port_key_3_3_7        (port_key_3_3_7              ), //i
    .port_key_4_0_0        (port_key_4_0_0              ), //i
    .port_key_4_0_1        (port_key_4_0_1              ), //i
    .port_key_4_0_2        (port_key_4_0_2              ), //i
    .port_key_4_0_3        (port_key_4_0_3              ), //i
    .port_key_4_0_4        (port_key_4_0_4              ), //i
    .port_key_4_0_5        (port_key_4_0_5              ), //i
    .port_key_4_0_6        (port_key_4_0_6              ), //i
    .port_key_4_0_7        (port_key_4_0_7              ), //i
    .port_key_4_1_0        (port_key_4_1_0              ), //i
    .port_key_4_1_1        (port_key_4_1_1              ), //i
    .port_key_4_1_2        (port_key_4_1_2              ), //i
    .port_key_4_1_3        (port_key_4_1_3              ), //i
    .port_key_4_1_4        (port_key_4_1_4              ), //i
    .port_key_4_1_5        (port_key_4_1_5              ), //i
    .port_key_4_1_6        (port_key_4_1_6              ), //i
    .port_key_4_1_7        (port_key_4_1_7              ), //i
    .port_key_4_2_0        (port_key_4_2_0              ), //i
    .port_key_4_2_1        (port_key_4_2_1              ), //i
    .port_key_4_2_2        (port_key_4_2_2              ), //i
    .port_key_4_2_3        (port_key_4_2_3              ), //i
    .port_key_4_2_4        (port_key_4_2_4              ), //i
    .port_key_4_2_5        (port_key_4_2_5              ), //i
    .port_key_4_2_6        (port_key_4_2_6              ), //i
    .port_key_4_2_7        (port_key_4_2_7              ), //i
    .port_key_4_3_0        (port_key_4_3_0              ), //i
    .port_key_4_3_1        (port_key_4_3_1              ), //i
    .port_key_4_3_2        (port_key_4_3_2              ), //i
    .port_key_4_3_3        (port_key_4_3_3              ), //i
    .port_key_4_3_4        (port_key_4_3_4              ), //i
    .port_key_4_3_5        (port_key_4_3_5              ), //i
    .port_key_4_3_6        (port_key_4_3_6              ), //i
    .port_key_4_3_7        (port_key_4_3_7              ), //i
    .port_key_5_0_0        (port_key_5_0_0              ), //i
    .port_key_5_0_1        (port_key_5_0_1              ), //i
    .port_key_5_0_2        (port_key_5_0_2              ), //i
    .port_key_5_0_3        (port_key_5_0_3              ), //i
    .port_key_5_0_4        (port_key_5_0_4              ), //i
    .port_key_5_0_5        (port_key_5_0_5              ), //i
    .port_key_5_0_6        (port_key_5_0_6              ), //i
    .port_key_5_0_7        (port_key_5_0_7              ), //i
    .port_key_5_1_0        (port_key_5_1_0              ), //i
    .port_key_5_1_1        (port_key_5_1_1              ), //i
    .port_key_5_1_2        (port_key_5_1_2              ), //i
    .port_key_5_1_3        (port_key_5_1_3              ), //i
    .port_key_5_1_4        (port_key_5_1_4              ), //i
    .port_key_5_1_5        (port_key_5_1_5              ), //i
    .port_key_5_1_6        (port_key_5_1_6              ), //i
    .port_key_5_1_7        (port_key_5_1_7              ), //i
    .port_key_5_2_0        (port_key_5_2_0              ), //i
    .port_key_5_2_1        (port_key_5_2_1              ), //i
    .port_key_5_2_2        (port_key_5_2_2              ), //i
    .port_key_5_2_3        (port_key_5_2_3              ), //i
    .port_key_5_2_4        (port_key_5_2_4              ), //i
    .port_key_5_2_5        (port_key_5_2_5              ), //i
    .port_key_5_2_6        (port_key_5_2_6              ), //i
    .port_key_5_2_7        (port_key_5_2_7              ), //i
    .port_key_5_3_0        (port_key_5_3_0              ), //i
    .port_key_5_3_1        (port_key_5_3_1              ), //i
    .port_key_5_3_2        (port_key_5_3_2              ), //i
    .port_key_5_3_3        (port_key_5_3_3              ), //i
    .port_key_5_3_4        (port_key_5_3_4              ), //i
    .port_key_5_3_5        (port_key_5_3_5              ), //i
    .port_key_5_3_6        (port_key_5_3_6              ), //i
    .port_key_5_3_7        (port_key_5_3_7              ), //i
    .port_key_6_0_0        (port_key_6_0_0              ), //i
    .port_key_6_0_1        (port_key_6_0_1              ), //i
    .port_key_6_0_2        (port_key_6_0_2              ), //i
    .port_key_6_0_3        (port_key_6_0_3              ), //i
    .port_key_6_0_4        (port_key_6_0_4              ), //i
    .port_key_6_0_5        (port_key_6_0_5              ), //i
    .port_key_6_0_6        (port_key_6_0_6              ), //i
    .port_key_6_0_7        (port_key_6_0_7              ), //i
    .port_key_6_1_0        (port_key_6_1_0              ), //i
    .port_key_6_1_1        (port_key_6_1_1              ), //i
    .port_key_6_1_2        (port_key_6_1_2              ), //i
    .port_key_6_1_3        (port_key_6_1_3              ), //i
    .port_key_6_1_4        (port_key_6_1_4              ), //i
    .port_key_6_1_5        (port_key_6_1_5              ), //i
    .port_key_6_1_6        (port_key_6_1_6              ), //i
    .port_key_6_1_7        (port_key_6_1_7              ), //i
    .port_key_6_2_0        (port_key_6_2_0              ), //i
    .port_key_6_2_1        (port_key_6_2_1              ), //i
    .port_key_6_2_2        (port_key_6_2_2              ), //i
    .port_key_6_2_3        (port_key_6_2_3              ), //i
    .port_key_6_2_4        (port_key_6_2_4              ), //i
    .port_key_6_2_5        (port_key_6_2_5              ), //i
    .port_key_6_2_6        (port_key_6_2_6              ), //i
    .port_key_6_2_7        (port_key_6_2_7              ), //i
    .port_key_6_3_0        (port_key_6_3_0              ), //i
    .port_key_6_3_1        (port_key_6_3_1              ), //i
    .port_key_6_3_2        (port_key_6_3_2              ), //i
    .port_key_6_3_3        (port_key_6_3_3              ), //i
    .port_key_6_3_4        (port_key_6_3_4              ), //i
    .port_key_6_3_5        (port_key_6_3_5              ), //i
    .port_key_6_3_6        (port_key_6_3_6              ), //i
    .port_key_6_3_7        (port_key_6_3_7              ), //i
    .port_key_7_0_0        (port_key_7_0_0              ), //i
    .port_key_7_0_1        (port_key_7_0_1              ), //i
    .port_key_7_0_2        (port_key_7_0_2              ), //i
    .port_key_7_0_3        (port_key_7_0_3              ), //i
    .port_key_7_0_4        (port_key_7_0_4              ), //i
    .port_key_7_0_5        (port_key_7_0_5              ), //i
    .port_key_7_0_6        (port_key_7_0_6              ), //i
    .port_key_7_0_7        (port_key_7_0_7              ), //i
    .port_key_7_1_0        (port_key_7_1_0              ), //i
    .port_key_7_1_1        (port_key_7_1_1              ), //i
    .port_key_7_1_2        (port_key_7_1_2              ), //i
    .port_key_7_1_3        (port_key_7_1_3              ), //i
    .port_key_7_1_4        (port_key_7_1_4              ), //i
    .port_key_7_1_5        (port_key_7_1_5              ), //i
    .port_key_7_1_6        (port_key_7_1_6              ), //i
    .port_key_7_1_7        (port_key_7_1_7              ), //i
    .port_key_7_2_0        (port_key_7_2_0              ), //i
    .port_key_7_2_1        (port_key_7_2_1              ), //i
    .port_key_7_2_2        (port_key_7_2_2              ), //i
    .port_key_7_2_3        (port_key_7_2_3              ), //i
    .port_key_7_2_4        (port_key_7_2_4              ), //i
    .port_key_7_2_5        (port_key_7_2_5              ), //i
    .port_key_7_2_6        (port_key_7_2_6              ), //i
    .port_key_7_2_7        (port_key_7_2_7              ), //i
    .port_key_7_3_0        (port_key_7_3_0              ), //i
    .port_key_7_3_1        (port_key_7_3_1              ), //i
    .port_key_7_3_2        (port_key_7_3_2              ), //i
    .port_key_7_3_3        (port_key_7_3_3              ), //i
    .port_key_7_3_4        (port_key_7_3_4              ), //i
    .port_key_7_3_5        (port_key_7_3_5              ), //i
    .port_key_7_3_6        (port_key_7_3_6              ), //i
    .port_key_7_3_7        (port_key_7_3_7              ), //i
    .port_key_8_0_0        (port_key_8_0_0              ), //i
    .port_key_8_0_1        (port_key_8_0_1              ), //i
    .port_key_8_0_2        (port_key_8_0_2              ), //i
    .port_key_8_0_3        (port_key_8_0_3              ), //i
    .port_key_8_0_4        (port_key_8_0_4              ), //i
    .port_key_8_0_5        (port_key_8_0_5              ), //i
    .port_key_8_0_6        (port_key_8_0_6              ), //i
    .port_key_8_0_7        (port_key_8_0_7              ), //i
    .port_key_8_1_0        (port_key_8_1_0              ), //i
    .port_key_8_1_1        (port_key_8_1_1              ), //i
    .port_key_8_1_2        (port_key_8_1_2              ), //i
    .port_key_8_1_3        (port_key_8_1_3              ), //i
    .port_key_8_1_4        (port_key_8_1_4              ), //i
    .port_key_8_1_5        (port_key_8_1_5              ), //i
    .port_key_8_1_6        (port_key_8_1_6              ), //i
    .port_key_8_1_7        (port_key_8_1_7              ), //i
    .port_key_8_2_0        (port_key_8_2_0              ), //i
    .port_key_8_2_1        (port_key_8_2_1              ), //i
    .port_key_8_2_2        (port_key_8_2_2              ), //i
    .port_key_8_2_3        (port_key_8_2_3              ), //i
    .port_key_8_2_4        (port_key_8_2_4              ), //i
    .port_key_8_2_5        (port_key_8_2_5              ), //i
    .port_key_8_2_6        (port_key_8_2_6              ), //i
    .port_key_8_2_7        (port_key_8_2_7              ), //i
    .port_key_8_3_0        (port_key_8_3_0              ), //i
    .port_key_8_3_1        (port_key_8_3_1              ), //i
    .port_key_8_3_2        (port_key_8_3_2              ), //i
    .port_key_8_3_3        (port_key_8_3_3              ), //i
    .port_key_8_3_4        (port_key_8_3_4              ), //i
    .port_key_8_3_5        (port_key_8_3_5              ), //i
    .port_key_8_3_6        (port_key_8_3_6              ), //i
    .port_key_8_3_7        (port_key_8_3_7              ), //i
    .port_key_9_0_0        (port_key_9_0_0              ), //i
    .port_key_9_0_1        (port_key_9_0_1              ), //i
    .port_key_9_0_2        (port_key_9_0_2              ), //i
    .port_key_9_0_3        (port_key_9_0_3              ), //i
    .port_key_9_0_4        (port_key_9_0_4              ), //i
    .port_key_9_0_5        (port_key_9_0_5              ), //i
    .port_key_9_0_6        (port_key_9_0_6              ), //i
    .port_key_9_0_7        (port_key_9_0_7              ), //i
    .port_key_9_1_0        (port_key_9_1_0              ), //i
    .port_key_9_1_1        (port_key_9_1_1              ), //i
    .port_key_9_1_2        (port_key_9_1_2              ), //i
    .port_key_9_1_3        (port_key_9_1_3              ), //i
    .port_key_9_1_4        (port_key_9_1_4              ), //i
    .port_key_9_1_5        (port_key_9_1_5              ), //i
    .port_key_9_1_6        (port_key_9_1_6              ), //i
    .port_key_9_1_7        (port_key_9_1_7              ), //i
    .port_key_9_2_0        (port_key_9_2_0              ), //i
    .port_key_9_2_1        (port_key_9_2_1              ), //i
    .port_key_9_2_2        (port_key_9_2_2              ), //i
    .port_key_9_2_3        (port_key_9_2_3              ), //i
    .port_key_9_2_4        (port_key_9_2_4              ), //i
    .port_key_9_2_5        (port_key_9_2_5              ), //i
    .port_key_9_2_6        (port_key_9_2_6              ), //i
    .port_key_9_2_7        (port_key_9_2_7              ), //i
    .port_key_9_3_0        (port_key_9_3_0              ), //i
    .port_key_9_3_1        (port_key_9_3_1              ), //i
    .port_key_9_3_2        (port_key_9_3_2              ), //i
    .port_key_9_3_3        (port_key_9_3_3              ), //i
    .port_key_9_3_4        (port_key_9_3_4              ), //i
    .port_key_9_3_5        (port_key_9_3_5              ), //i
    .port_key_9_3_6        (port_key_9_3_6              ), //i
    .port_key_9_3_7        (port_key_9_3_7              ), //i
    .port_key_10_0_0       (port_key_10_0_0             ), //i
    .port_key_10_0_1       (port_key_10_0_1             ), //i
    .port_key_10_0_2       (port_key_10_0_2             ), //i
    .port_key_10_0_3       (port_key_10_0_3             ), //i
    .port_key_10_0_4       (port_key_10_0_4             ), //i
    .port_key_10_0_5       (port_key_10_0_5             ), //i
    .port_key_10_0_6       (port_key_10_0_6             ), //i
    .port_key_10_0_7       (port_key_10_0_7             ), //i
    .port_key_10_1_0       (port_key_10_1_0             ), //i
    .port_key_10_1_1       (port_key_10_1_1             ), //i
    .port_key_10_1_2       (port_key_10_1_2             ), //i
    .port_key_10_1_3       (port_key_10_1_3             ), //i
    .port_key_10_1_4       (port_key_10_1_4             ), //i
    .port_key_10_1_5       (port_key_10_1_5             ), //i
    .port_key_10_1_6       (port_key_10_1_6             ), //i
    .port_key_10_1_7       (port_key_10_1_7             ), //i
    .port_key_10_2_0       (port_key_10_2_0             ), //i
    .port_key_10_2_1       (port_key_10_2_1             ), //i
    .port_key_10_2_2       (port_key_10_2_2             ), //i
    .port_key_10_2_3       (port_key_10_2_3             ), //i
    .port_key_10_2_4       (port_key_10_2_4             ), //i
    .port_key_10_2_5       (port_key_10_2_5             ), //i
    .port_key_10_2_6       (port_key_10_2_6             ), //i
    .port_key_10_2_7       (port_key_10_2_7             ), //i
    .port_key_10_3_0       (port_key_10_3_0             ), //i
    .port_key_10_3_1       (port_key_10_3_1             ), //i
    .port_key_10_3_2       (port_key_10_3_2             ), //i
    .port_key_10_3_3       (port_key_10_3_3             ), //i
    .port_key_10_3_4       (port_key_10_3_4             ), //i
    .port_key_10_3_5       (port_key_10_3_5             ), //i
    .port_key_10_3_6       (port_key_10_3_6             ), //i
    .port_key_10_3_7       (port_key_10_3_7             ), //i
    .port_key_11_0_0       (port_key_11_0_0             ), //i
    .port_key_11_0_1       (port_key_11_0_1             ), //i
    .port_key_11_0_2       (port_key_11_0_2             ), //i
    .port_key_11_0_3       (port_key_11_0_3             ), //i
    .port_key_11_0_4       (port_key_11_0_4             ), //i
    .port_key_11_0_5       (port_key_11_0_5             ), //i
    .port_key_11_0_6       (port_key_11_0_6             ), //i
    .port_key_11_0_7       (port_key_11_0_7             ), //i
    .port_key_11_1_0       (port_key_11_1_0             ), //i
    .port_key_11_1_1       (port_key_11_1_1             ), //i
    .port_key_11_1_2       (port_key_11_1_2             ), //i
    .port_key_11_1_3       (port_key_11_1_3             ), //i
    .port_key_11_1_4       (port_key_11_1_4             ), //i
    .port_key_11_1_5       (port_key_11_1_5             ), //i
    .port_key_11_1_6       (port_key_11_1_6             ), //i
    .port_key_11_1_7       (port_key_11_1_7             ), //i
    .port_key_11_2_0       (port_key_11_2_0             ), //i
    .port_key_11_2_1       (port_key_11_2_1             ), //i
    .port_key_11_2_2       (port_key_11_2_2             ), //i
    .port_key_11_2_3       (port_key_11_2_3             ), //i
    .port_key_11_2_4       (port_key_11_2_4             ), //i
    .port_key_11_2_5       (port_key_11_2_5             ), //i
    .port_key_11_2_6       (port_key_11_2_6             ), //i
    .port_key_11_2_7       (port_key_11_2_7             ), //i
    .port_key_11_3_0       (port_key_11_3_0             ), //i
    .port_key_11_3_1       (port_key_11_3_1             ), //i
    .port_key_11_3_2       (port_key_11_3_2             ), //i
    .port_key_11_3_3       (port_key_11_3_3             ), //i
    .port_key_11_3_4       (port_key_11_3_4             ), //i
    .port_key_11_3_5       (port_key_11_3_5             ), //i
    .port_key_11_3_6       (port_key_11_3_6             ), //i
    .port_key_11_3_7       (port_key_11_3_7             ), //i
    .port_key_12_0_0       (port_key_12_0_0             ), //i
    .port_key_12_0_1       (port_key_12_0_1             ), //i
    .port_key_12_0_2       (port_key_12_0_2             ), //i
    .port_key_12_0_3       (port_key_12_0_3             ), //i
    .port_key_12_0_4       (port_key_12_0_4             ), //i
    .port_key_12_0_5       (port_key_12_0_5             ), //i
    .port_key_12_0_6       (port_key_12_0_6             ), //i
    .port_key_12_0_7       (port_key_12_0_7             ), //i
    .port_key_12_1_0       (port_key_12_1_0             ), //i
    .port_key_12_1_1       (port_key_12_1_1             ), //i
    .port_key_12_1_2       (port_key_12_1_2             ), //i
    .port_key_12_1_3       (port_key_12_1_3             ), //i
    .port_key_12_1_4       (port_key_12_1_4             ), //i
    .port_key_12_1_5       (port_key_12_1_5             ), //i
    .port_key_12_1_6       (port_key_12_1_6             ), //i
    .port_key_12_1_7       (port_key_12_1_7             ), //i
    .port_key_12_2_0       (port_key_12_2_0             ), //i
    .port_key_12_2_1       (port_key_12_2_1             ), //i
    .port_key_12_2_2       (port_key_12_2_2             ), //i
    .port_key_12_2_3       (port_key_12_2_3             ), //i
    .port_key_12_2_4       (port_key_12_2_4             ), //i
    .port_key_12_2_5       (port_key_12_2_5             ), //i
    .port_key_12_2_6       (port_key_12_2_6             ), //i
    .port_key_12_2_7       (port_key_12_2_7             ), //i
    .port_key_12_3_0       (port_key_12_3_0             ), //i
    .port_key_12_3_1       (port_key_12_3_1             ), //i
    .port_key_12_3_2       (port_key_12_3_2             ), //i
    .port_key_12_3_3       (port_key_12_3_3             ), //i
    .port_key_12_3_4       (port_key_12_3_4             ), //i
    .port_key_12_3_5       (port_key_12_3_5             ), //i
    .port_key_12_3_6       (port_key_12_3_6             ), //i
    .port_key_12_3_7       (port_key_12_3_7             ), //i
    .port_key_13_0_0       (port_key_13_0_0             ), //i
    .port_key_13_0_1       (port_key_13_0_1             ), //i
    .port_key_13_0_2       (port_key_13_0_2             ), //i
    .port_key_13_0_3       (port_key_13_0_3             ), //i
    .port_key_13_0_4       (port_key_13_0_4             ), //i
    .port_key_13_0_5       (port_key_13_0_5             ), //i
    .port_key_13_0_6       (port_key_13_0_6             ), //i
    .port_key_13_0_7       (port_key_13_0_7             ), //i
    .port_key_13_1_0       (port_key_13_1_0             ), //i
    .port_key_13_1_1       (port_key_13_1_1             ), //i
    .port_key_13_1_2       (port_key_13_1_2             ), //i
    .port_key_13_1_3       (port_key_13_1_3             ), //i
    .port_key_13_1_4       (port_key_13_1_4             ), //i
    .port_key_13_1_5       (port_key_13_1_5             ), //i
    .port_key_13_1_6       (port_key_13_1_6             ), //i
    .port_key_13_1_7       (port_key_13_1_7             ), //i
    .port_key_13_2_0       (port_key_13_2_0             ), //i
    .port_key_13_2_1       (port_key_13_2_1             ), //i
    .port_key_13_2_2       (port_key_13_2_2             ), //i
    .port_key_13_2_3       (port_key_13_2_3             ), //i
    .port_key_13_2_4       (port_key_13_2_4             ), //i
    .port_key_13_2_5       (port_key_13_2_5             ), //i
    .port_key_13_2_6       (port_key_13_2_6             ), //i
    .port_key_13_2_7       (port_key_13_2_7             ), //i
    .port_key_13_3_0       (port_key_13_3_0             ), //i
    .port_key_13_3_1       (port_key_13_3_1             ), //i
    .port_key_13_3_2       (port_key_13_3_2             ), //i
    .port_key_13_3_3       (port_key_13_3_3             ), //i
    .port_key_13_3_4       (port_key_13_3_4             ), //i
    .port_key_13_3_5       (port_key_13_3_5             ), //i
    .port_key_13_3_6       (port_key_13_3_6             ), //i
    .port_key_13_3_7       (port_key_13_3_7             ), //i
    .port_key_14_0_0       (port_key_14_0_0             ), //i
    .port_key_14_0_1       (port_key_14_0_1             ), //i
    .port_key_14_0_2       (port_key_14_0_2             ), //i
    .port_key_14_0_3       (port_key_14_0_3             ), //i
    .port_key_14_0_4       (port_key_14_0_4             ), //i
    .port_key_14_0_5       (port_key_14_0_5             ), //i
    .port_key_14_0_6       (port_key_14_0_6             ), //i
    .port_key_14_0_7       (port_key_14_0_7             ), //i
    .port_key_14_1_0       (port_key_14_1_0             ), //i
    .port_key_14_1_1       (port_key_14_1_1             ), //i
    .port_key_14_1_2       (port_key_14_1_2             ), //i
    .port_key_14_1_3       (port_key_14_1_3             ), //i
    .port_key_14_1_4       (port_key_14_1_4             ), //i
    .port_key_14_1_5       (port_key_14_1_5             ), //i
    .port_key_14_1_6       (port_key_14_1_6             ), //i
    .port_key_14_1_7       (port_key_14_1_7             ), //i
    .port_key_14_2_0       (port_key_14_2_0             ), //i
    .port_key_14_2_1       (port_key_14_2_1             ), //i
    .port_key_14_2_2       (port_key_14_2_2             ), //i
    .port_key_14_2_3       (port_key_14_2_3             ), //i
    .port_key_14_2_4       (port_key_14_2_4             ), //i
    .port_key_14_2_5       (port_key_14_2_5             ), //i
    .port_key_14_2_6       (port_key_14_2_6             ), //i
    .port_key_14_2_7       (port_key_14_2_7             ), //i
    .port_key_14_3_0       (port_key_14_3_0             ), //i
    .port_key_14_3_1       (port_key_14_3_1             ), //i
    .port_key_14_3_2       (port_key_14_3_2             ), //i
    .port_key_14_3_3       (port_key_14_3_3             ), //i
    .port_key_14_3_4       (port_key_14_3_4             ), //i
    .port_key_14_3_5       (port_key_14_3_5             ), //i
    .port_key_14_3_6       (port_key_14_3_6             ), //i
    .port_key_14_3_7       (port_key_14_3_7             ), //i
    .port_key_15_0_0       (port_key_15_0_0             ), //i
    .port_key_15_0_1       (port_key_15_0_1             ), //i
    .port_key_15_0_2       (port_key_15_0_2             ), //i
    .port_key_15_0_3       (port_key_15_0_3             ), //i
    .port_key_15_0_4       (port_key_15_0_4             ), //i
    .port_key_15_0_5       (port_key_15_0_5             ), //i
    .port_key_15_0_6       (port_key_15_0_6             ), //i
    .port_key_15_0_7       (port_key_15_0_7             ), //i
    .port_key_15_1_0       (port_key_15_1_0             ), //i
    .port_key_15_1_1       (port_key_15_1_1             ), //i
    .port_key_15_1_2       (port_key_15_1_2             ), //i
    .port_key_15_1_3       (port_key_15_1_3             ), //i
    .port_key_15_1_4       (port_key_15_1_4             ), //i
    .port_key_15_1_5       (port_key_15_1_5             ), //i
    .port_key_15_1_6       (port_key_15_1_6             ), //i
    .port_key_15_1_7       (port_key_15_1_7             ), //i
    .port_key_15_2_0       (port_key_15_2_0             ), //i
    .port_key_15_2_1       (port_key_15_2_1             ), //i
    .port_key_15_2_2       (port_key_15_2_2             ), //i
    .port_key_15_2_3       (port_key_15_2_3             ), //i
    .port_key_15_2_4       (port_key_15_2_4             ), //i
    .port_key_15_2_5       (port_key_15_2_5             ), //i
    .port_key_15_2_6       (port_key_15_2_6             ), //i
    .port_key_15_2_7       (port_key_15_2_7             ), //i
    .port_key_15_3_0       (port_key_15_3_0             ), //i
    .port_key_15_3_1       (port_key_15_3_1             ), //i
    .port_key_15_3_2       (port_key_15_3_2             ), //i
    .port_key_15_3_3       (port_key_15_3_3             ), //i
    .port_key_15_3_4       (port_key_15_3_4             ), //i
    .port_key_15_3_5       (port_key_15_3_5             ), //i
    .port_key_15_3_6       (port_key_15_3_6             ), //i
    .port_key_15_3_7       (port_key_15_3_7             ), //i
    .port_state_out_0_0_0  (keyAdd_port_state_out_0_0_0 ), //o
    .port_state_out_0_0_1  (keyAdd_port_state_out_0_0_1 ), //o
    .port_state_out_0_0_2  (keyAdd_port_state_out_0_0_2 ), //o
    .port_state_out_0_0_3  (keyAdd_port_state_out_0_0_3 ), //o
    .port_state_out_0_0_4  (keyAdd_port_state_out_0_0_4 ), //o
    .port_state_out_0_0_5  (keyAdd_port_state_out_0_0_5 ), //o
    .port_state_out_0_0_6  (keyAdd_port_state_out_0_0_6 ), //o
    .port_state_out_0_0_7  (keyAdd_port_state_out_0_0_7 ), //o
    .port_state_out_0_1_0  (keyAdd_port_state_out_0_1_0 ), //o
    .port_state_out_0_1_1  (keyAdd_port_state_out_0_1_1 ), //o
    .port_state_out_0_1_2  (keyAdd_port_state_out_0_1_2 ), //o
    .port_state_out_0_1_3  (keyAdd_port_state_out_0_1_3 ), //o
    .port_state_out_0_1_4  (keyAdd_port_state_out_0_1_4 ), //o
    .port_state_out_0_1_5  (keyAdd_port_state_out_0_1_5 ), //o
    .port_state_out_0_1_6  (keyAdd_port_state_out_0_1_6 ), //o
    .port_state_out_0_1_7  (keyAdd_port_state_out_0_1_7 ), //o
    .port_state_out_0_2_0  (keyAdd_port_state_out_0_2_0 ), //o
    .port_state_out_0_2_1  (keyAdd_port_state_out_0_2_1 ), //o
    .port_state_out_0_2_2  (keyAdd_port_state_out_0_2_2 ), //o
    .port_state_out_0_2_3  (keyAdd_port_state_out_0_2_3 ), //o
    .port_state_out_0_2_4  (keyAdd_port_state_out_0_2_4 ), //o
    .port_state_out_0_2_5  (keyAdd_port_state_out_0_2_5 ), //o
    .port_state_out_0_2_6  (keyAdd_port_state_out_0_2_6 ), //o
    .port_state_out_0_2_7  (keyAdd_port_state_out_0_2_7 ), //o
    .port_state_out_0_3_0  (keyAdd_port_state_out_0_3_0 ), //o
    .port_state_out_0_3_1  (keyAdd_port_state_out_0_3_1 ), //o
    .port_state_out_0_3_2  (keyAdd_port_state_out_0_3_2 ), //o
    .port_state_out_0_3_3  (keyAdd_port_state_out_0_3_3 ), //o
    .port_state_out_0_3_4  (keyAdd_port_state_out_0_3_4 ), //o
    .port_state_out_0_3_5  (keyAdd_port_state_out_0_3_5 ), //o
    .port_state_out_0_3_6  (keyAdd_port_state_out_0_3_6 ), //o
    .port_state_out_0_3_7  (keyAdd_port_state_out_0_3_7 ), //o
    .port_state_out_1_0_0  (keyAdd_port_state_out_1_0_0 ), //o
    .port_state_out_1_0_1  (keyAdd_port_state_out_1_0_1 ), //o
    .port_state_out_1_0_2  (keyAdd_port_state_out_1_0_2 ), //o
    .port_state_out_1_0_3  (keyAdd_port_state_out_1_0_3 ), //o
    .port_state_out_1_0_4  (keyAdd_port_state_out_1_0_4 ), //o
    .port_state_out_1_0_5  (keyAdd_port_state_out_1_0_5 ), //o
    .port_state_out_1_0_6  (keyAdd_port_state_out_1_0_6 ), //o
    .port_state_out_1_0_7  (keyAdd_port_state_out_1_0_7 ), //o
    .port_state_out_1_1_0  (keyAdd_port_state_out_1_1_0 ), //o
    .port_state_out_1_1_1  (keyAdd_port_state_out_1_1_1 ), //o
    .port_state_out_1_1_2  (keyAdd_port_state_out_1_1_2 ), //o
    .port_state_out_1_1_3  (keyAdd_port_state_out_1_1_3 ), //o
    .port_state_out_1_1_4  (keyAdd_port_state_out_1_1_4 ), //o
    .port_state_out_1_1_5  (keyAdd_port_state_out_1_1_5 ), //o
    .port_state_out_1_1_6  (keyAdd_port_state_out_1_1_6 ), //o
    .port_state_out_1_1_7  (keyAdd_port_state_out_1_1_7 ), //o
    .port_state_out_1_2_0  (keyAdd_port_state_out_1_2_0 ), //o
    .port_state_out_1_2_1  (keyAdd_port_state_out_1_2_1 ), //o
    .port_state_out_1_2_2  (keyAdd_port_state_out_1_2_2 ), //o
    .port_state_out_1_2_3  (keyAdd_port_state_out_1_2_3 ), //o
    .port_state_out_1_2_4  (keyAdd_port_state_out_1_2_4 ), //o
    .port_state_out_1_2_5  (keyAdd_port_state_out_1_2_5 ), //o
    .port_state_out_1_2_6  (keyAdd_port_state_out_1_2_6 ), //o
    .port_state_out_1_2_7  (keyAdd_port_state_out_1_2_7 ), //o
    .port_state_out_1_3_0  (keyAdd_port_state_out_1_3_0 ), //o
    .port_state_out_1_3_1  (keyAdd_port_state_out_1_3_1 ), //o
    .port_state_out_1_3_2  (keyAdd_port_state_out_1_3_2 ), //o
    .port_state_out_1_3_3  (keyAdd_port_state_out_1_3_3 ), //o
    .port_state_out_1_3_4  (keyAdd_port_state_out_1_3_4 ), //o
    .port_state_out_1_3_5  (keyAdd_port_state_out_1_3_5 ), //o
    .port_state_out_1_3_6  (keyAdd_port_state_out_1_3_6 ), //o
    .port_state_out_1_3_7  (keyAdd_port_state_out_1_3_7 ), //o
    .port_state_out_2_0_0  (keyAdd_port_state_out_2_0_0 ), //o
    .port_state_out_2_0_1  (keyAdd_port_state_out_2_0_1 ), //o
    .port_state_out_2_0_2  (keyAdd_port_state_out_2_0_2 ), //o
    .port_state_out_2_0_3  (keyAdd_port_state_out_2_0_3 ), //o
    .port_state_out_2_0_4  (keyAdd_port_state_out_2_0_4 ), //o
    .port_state_out_2_0_5  (keyAdd_port_state_out_2_0_5 ), //o
    .port_state_out_2_0_6  (keyAdd_port_state_out_2_0_6 ), //o
    .port_state_out_2_0_7  (keyAdd_port_state_out_2_0_7 ), //o
    .port_state_out_2_1_0  (keyAdd_port_state_out_2_1_0 ), //o
    .port_state_out_2_1_1  (keyAdd_port_state_out_2_1_1 ), //o
    .port_state_out_2_1_2  (keyAdd_port_state_out_2_1_2 ), //o
    .port_state_out_2_1_3  (keyAdd_port_state_out_2_1_3 ), //o
    .port_state_out_2_1_4  (keyAdd_port_state_out_2_1_4 ), //o
    .port_state_out_2_1_5  (keyAdd_port_state_out_2_1_5 ), //o
    .port_state_out_2_1_6  (keyAdd_port_state_out_2_1_6 ), //o
    .port_state_out_2_1_7  (keyAdd_port_state_out_2_1_7 ), //o
    .port_state_out_2_2_0  (keyAdd_port_state_out_2_2_0 ), //o
    .port_state_out_2_2_1  (keyAdd_port_state_out_2_2_1 ), //o
    .port_state_out_2_2_2  (keyAdd_port_state_out_2_2_2 ), //o
    .port_state_out_2_2_3  (keyAdd_port_state_out_2_2_3 ), //o
    .port_state_out_2_2_4  (keyAdd_port_state_out_2_2_4 ), //o
    .port_state_out_2_2_5  (keyAdd_port_state_out_2_2_5 ), //o
    .port_state_out_2_2_6  (keyAdd_port_state_out_2_2_6 ), //o
    .port_state_out_2_2_7  (keyAdd_port_state_out_2_2_7 ), //o
    .port_state_out_2_3_0  (keyAdd_port_state_out_2_3_0 ), //o
    .port_state_out_2_3_1  (keyAdd_port_state_out_2_3_1 ), //o
    .port_state_out_2_3_2  (keyAdd_port_state_out_2_3_2 ), //o
    .port_state_out_2_3_3  (keyAdd_port_state_out_2_3_3 ), //o
    .port_state_out_2_3_4  (keyAdd_port_state_out_2_3_4 ), //o
    .port_state_out_2_3_5  (keyAdd_port_state_out_2_3_5 ), //o
    .port_state_out_2_3_6  (keyAdd_port_state_out_2_3_6 ), //o
    .port_state_out_2_3_7  (keyAdd_port_state_out_2_3_7 ), //o
    .port_state_out_3_0_0  (keyAdd_port_state_out_3_0_0 ), //o
    .port_state_out_3_0_1  (keyAdd_port_state_out_3_0_1 ), //o
    .port_state_out_3_0_2  (keyAdd_port_state_out_3_0_2 ), //o
    .port_state_out_3_0_3  (keyAdd_port_state_out_3_0_3 ), //o
    .port_state_out_3_0_4  (keyAdd_port_state_out_3_0_4 ), //o
    .port_state_out_3_0_5  (keyAdd_port_state_out_3_0_5 ), //o
    .port_state_out_3_0_6  (keyAdd_port_state_out_3_0_6 ), //o
    .port_state_out_3_0_7  (keyAdd_port_state_out_3_0_7 ), //o
    .port_state_out_3_1_0  (keyAdd_port_state_out_3_1_0 ), //o
    .port_state_out_3_1_1  (keyAdd_port_state_out_3_1_1 ), //o
    .port_state_out_3_1_2  (keyAdd_port_state_out_3_1_2 ), //o
    .port_state_out_3_1_3  (keyAdd_port_state_out_3_1_3 ), //o
    .port_state_out_3_1_4  (keyAdd_port_state_out_3_1_4 ), //o
    .port_state_out_3_1_5  (keyAdd_port_state_out_3_1_5 ), //o
    .port_state_out_3_1_6  (keyAdd_port_state_out_3_1_6 ), //o
    .port_state_out_3_1_7  (keyAdd_port_state_out_3_1_7 ), //o
    .port_state_out_3_2_0  (keyAdd_port_state_out_3_2_0 ), //o
    .port_state_out_3_2_1  (keyAdd_port_state_out_3_2_1 ), //o
    .port_state_out_3_2_2  (keyAdd_port_state_out_3_2_2 ), //o
    .port_state_out_3_2_3  (keyAdd_port_state_out_3_2_3 ), //o
    .port_state_out_3_2_4  (keyAdd_port_state_out_3_2_4 ), //o
    .port_state_out_3_2_5  (keyAdd_port_state_out_3_2_5 ), //o
    .port_state_out_3_2_6  (keyAdd_port_state_out_3_2_6 ), //o
    .port_state_out_3_2_7  (keyAdd_port_state_out_3_2_7 ), //o
    .port_state_out_3_3_0  (keyAdd_port_state_out_3_3_0 ), //o
    .port_state_out_3_3_1  (keyAdd_port_state_out_3_3_1 ), //o
    .port_state_out_3_3_2  (keyAdd_port_state_out_3_3_2 ), //o
    .port_state_out_3_3_3  (keyAdd_port_state_out_3_3_3 ), //o
    .port_state_out_3_3_4  (keyAdd_port_state_out_3_3_4 ), //o
    .port_state_out_3_3_5  (keyAdd_port_state_out_3_3_5 ), //o
    .port_state_out_3_3_6  (keyAdd_port_state_out_3_3_6 ), //o
    .port_state_out_3_3_7  (keyAdd_port_state_out_3_3_7 ), //o
    .port_state_out_4_0_0  (keyAdd_port_state_out_4_0_0 ), //o
    .port_state_out_4_0_1  (keyAdd_port_state_out_4_0_1 ), //o
    .port_state_out_4_0_2  (keyAdd_port_state_out_4_0_2 ), //o
    .port_state_out_4_0_3  (keyAdd_port_state_out_4_0_3 ), //o
    .port_state_out_4_0_4  (keyAdd_port_state_out_4_0_4 ), //o
    .port_state_out_4_0_5  (keyAdd_port_state_out_4_0_5 ), //o
    .port_state_out_4_0_6  (keyAdd_port_state_out_4_0_6 ), //o
    .port_state_out_4_0_7  (keyAdd_port_state_out_4_0_7 ), //o
    .port_state_out_4_1_0  (keyAdd_port_state_out_4_1_0 ), //o
    .port_state_out_4_1_1  (keyAdd_port_state_out_4_1_1 ), //o
    .port_state_out_4_1_2  (keyAdd_port_state_out_4_1_2 ), //o
    .port_state_out_4_1_3  (keyAdd_port_state_out_4_1_3 ), //o
    .port_state_out_4_1_4  (keyAdd_port_state_out_4_1_4 ), //o
    .port_state_out_4_1_5  (keyAdd_port_state_out_4_1_5 ), //o
    .port_state_out_4_1_6  (keyAdd_port_state_out_4_1_6 ), //o
    .port_state_out_4_1_7  (keyAdd_port_state_out_4_1_7 ), //o
    .port_state_out_4_2_0  (keyAdd_port_state_out_4_2_0 ), //o
    .port_state_out_4_2_1  (keyAdd_port_state_out_4_2_1 ), //o
    .port_state_out_4_2_2  (keyAdd_port_state_out_4_2_2 ), //o
    .port_state_out_4_2_3  (keyAdd_port_state_out_4_2_3 ), //o
    .port_state_out_4_2_4  (keyAdd_port_state_out_4_2_4 ), //o
    .port_state_out_4_2_5  (keyAdd_port_state_out_4_2_5 ), //o
    .port_state_out_4_2_6  (keyAdd_port_state_out_4_2_6 ), //o
    .port_state_out_4_2_7  (keyAdd_port_state_out_4_2_7 ), //o
    .port_state_out_4_3_0  (keyAdd_port_state_out_4_3_0 ), //o
    .port_state_out_4_3_1  (keyAdd_port_state_out_4_3_1 ), //o
    .port_state_out_4_3_2  (keyAdd_port_state_out_4_3_2 ), //o
    .port_state_out_4_3_3  (keyAdd_port_state_out_4_3_3 ), //o
    .port_state_out_4_3_4  (keyAdd_port_state_out_4_3_4 ), //o
    .port_state_out_4_3_5  (keyAdd_port_state_out_4_3_5 ), //o
    .port_state_out_4_3_6  (keyAdd_port_state_out_4_3_6 ), //o
    .port_state_out_4_3_7  (keyAdd_port_state_out_4_3_7 ), //o
    .port_state_out_5_0_0  (keyAdd_port_state_out_5_0_0 ), //o
    .port_state_out_5_0_1  (keyAdd_port_state_out_5_0_1 ), //o
    .port_state_out_5_0_2  (keyAdd_port_state_out_5_0_2 ), //o
    .port_state_out_5_0_3  (keyAdd_port_state_out_5_0_3 ), //o
    .port_state_out_5_0_4  (keyAdd_port_state_out_5_0_4 ), //o
    .port_state_out_5_0_5  (keyAdd_port_state_out_5_0_5 ), //o
    .port_state_out_5_0_6  (keyAdd_port_state_out_5_0_6 ), //o
    .port_state_out_5_0_7  (keyAdd_port_state_out_5_0_7 ), //o
    .port_state_out_5_1_0  (keyAdd_port_state_out_5_1_0 ), //o
    .port_state_out_5_1_1  (keyAdd_port_state_out_5_1_1 ), //o
    .port_state_out_5_1_2  (keyAdd_port_state_out_5_1_2 ), //o
    .port_state_out_5_1_3  (keyAdd_port_state_out_5_1_3 ), //o
    .port_state_out_5_1_4  (keyAdd_port_state_out_5_1_4 ), //o
    .port_state_out_5_1_5  (keyAdd_port_state_out_5_1_5 ), //o
    .port_state_out_5_1_6  (keyAdd_port_state_out_5_1_6 ), //o
    .port_state_out_5_1_7  (keyAdd_port_state_out_5_1_7 ), //o
    .port_state_out_5_2_0  (keyAdd_port_state_out_5_2_0 ), //o
    .port_state_out_5_2_1  (keyAdd_port_state_out_5_2_1 ), //o
    .port_state_out_5_2_2  (keyAdd_port_state_out_5_2_2 ), //o
    .port_state_out_5_2_3  (keyAdd_port_state_out_5_2_3 ), //o
    .port_state_out_5_2_4  (keyAdd_port_state_out_5_2_4 ), //o
    .port_state_out_5_2_5  (keyAdd_port_state_out_5_2_5 ), //o
    .port_state_out_5_2_6  (keyAdd_port_state_out_5_2_6 ), //o
    .port_state_out_5_2_7  (keyAdd_port_state_out_5_2_7 ), //o
    .port_state_out_5_3_0  (keyAdd_port_state_out_5_3_0 ), //o
    .port_state_out_5_3_1  (keyAdd_port_state_out_5_3_1 ), //o
    .port_state_out_5_3_2  (keyAdd_port_state_out_5_3_2 ), //o
    .port_state_out_5_3_3  (keyAdd_port_state_out_5_3_3 ), //o
    .port_state_out_5_3_4  (keyAdd_port_state_out_5_3_4 ), //o
    .port_state_out_5_3_5  (keyAdd_port_state_out_5_3_5 ), //o
    .port_state_out_5_3_6  (keyAdd_port_state_out_5_3_6 ), //o
    .port_state_out_5_3_7  (keyAdd_port_state_out_5_3_7 ), //o
    .port_state_out_6_0_0  (keyAdd_port_state_out_6_0_0 ), //o
    .port_state_out_6_0_1  (keyAdd_port_state_out_6_0_1 ), //o
    .port_state_out_6_0_2  (keyAdd_port_state_out_6_0_2 ), //o
    .port_state_out_6_0_3  (keyAdd_port_state_out_6_0_3 ), //o
    .port_state_out_6_0_4  (keyAdd_port_state_out_6_0_4 ), //o
    .port_state_out_6_0_5  (keyAdd_port_state_out_6_0_5 ), //o
    .port_state_out_6_0_6  (keyAdd_port_state_out_6_0_6 ), //o
    .port_state_out_6_0_7  (keyAdd_port_state_out_6_0_7 ), //o
    .port_state_out_6_1_0  (keyAdd_port_state_out_6_1_0 ), //o
    .port_state_out_6_1_1  (keyAdd_port_state_out_6_1_1 ), //o
    .port_state_out_6_1_2  (keyAdd_port_state_out_6_1_2 ), //o
    .port_state_out_6_1_3  (keyAdd_port_state_out_6_1_3 ), //o
    .port_state_out_6_1_4  (keyAdd_port_state_out_6_1_4 ), //o
    .port_state_out_6_1_5  (keyAdd_port_state_out_6_1_5 ), //o
    .port_state_out_6_1_6  (keyAdd_port_state_out_6_1_6 ), //o
    .port_state_out_6_1_7  (keyAdd_port_state_out_6_1_7 ), //o
    .port_state_out_6_2_0  (keyAdd_port_state_out_6_2_0 ), //o
    .port_state_out_6_2_1  (keyAdd_port_state_out_6_2_1 ), //o
    .port_state_out_6_2_2  (keyAdd_port_state_out_6_2_2 ), //o
    .port_state_out_6_2_3  (keyAdd_port_state_out_6_2_3 ), //o
    .port_state_out_6_2_4  (keyAdd_port_state_out_6_2_4 ), //o
    .port_state_out_6_2_5  (keyAdd_port_state_out_6_2_5 ), //o
    .port_state_out_6_2_6  (keyAdd_port_state_out_6_2_6 ), //o
    .port_state_out_6_2_7  (keyAdd_port_state_out_6_2_7 ), //o
    .port_state_out_6_3_0  (keyAdd_port_state_out_6_3_0 ), //o
    .port_state_out_6_3_1  (keyAdd_port_state_out_6_3_1 ), //o
    .port_state_out_6_3_2  (keyAdd_port_state_out_6_3_2 ), //o
    .port_state_out_6_3_3  (keyAdd_port_state_out_6_3_3 ), //o
    .port_state_out_6_3_4  (keyAdd_port_state_out_6_3_4 ), //o
    .port_state_out_6_3_5  (keyAdd_port_state_out_6_3_5 ), //o
    .port_state_out_6_3_6  (keyAdd_port_state_out_6_3_6 ), //o
    .port_state_out_6_3_7  (keyAdd_port_state_out_6_3_7 ), //o
    .port_state_out_7_0_0  (keyAdd_port_state_out_7_0_0 ), //o
    .port_state_out_7_0_1  (keyAdd_port_state_out_7_0_1 ), //o
    .port_state_out_7_0_2  (keyAdd_port_state_out_7_0_2 ), //o
    .port_state_out_7_0_3  (keyAdd_port_state_out_7_0_3 ), //o
    .port_state_out_7_0_4  (keyAdd_port_state_out_7_0_4 ), //o
    .port_state_out_7_0_5  (keyAdd_port_state_out_7_0_5 ), //o
    .port_state_out_7_0_6  (keyAdd_port_state_out_7_0_6 ), //o
    .port_state_out_7_0_7  (keyAdd_port_state_out_7_0_7 ), //o
    .port_state_out_7_1_0  (keyAdd_port_state_out_7_1_0 ), //o
    .port_state_out_7_1_1  (keyAdd_port_state_out_7_1_1 ), //o
    .port_state_out_7_1_2  (keyAdd_port_state_out_7_1_2 ), //o
    .port_state_out_7_1_3  (keyAdd_port_state_out_7_1_3 ), //o
    .port_state_out_7_1_4  (keyAdd_port_state_out_7_1_4 ), //o
    .port_state_out_7_1_5  (keyAdd_port_state_out_7_1_5 ), //o
    .port_state_out_7_1_6  (keyAdd_port_state_out_7_1_6 ), //o
    .port_state_out_7_1_7  (keyAdd_port_state_out_7_1_7 ), //o
    .port_state_out_7_2_0  (keyAdd_port_state_out_7_2_0 ), //o
    .port_state_out_7_2_1  (keyAdd_port_state_out_7_2_1 ), //o
    .port_state_out_7_2_2  (keyAdd_port_state_out_7_2_2 ), //o
    .port_state_out_7_2_3  (keyAdd_port_state_out_7_2_3 ), //o
    .port_state_out_7_2_4  (keyAdd_port_state_out_7_2_4 ), //o
    .port_state_out_7_2_5  (keyAdd_port_state_out_7_2_5 ), //o
    .port_state_out_7_2_6  (keyAdd_port_state_out_7_2_6 ), //o
    .port_state_out_7_2_7  (keyAdd_port_state_out_7_2_7 ), //o
    .port_state_out_7_3_0  (keyAdd_port_state_out_7_3_0 ), //o
    .port_state_out_7_3_1  (keyAdd_port_state_out_7_3_1 ), //o
    .port_state_out_7_3_2  (keyAdd_port_state_out_7_3_2 ), //o
    .port_state_out_7_3_3  (keyAdd_port_state_out_7_3_3 ), //o
    .port_state_out_7_3_4  (keyAdd_port_state_out_7_3_4 ), //o
    .port_state_out_7_3_5  (keyAdd_port_state_out_7_3_5 ), //o
    .port_state_out_7_3_6  (keyAdd_port_state_out_7_3_6 ), //o
    .port_state_out_7_3_7  (keyAdd_port_state_out_7_3_7 ), //o
    .port_state_out_8_0_0  (keyAdd_port_state_out_8_0_0 ), //o
    .port_state_out_8_0_1  (keyAdd_port_state_out_8_0_1 ), //o
    .port_state_out_8_0_2  (keyAdd_port_state_out_8_0_2 ), //o
    .port_state_out_8_0_3  (keyAdd_port_state_out_8_0_3 ), //o
    .port_state_out_8_0_4  (keyAdd_port_state_out_8_0_4 ), //o
    .port_state_out_8_0_5  (keyAdd_port_state_out_8_0_5 ), //o
    .port_state_out_8_0_6  (keyAdd_port_state_out_8_0_6 ), //o
    .port_state_out_8_0_7  (keyAdd_port_state_out_8_0_7 ), //o
    .port_state_out_8_1_0  (keyAdd_port_state_out_8_1_0 ), //o
    .port_state_out_8_1_1  (keyAdd_port_state_out_8_1_1 ), //o
    .port_state_out_8_1_2  (keyAdd_port_state_out_8_1_2 ), //o
    .port_state_out_8_1_3  (keyAdd_port_state_out_8_1_3 ), //o
    .port_state_out_8_1_4  (keyAdd_port_state_out_8_1_4 ), //o
    .port_state_out_8_1_5  (keyAdd_port_state_out_8_1_5 ), //o
    .port_state_out_8_1_6  (keyAdd_port_state_out_8_1_6 ), //o
    .port_state_out_8_1_7  (keyAdd_port_state_out_8_1_7 ), //o
    .port_state_out_8_2_0  (keyAdd_port_state_out_8_2_0 ), //o
    .port_state_out_8_2_1  (keyAdd_port_state_out_8_2_1 ), //o
    .port_state_out_8_2_2  (keyAdd_port_state_out_8_2_2 ), //o
    .port_state_out_8_2_3  (keyAdd_port_state_out_8_2_3 ), //o
    .port_state_out_8_2_4  (keyAdd_port_state_out_8_2_4 ), //o
    .port_state_out_8_2_5  (keyAdd_port_state_out_8_2_5 ), //o
    .port_state_out_8_2_6  (keyAdd_port_state_out_8_2_6 ), //o
    .port_state_out_8_2_7  (keyAdd_port_state_out_8_2_7 ), //o
    .port_state_out_8_3_0  (keyAdd_port_state_out_8_3_0 ), //o
    .port_state_out_8_3_1  (keyAdd_port_state_out_8_3_1 ), //o
    .port_state_out_8_3_2  (keyAdd_port_state_out_8_3_2 ), //o
    .port_state_out_8_3_3  (keyAdd_port_state_out_8_3_3 ), //o
    .port_state_out_8_3_4  (keyAdd_port_state_out_8_3_4 ), //o
    .port_state_out_8_3_5  (keyAdd_port_state_out_8_3_5 ), //o
    .port_state_out_8_3_6  (keyAdd_port_state_out_8_3_6 ), //o
    .port_state_out_8_3_7  (keyAdd_port_state_out_8_3_7 ), //o
    .port_state_out_9_0_0  (keyAdd_port_state_out_9_0_0 ), //o
    .port_state_out_9_0_1  (keyAdd_port_state_out_9_0_1 ), //o
    .port_state_out_9_0_2  (keyAdd_port_state_out_9_0_2 ), //o
    .port_state_out_9_0_3  (keyAdd_port_state_out_9_0_3 ), //o
    .port_state_out_9_0_4  (keyAdd_port_state_out_9_0_4 ), //o
    .port_state_out_9_0_5  (keyAdd_port_state_out_9_0_5 ), //o
    .port_state_out_9_0_6  (keyAdd_port_state_out_9_0_6 ), //o
    .port_state_out_9_0_7  (keyAdd_port_state_out_9_0_7 ), //o
    .port_state_out_9_1_0  (keyAdd_port_state_out_9_1_0 ), //o
    .port_state_out_9_1_1  (keyAdd_port_state_out_9_1_1 ), //o
    .port_state_out_9_1_2  (keyAdd_port_state_out_9_1_2 ), //o
    .port_state_out_9_1_3  (keyAdd_port_state_out_9_1_3 ), //o
    .port_state_out_9_1_4  (keyAdd_port_state_out_9_1_4 ), //o
    .port_state_out_9_1_5  (keyAdd_port_state_out_9_1_5 ), //o
    .port_state_out_9_1_6  (keyAdd_port_state_out_9_1_6 ), //o
    .port_state_out_9_1_7  (keyAdd_port_state_out_9_1_7 ), //o
    .port_state_out_9_2_0  (keyAdd_port_state_out_9_2_0 ), //o
    .port_state_out_9_2_1  (keyAdd_port_state_out_9_2_1 ), //o
    .port_state_out_9_2_2  (keyAdd_port_state_out_9_2_2 ), //o
    .port_state_out_9_2_3  (keyAdd_port_state_out_9_2_3 ), //o
    .port_state_out_9_2_4  (keyAdd_port_state_out_9_2_4 ), //o
    .port_state_out_9_2_5  (keyAdd_port_state_out_9_2_5 ), //o
    .port_state_out_9_2_6  (keyAdd_port_state_out_9_2_6 ), //o
    .port_state_out_9_2_7  (keyAdd_port_state_out_9_2_7 ), //o
    .port_state_out_9_3_0  (keyAdd_port_state_out_9_3_0 ), //o
    .port_state_out_9_3_1  (keyAdd_port_state_out_9_3_1 ), //o
    .port_state_out_9_3_2  (keyAdd_port_state_out_9_3_2 ), //o
    .port_state_out_9_3_3  (keyAdd_port_state_out_9_3_3 ), //o
    .port_state_out_9_3_4  (keyAdd_port_state_out_9_3_4 ), //o
    .port_state_out_9_3_5  (keyAdd_port_state_out_9_3_5 ), //o
    .port_state_out_9_3_6  (keyAdd_port_state_out_9_3_6 ), //o
    .port_state_out_9_3_7  (keyAdd_port_state_out_9_3_7 ), //o
    .port_state_out_10_0_0 (keyAdd_port_state_out_10_0_0), //o
    .port_state_out_10_0_1 (keyAdd_port_state_out_10_0_1), //o
    .port_state_out_10_0_2 (keyAdd_port_state_out_10_0_2), //o
    .port_state_out_10_0_3 (keyAdd_port_state_out_10_0_3), //o
    .port_state_out_10_0_4 (keyAdd_port_state_out_10_0_4), //o
    .port_state_out_10_0_5 (keyAdd_port_state_out_10_0_5), //o
    .port_state_out_10_0_6 (keyAdd_port_state_out_10_0_6), //o
    .port_state_out_10_0_7 (keyAdd_port_state_out_10_0_7), //o
    .port_state_out_10_1_0 (keyAdd_port_state_out_10_1_0), //o
    .port_state_out_10_1_1 (keyAdd_port_state_out_10_1_1), //o
    .port_state_out_10_1_2 (keyAdd_port_state_out_10_1_2), //o
    .port_state_out_10_1_3 (keyAdd_port_state_out_10_1_3), //o
    .port_state_out_10_1_4 (keyAdd_port_state_out_10_1_4), //o
    .port_state_out_10_1_5 (keyAdd_port_state_out_10_1_5), //o
    .port_state_out_10_1_6 (keyAdd_port_state_out_10_1_6), //o
    .port_state_out_10_1_7 (keyAdd_port_state_out_10_1_7), //o
    .port_state_out_10_2_0 (keyAdd_port_state_out_10_2_0), //o
    .port_state_out_10_2_1 (keyAdd_port_state_out_10_2_1), //o
    .port_state_out_10_2_2 (keyAdd_port_state_out_10_2_2), //o
    .port_state_out_10_2_3 (keyAdd_port_state_out_10_2_3), //o
    .port_state_out_10_2_4 (keyAdd_port_state_out_10_2_4), //o
    .port_state_out_10_2_5 (keyAdd_port_state_out_10_2_5), //o
    .port_state_out_10_2_6 (keyAdd_port_state_out_10_2_6), //o
    .port_state_out_10_2_7 (keyAdd_port_state_out_10_2_7), //o
    .port_state_out_10_3_0 (keyAdd_port_state_out_10_3_0), //o
    .port_state_out_10_3_1 (keyAdd_port_state_out_10_3_1), //o
    .port_state_out_10_3_2 (keyAdd_port_state_out_10_3_2), //o
    .port_state_out_10_3_3 (keyAdd_port_state_out_10_3_3), //o
    .port_state_out_10_3_4 (keyAdd_port_state_out_10_3_4), //o
    .port_state_out_10_3_5 (keyAdd_port_state_out_10_3_5), //o
    .port_state_out_10_3_6 (keyAdd_port_state_out_10_3_6), //o
    .port_state_out_10_3_7 (keyAdd_port_state_out_10_3_7), //o
    .port_state_out_11_0_0 (keyAdd_port_state_out_11_0_0), //o
    .port_state_out_11_0_1 (keyAdd_port_state_out_11_0_1), //o
    .port_state_out_11_0_2 (keyAdd_port_state_out_11_0_2), //o
    .port_state_out_11_0_3 (keyAdd_port_state_out_11_0_3), //o
    .port_state_out_11_0_4 (keyAdd_port_state_out_11_0_4), //o
    .port_state_out_11_0_5 (keyAdd_port_state_out_11_0_5), //o
    .port_state_out_11_0_6 (keyAdd_port_state_out_11_0_6), //o
    .port_state_out_11_0_7 (keyAdd_port_state_out_11_0_7), //o
    .port_state_out_11_1_0 (keyAdd_port_state_out_11_1_0), //o
    .port_state_out_11_1_1 (keyAdd_port_state_out_11_1_1), //o
    .port_state_out_11_1_2 (keyAdd_port_state_out_11_1_2), //o
    .port_state_out_11_1_3 (keyAdd_port_state_out_11_1_3), //o
    .port_state_out_11_1_4 (keyAdd_port_state_out_11_1_4), //o
    .port_state_out_11_1_5 (keyAdd_port_state_out_11_1_5), //o
    .port_state_out_11_1_6 (keyAdd_port_state_out_11_1_6), //o
    .port_state_out_11_1_7 (keyAdd_port_state_out_11_1_7), //o
    .port_state_out_11_2_0 (keyAdd_port_state_out_11_2_0), //o
    .port_state_out_11_2_1 (keyAdd_port_state_out_11_2_1), //o
    .port_state_out_11_2_2 (keyAdd_port_state_out_11_2_2), //o
    .port_state_out_11_2_3 (keyAdd_port_state_out_11_2_3), //o
    .port_state_out_11_2_4 (keyAdd_port_state_out_11_2_4), //o
    .port_state_out_11_2_5 (keyAdd_port_state_out_11_2_5), //o
    .port_state_out_11_2_6 (keyAdd_port_state_out_11_2_6), //o
    .port_state_out_11_2_7 (keyAdd_port_state_out_11_2_7), //o
    .port_state_out_11_3_0 (keyAdd_port_state_out_11_3_0), //o
    .port_state_out_11_3_1 (keyAdd_port_state_out_11_3_1), //o
    .port_state_out_11_3_2 (keyAdd_port_state_out_11_3_2), //o
    .port_state_out_11_3_3 (keyAdd_port_state_out_11_3_3), //o
    .port_state_out_11_3_4 (keyAdd_port_state_out_11_3_4), //o
    .port_state_out_11_3_5 (keyAdd_port_state_out_11_3_5), //o
    .port_state_out_11_3_6 (keyAdd_port_state_out_11_3_6), //o
    .port_state_out_11_3_7 (keyAdd_port_state_out_11_3_7), //o
    .port_state_out_12_0_0 (keyAdd_port_state_out_12_0_0), //o
    .port_state_out_12_0_1 (keyAdd_port_state_out_12_0_1), //o
    .port_state_out_12_0_2 (keyAdd_port_state_out_12_0_2), //o
    .port_state_out_12_0_3 (keyAdd_port_state_out_12_0_3), //o
    .port_state_out_12_0_4 (keyAdd_port_state_out_12_0_4), //o
    .port_state_out_12_0_5 (keyAdd_port_state_out_12_0_5), //o
    .port_state_out_12_0_6 (keyAdd_port_state_out_12_0_6), //o
    .port_state_out_12_0_7 (keyAdd_port_state_out_12_0_7), //o
    .port_state_out_12_1_0 (keyAdd_port_state_out_12_1_0), //o
    .port_state_out_12_1_1 (keyAdd_port_state_out_12_1_1), //o
    .port_state_out_12_1_2 (keyAdd_port_state_out_12_1_2), //o
    .port_state_out_12_1_3 (keyAdd_port_state_out_12_1_3), //o
    .port_state_out_12_1_4 (keyAdd_port_state_out_12_1_4), //o
    .port_state_out_12_1_5 (keyAdd_port_state_out_12_1_5), //o
    .port_state_out_12_1_6 (keyAdd_port_state_out_12_1_6), //o
    .port_state_out_12_1_7 (keyAdd_port_state_out_12_1_7), //o
    .port_state_out_12_2_0 (keyAdd_port_state_out_12_2_0), //o
    .port_state_out_12_2_1 (keyAdd_port_state_out_12_2_1), //o
    .port_state_out_12_2_2 (keyAdd_port_state_out_12_2_2), //o
    .port_state_out_12_2_3 (keyAdd_port_state_out_12_2_3), //o
    .port_state_out_12_2_4 (keyAdd_port_state_out_12_2_4), //o
    .port_state_out_12_2_5 (keyAdd_port_state_out_12_2_5), //o
    .port_state_out_12_2_6 (keyAdd_port_state_out_12_2_6), //o
    .port_state_out_12_2_7 (keyAdd_port_state_out_12_2_7), //o
    .port_state_out_12_3_0 (keyAdd_port_state_out_12_3_0), //o
    .port_state_out_12_3_1 (keyAdd_port_state_out_12_3_1), //o
    .port_state_out_12_3_2 (keyAdd_port_state_out_12_3_2), //o
    .port_state_out_12_3_3 (keyAdd_port_state_out_12_3_3), //o
    .port_state_out_12_3_4 (keyAdd_port_state_out_12_3_4), //o
    .port_state_out_12_3_5 (keyAdd_port_state_out_12_3_5), //o
    .port_state_out_12_3_6 (keyAdd_port_state_out_12_3_6), //o
    .port_state_out_12_3_7 (keyAdd_port_state_out_12_3_7), //o
    .port_state_out_13_0_0 (keyAdd_port_state_out_13_0_0), //o
    .port_state_out_13_0_1 (keyAdd_port_state_out_13_0_1), //o
    .port_state_out_13_0_2 (keyAdd_port_state_out_13_0_2), //o
    .port_state_out_13_0_3 (keyAdd_port_state_out_13_0_3), //o
    .port_state_out_13_0_4 (keyAdd_port_state_out_13_0_4), //o
    .port_state_out_13_0_5 (keyAdd_port_state_out_13_0_5), //o
    .port_state_out_13_0_6 (keyAdd_port_state_out_13_0_6), //o
    .port_state_out_13_0_7 (keyAdd_port_state_out_13_0_7), //o
    .port_state_out_13_1_0 (keyAdd_port_state_out_13_1_0), //o
    .port_state_out_13_1_1 (keyAdd_port_state_out_13_1_1), //o
    .port_state_out_13_1_2 (keyAdd_port_state_out_13_1_2), //o
    .port_state_out_13_1_3 (keyAdd_port_state_out_13_1_3), //o
    .port_state_out_13_1_4 (keyAdd_port_state_out_13_1_4), //o
    .port_state_out_13_1_5 (keyAdd_port_state_out_13_1_5), //o
    .port_state_out_13_1_6 (keyAdd_port_state_out_13_1_6), //o
    .port_state_out_13_1_7 (keyAdd_port_state_out_13_1_7), //o
    .port_state_out_13_2_0 (keyAdd_port_state_out_13_2_0), //o
    .port_state_out_13_2_1 (keyAdd_port_state_out_13_2_1), //o
    .port_state_out_13_2_2 (keyAdd_port_state_out_13_2_2), //o
    .port_state_out_13_2_3 (keyAdd_port_state_out_13_2_3), //o
    .port_state_out_13_2_4 (keyAdd_port_state_out_13_2_4), //o
    .port_state_out_13_2_5 (keyAdd_port_state_out_13_2_5), //o
    .port_state_out_13_2_6 (keyAdd_port_state_out_13_2_6), //o
    .port_state_out_13_2_7 (keyAdd_port_state_out_13_2_7), //o
    .port_state_out_13_3_0 (keyAdd_port_state_out_13_3_0), //o
    .port_state_out_13_3_1 (keyAdd_port_state_out_13_3_1), //o
    .port_state_out_13_3_2 (keyAdd_port_state_out_13_3_2), //o
    .port_state_out_13_3_3 (keyAdd_port_state_out_13_3_3), //o
    .port_state_out_13_3_4 (keyAdd_port_state_out_13_3_4), //o
    .port_state_out_13_3_5 (keyAdd_port_state_out_13_3_5), //o
    .port_state_out_13_3_6 (keyAdd_port_state_out_13_3_6), //o
    .port_state_out_13_3_7 (keyAdd_port_state_out_13_3_7), //o
    .port_state_out_14_0_0 (keyAdd_port_state_out_14_0_0), //o
    .port_state_out_14_0_1 (keyAdd_port_state_out_14_0_1), //o
    .port_state_out_14_0_2 (keyAdd_port_state_out_14_0_2), //o
    .port_state_out_14_0_3 (keyAdd_port_state_out_14_0_3), //o
    .port_state_out_14_0_4 (keyAdd_port_state_out_14_0_4), //o
    .port_state_out_14_0_5 (keyAdd_port_state_out_14_0_5), //o
    .port_state_out_14_0_6 (keyAdd_port_state_out_14_0_6), //o
    .port_state_out_14_0_7 (keyAdd_port_state_out_14_0_7), //o
    .port_state_out_14_1_0 (keyAdd_port_state_out_14_1_0), //o
    .port_state_out_14_1_1 (keyAdd_port_state_out_14_1_1), //o
    .port_state_out_14_1_2 (keyAdd_port_state_out_14_1_2), //o
    .port_state_out_14_1_3 (keyAdd_port_state_out_14_1_3), //o
    .port_state_out_14_1_4 (keyAdd_port_state_out_14_1_4), //o
    .port_state_out_14_1_5 (keyAdd_port_state_out_14_1_5), //o
    .port_state_out_14_1_6 (keyAdd_port_state_out_14_1_6), //o
    .port_state_out_14_1_7 (keyAdd_port_state_out_14_1_7), //o
    .port_state_out_14_2_0 (keyAdd_port_state_out_14_2_0), //o
    .port_state_out_14_2_1 (keyAdd_port_state_out_14_2_1), //o
    .port_state_out_14_2_2 (keyAdd_port_state_out_14_2_2), //o
    .port_state_out_14_2_3 (keyAdd_port_state_out_14_2_3), //o
    .port_state_out_14_2_4 (keyAdd_port_state_out_14_2_4), //o
    .port_state_out_14_2_5 (keyAdd_port_state_out_14_2_5), //o
    .port_state_out_14_2_6 (keyAdd_port_state_out_14_2_6), //o
    .port_state_out_14_2_7 (keyAdd_port_state_out_14_2_7), //o
    .port_state_out_14_3_0 (keyAdd_port_state_out_14_3_0), //o
    .port_state_out_14_3_1 (keyAdd_port_state_out_14_3_1), //o
    .port_state_out_14_3_2 (keyAdd_port_state_out_14_3_2), //o
    .port_state_out_14_3_3 (keyAdd_port_state_out_14_3_3), //o
    .port_state_out_14_3_4 (keyAdd_port_state_out_14_3_4), //o
    .port_state_out_14_3_5 (keyAdd_port_state_out_14_3_5), //o
    .port_state_out_14_3_6 (keyAdd_port_state_out_14_3_6), //o
    .port_state_out_14_3_7 (keyAdd_port_state_out_14_3_7), //o
    .port_state_out_15_0_0 (keyAdd_port_state_out_15_0_0), //o
    .port_state_out_15_0_1 (keyAdd_port_state_out_15_0_1), //o
    .port_state_out_15_0_2 (keyAdd_port_state_out_15_0_2), //o
    .port_state_out_15_0_3 (keyAdd_port_state_out_15_0_3), //o
    .port_state_out_15_0_4 (keyAdd_port_state_out_15_0_4), //o
    .port_state_out_15_0_5 (keyAdd_port_state_out_15_0_5), //o
    .port_state_out_15_0_6 (keyAdd_port_state_out_15_0_6), //o
    .port_state_out_15_0_7 (keyAdd_port_state_out_15_0_7), //o
    .port_state_out_15_1_0 (keyAdd_port_state_out_15_1_0), //o
    .port_state_out_15_1_1 (keyAdd_port_state_out_15_1_1), //o
    .port_state_out_15_1_2 (keyAdd_port_state_out_15_1_2), //o
    .port_state_out_15_1_3 (keyAdd_port_state_out_15_1_3), //o
    .port_state_out_15_1_4 (keyAdd_port_state_out_15_1_4), //o
    .port_state_out_15_1_5 (keyAdd_port_state_out_15_1_5), //o
    .port_state_out_15_1_6 (keyAdd_port_state_out_15_1_6), //o
    .port_state_out_15_1_7 (keyAdd_port_state_out_15_1_7), //o
    .port_state_out_15_2_0 (keyAdd_port_state_out_15_2_0), //o
    .port_state_out_15_2_1 (keyAdd_port_state_out_15_2_1), //o
    .port_state_out_15_2_2 (keyAdd_port_state_out_15_2_2), //o
    .port_state_out_15_2_3 (keyAdd_port_state_out_15_2_3), //o
    .port_state_out_15_2_4 (keyAdd_port_state_out_15_2_4), //o
    .port_state_out_15_2_5 (keyAdd_port_state_out_15_2_5), //o
    .port_state_out_15_2_6 (keyAdd_port_state_out_15_2_6), //o
    .port_state_out_15_2_7 (keyAdd_port_state_out_15_2_7), //o
    .port_state_out_15_3_0 (keyAdd_port_state_out_15_3_0), //o
    .port_state_out_15_3_1 (keyAdd_port_state_out_15_3_1), //o
    .port_state_out_15_3_2 (keyAdd_port_state_out_15_3_2), //o
    .port_state_out_15_3_3 (keyAdd_port_state_out_15_3_3), //o
    .port_state_out_15_3_4 (keyAdd_port_state_out_15_3_4), //o
    .port_state_out_15_3_5 (keyAdd_port_state_out_15_3_5), //o
    .port_state_out_15_3_6 (keyAdd_port_state_out_15_3_6), //o
    .port_state_out_15_3_7 (keyAdd_port_state_out_15_3_7)  //o
  );
  Sbox_AES_BoyarPeralta sbox_AES_BoyarPeralta_16 (
    .port_i_0_0 (keyAdd_port_state_out_0_0_0        ), //i
    .port_i_0_1 (keyAdd_port_state_out_0_0_1        ), //i
    .port_i_0_2 (keyAdd_port_state_out_0_0_2        ), //i
    .port_i_0_3 (keyAdd_port_state_out_0_0_3        ), //i
    .port_i_0_4 (keyAdd_port_state_out_0_0_4        ), //i
    .port_i_0_5 (keyAdd_port_state_out_0_0_5        ), //i
    .port_i_0_6 (keyAdd_port_state_out_0_0_6        ), //i
    .port_i_0_7 (keyAdd_port_state_out_0_0_7        ), //i
    .port_i_1_0 (keyAdd_port_state_out_0_1_0        ), //i
    .port_i_1_1 (keyAdd_port_state_out_0_1_1        ), //i
    .port_i_1_2 (keyAdd_port_state_out_0_1_2        ), //i
    .port_i_1_3 (keyAdd_port_state_out_0_1_3        ), //i
    .port_i_1_4 (keyAdd_port_state_out_0_1_4        ), //i
    .port_i_1_5 (keyAdd_port_state_out_0_1_5        ), //i
    .port_i_1_6 (keyAdd_port_state_out_0_1_6        ), //i
    .port_i_1_7 (keyAdd_port_state_out_0_1_7        ), //i
    .port_i_2_0 (keyAdd_port_state_out_0_2_0        ), //i
    .port_i_2_1 (keyAdd_port_state_out_0_2_1        ), //i
    .port_i_2_2 (keyAdd_port_state_out_0_2_2        ), //i
    .port_i_2_3 (keyAdd_port_state_out_0_2_3        ), //i
    .port_i_2_4 (keyAdd_port_state_out_0_2_4        ), //i
    .port_i_2_5 (keyAdd_port_state_out_0_2_5        ), //i
    .port_i_2_6 (keyAdd_port_state_out_0_2_6        ), //i
    .port_i_2_7 (keyAdd_port_state_out_0_2_7        ), //i
    .port_i_3_0 (keyAdd_port_state_out_0_3_0        ), //i
    .port_i_3_1 (keyAdd_port_state_out_0_3_1        ), //i
    .port_i_3_2 (keyAdd_port_state_out_0_3_2        ), //i
    .port_i_3_3 (keyAdd_port_state_out_0_3_3        ), //i
    .port_i_3_4 (keyAdd_port_state_out_0_3_4        ), //i
    .port_i_3_5 (keyAdd_port_state_out_0_3_5        ), //i
    .port_i_3_6 (keyAdd_port_state_out_0_3_6        ), //i
    .port_i_3_7 (keyAdd_port_state_out_0_3_7        ), //i
    .port_o_0_0 (sbox_AES_BoyarPeralta_16_port_o_0_0), //o
    .port_o_0_1 (sbox_AES_BoyarPeralta_16_port_o_0_1), //o
    .port_o_0_2 (sbox_AES_BoyarPeralta_16_port_o_0_2), //o
    .port_o_0_3 (sbox_AES_BoyarPeralta_16_port_o_0_3), //o
    .port_o_0_4 (sbox_AES_BoyarPeralta_16_port_o_0_4), //o
    .port_o_0_5 (sbox_AES_BoyarPeralta_16_port_o_0_5), //o
    .port_o_0_6 (sbox_AES_BoyarPeralta_16_port_o_0_6), //o
    .port_o_0_7 (sbox_AES_BoyarPeralta_16_port_o_0_7), //o
    .port_o_1_0 (sbox_AES_BoyarPeralta_16_port_o_1_0), //o
    .port_o_1_1 (sbox_AES_BoyarPeralta_16_port_o_1_1), //o
    .port_o_1_2 (sbox_AES_BoyarPeralta_16_port_o_1_2), //o
    .port_o_1_3 (sbox_AES_BoyarPeralta_16_port_o_1_3), //o
    .port_o_1_4 (sbox_AES_BoyarPeralta_16_port_o_1_4), //o
    .port_o_1_5 (sbox_AES_BoyarPeralta_16_port_o_1_5), //o
    .port_o_1_6 (sbox_AES_BoyarPeralta_16_port_o_1_6), //o
    .port_o_1_7 (sbox_AES_BoyarPeralta_16_port_o_1_7), //o
    .port_o_2_0 (sbox_AES_BoyarPeralta_16_port_o_2_0), //o
    .port_o_2_1 (sbox_AES_BoyarPeralta_16_port_o_2_1), //o
    .port_o_2_2 (sbox_AES_BoyarPeralta_16_port_o_2_2), //o
    .port_o_2_3 (sbox_AES_BoyarPeralta_16_port_o_2_3), //o
    .port_o_2_4 (sbox_AES_BoyarPeralta_16_port_o_2_4), //o
    .port_o_2_5 (sbox_AES_BoyarPeralta_16_port_o_2_5), //o
    .port_o_2_6 (sbox_AES_BoyarPeralta_16_port_o_2_6), //o
    .port_o_2_7 (sbox_AES_BoyarPeralta_16_port_o_2_7), //o
    .port_o_3_0 (sbox_AES_BoyarPeralta_16_port_o_3_0), //o
    .port_o_3_1 (sbox_AES_BoyarPeralta_16_port_o_3_1), //o
    .port_o_3_2 (sbox_AES_BoyarPeralta_16_port_o_3_2), //o
    .port_o_3_3 (sbox_AES_BoyarPeralta_16_port_o_3_3), //o
    .port_o_3_4 (sbox_AES_BoyarPeralta_16_port_o_3_4), //o
    .port_o_3_5 (sbox_AES_BoyarPeralta_16_port_o_3_5), //o
    .port_o_3_6 (sbox_AES_BoyarPeralta_16_port_o_3_6), //o
    .port_o_3_7 (sbox_AES_BoyarPeralta_16_port_o_3_7), //o
    .clk        (clk                                ), //i
    .reset      (reset                              )  //i
  );
  Sbox_AES_BoyarPeralta sbox_AES_BoyarPeralta_17 (
    .port_i_0_0 (keyAdd_port_state_out_1_0_0        ), //i
    .port_i_0_1 (keyAdd_port_state_out_1_0_1        ), //i
    .port_i_0_2 (keyAdd_port_state_out_1_0_2        ), //i
    .port_i_0_3 (keyAdd_port_state_out_1_0_3        ), //i
    .port_i_0_4 (keyAdd_port_state_out_1_0_4        ), //i
    .port_i_0_5 (keyAdd_port_state_out_1_0_5        ), //i
    .port_i_0_6 (keyAdd_port_state_out_1_0_6        ), //i
    .port_i_0_7 (keyAdd_port_state_out_1_0_7        ), //i
    .port_i_1_0 (keyAdd_port_state_out_1_1_0        ), //i
    .port_i_1_1 (keyAdd_port_state_out_1_1_1        ), //i
    .port_i_1_2 (keyAdd_port_state_out_1_1_2        ), //i
    .port_i_1_3 (keyAdd_port_state_out_1_1_3        ), //i
    .port_i_1_4 (keyAdd_port_state_out_1_1_4        ), //i
    .port_i_1_5 (keyAdd_port_state_out_1_1_5        ), //i
    .port_i_1_6 (keyAdd_port_state_out_1_1_6        ), //i
    .port_i_1_7 (keyAdd_port_state_out_1_1_7        ), //i
    .port_i_2_0 (keyAdd_port_state_out_1_2_0        ), //i
    .port_i_2_1 (keyAdd_port_state_out_1_2_1        ), //i
    .port_i_2_2 (keyAdd_port_state_out_1_2_2        ), //i
    .port_i_2_3 (keyAdd_port_state_out_1_2_3        ), //i
    .port_i_2_4 (keyAdd_port_state_out_1_2_4        ), //i
    .port_i_2_5 (keyAdd_port_state_out_1_2_5        ), //i
    .port_i_2_6 (keyAdd_port_state_out_1_2_6        ), //i
    .port_i_2_7 (keyAdd_port_state_out_1_2_7        ), //i
    .port_i_3_0 (keyAdd_port_state_out_1_3_0        ), //i
    .port_i_3_1 (keyAdd_port_state_out_1_3_1        ), //i
    .port_i_3_2 (keyAdd_port_state_out_1_3_2        ), //i
    .port_i_3_3 (keyAdd_port_state_out_1_3_3        ), //i
    .port_i_3_4 (keyAdd_port_state_out_1_3_4        ), //i
    .port_i_3_5 (keyAdd_port_state_out_1_3_5        ), //i
    .port_i_3_6 (keyAdd_port_state_out_1_3_6        ), //i
    .port_i_3_7 (keyAdd_port_state_out_1_3_7        ), //i
    .port_o_0_0 (sbox_AES_BoyarPeralta_17_port_o_0_0), //o
    .port_o_0_1 (sbox_AES_BoyarPeralta_17_port_o_0_1), //o
    .port_o_0_2 (sbox_AES_BoyarPeralta_17_port_o_0_2), //o
    .port_o_0_3 (sbox_AES_BoyarPeralta_17_port_o_0_3), //o
    .port_o_0_4 (sbox_AES_BoyarPeralta_17_port_o_0_4), //o
    .port_o_0_5 (sbox_AES_BoyarPeralta_17_port_o_0_5), //o
    .port_o_0_6 (sbox_AES_BoyarPeralta_17_port_o_0_6), //o
    .port_o_0_7 (sbox_AES_BoyarPeralta_17_port_o_0_7), //o
    .port_o_1_0 (sbox_AES_BoyarPeralta_17_port_o_1_0), //o
    .port_o_1_1 (sbox_AES_BoyarPeralta_17_port_o_1_1), //o
    .port_o_1_2 (sbox_AES_BoyarPeralta_17_port_o_1_2), //o
    .port_o_1_3 (sbox_AES_BoyarPeralta_17_port_o_1_3), //o
    .port_o_1_4 (sbox_AES_BoyarPeralta_17_port_o_1_4), //o
    .port_o_1_5 (sbox_AES_BoyarPeralta_17_port_o_1_5), //o
    .port_o_1_6 (sbox_AES_BoyarPeralta_17_port_o_1_6), //o
    .port_o_1_7 (sbox_AES_BoyarPeralta_17_port_o_1_7), //o
    .port_o_2_0 (sbox_AES_BoyarPeralta_17_port_o_2_0), //o
    .port_o_2_1 (sbox_AES_BoyarPeralta_17_port_o_2_1), //o
    .port_o_2_2 (sbox_AES_BoyarPeralta_17_port_o_2_2), //o
    .port_o_2_3 (sbox_AES_BoyarPeralta_17_port_o_2_3), //o
    .port_o_2_4 (sbox_AES_BoyarPeralta_17_port_o_2_4), //o
    .port_o_2_5 (sbox_AES_BoyarPeralta_17_port_o_2_5), //o
    .port_o_2_6 (sbox_AES_BoyarPeralta_17_port_o_2_6), //o
    .port_o_2_7 (sbox_AES_BoyarPeralta_17_port_o_2_7), //o
    .port_o_3_0 (sbox_AES_BoyarPeralta_17_port_o_3_0), //o
    .port_o_3_1 (sbox_AES_BoyarPeralta_17_port_o_3_1), //o
    .port_o_3_2 (sbox_AES_BoyarPeralta_17_port_o_3_2), //o
    .port_o_3_3 (sbox_AES_BoyarPeralta_17_port_o_3_3), //o
    .port_o_3_4 (sbox_AES_BoyarPeralta_17_port_o_3_4), //o
    .port_o_3_5 (sbox_AES_BoyarPeralta_17_port_o_3_5), //o
    .port_o_3_6 (sbox_AES_BoyarPeralta_17_port_o_3_6), //o
    .port_o_3_7 (sbox_AES_BoyarPeralta_17_port_o_3_7), //o
    .clk        (clk                                ), //i
    .reset      (reset                              )  //i
  );
  Sbox_AES_BoyarPeralta sbox_AES_BoyarPeralta_18 (
    .port_i_0_0 (keyAdd_port_state_out_2_0_0        ), //i
    .port_i_0_1 (keyAdd_port_state_out_2_0_1        ), //i
    .port_i_0_2 (keyAdd_port_state_out_2_0_2        ), //i
    .port_i_0_3 (keyAdd_port_state_out_2_0_3        ), //i
    .port_i_0_4 (keyAdd_port_state_out_2_0_4        ), //i
    .port_i_0_5 (keyAdd_port_state_out_2_0_5        ), //i
    .port_i_0_6 (keyAdd_port_state_out_2_0_6        ), //i
    .port_i_0_7 (keyAdd_port_state_out_2_0_7        ), //i
    .port_i_1_0 (keyAdd_port_state_out_2_1_0        ), //i
    .port_i_1_1 (keyAdd_port_state_out_2_1_1        ), //i
    .port_i_1_2 (keyAdd_port_state_out_2_1_2        ), //i
    .port_i_1_3 (keyAdd_port_state_out_2_1_3        ), //i
    .port_i_1_4 (keyAdd_port_state_out_2_1_4        ), //i
    .port_i_1_5 (keyAdd_port_state_out_2_1_5        ), //i
    .port_i_1_6 (keyAdd_port_state_out_2_1_6        ), //i
    .port_i_1_7 (keyAdd_port_state_out_2_1_7        ), //i
    .port_i_2_0 (keyAdd_port_state_out_2_2_0        ), //i
    .port_i_2_1 (keyAdd_port_state_out_2_2_1        ), //i
    .port_i_2_2 (keyAdd_port_state_out_2_2_2        ), //i
    .port_i_2_3 (keyAdd_port_state_out_2_2_3        ), //i
    .port_i_2_4 (keyAdd_port_state_out_2_2_4        ), //i
    .port_i_2_5 (keyAdd_port_state_out_2_2_5        ), //i
    .port_i_2_6 (keyAdd_port_state_out_2_2_6        ), //i
    .port_i_2_7 (keyAdd_port_state_out_2_2_7        ), //i
    .port_i_3_0 (keyAdd_port_state_out_2_3_0        ), //i
    .port_i_3_1 (keyAdd_port_state_out_2_3_1        ), //i
    .port_i_3_2 (keyAdd_port_state_out_2_3_2        ), //i
    .port_i_3_3 (keyAdd_port_state_out_2_3_3        ), //i
    .port_i_3_4 (keyAdd_port_state_out_2_3_4        ), //i
    .port_i_3_5 (keyAdd_port_state_out_2_3_5        ), //i
    .port_i_3_6 (keyAdd_port_state_out_2_3_6        ), //i
    .port_i_3_7 (keyAdd_port_state_out_2_3_7        ), //i
    .port_o_0_0 (sbox_AES_BoyarPeralta_18_port_o_0_0), //o
    .port_o_0_1 (sbox_AES_BoyarPeralta_18_port_o_0_1), //o
    .port_o_0_2 (sbox_AES_BoyarPeralta_18_port_o_0_2), //o
    .port_o_0_3 (sbox_AES_BoyarPeralta_18_port_o_0_3), //o
    .port_o_0_4 (sbox_AES_BoyarPeralta_18_port_o_0_4), //o
    .port_o_0_5 (sbox_AES_BoyarPeralta_18_port_o_0_5), //o
    .port_o_0_6 (sbox_AES_BoyarPeralta_18_port_o_0_6), //o
    .port_o_0_7 (sbox_AES_BoyarPeralta_18_port_o_0_7), //o
    .port_o_1_0 (sbox_AES_BoyarPeralta_18_port_o_1_0), //o
    .port_o_1_1 (sbox_AES_BoyarPeralta_18_port_o_1_1), //o
    .port_o_1_2 (sbox_AES_BoyarPeralta_18_port_o_1_2), //o
    .port_o_1_3 (sbox_AES_BoyarPeralta_18_port_o_1_3), //o
    .port_o_1_4 (sbox_AES_BoyarPeralta_18_port_o_1_4), //o
    .port_o_1_5 (sbox_AES_BoyarPeralta_18_port_o_1_5), //o
    .port_o_1_6 (sbox_AES_BoyarPeralta_18_port_o_1_6), //o
    .port_o_1_7 (sbox_AES_BoyarPeralta_18_port_o_1_7), //o
    .port_o_2_0 (sbox_AES_BoyarPeralta_18_port_o_2_0), //o
    .port_o_2_1 (sbox_AES_BoyarPeralta_18_port_o_2_1), //o
    .port_o_2_2 (sbox_AES_BoyarPeralta_18_port_o_2_2), //o
    .port_o_2_3 (sbox_AES_BoyarPeralta_18_port_o_2_3), //o
    .port_o_2_4 (sbox_AES_BoyarPeralta_18_port_o_2_4), //o
    .port_o_2_5 (sbox_AES_BoyarPeralta_18_port_o_2_5), //o
    .port_o_2_6 (sbox_AES_BoyarPeralta_18_port_o_2_6), //o
    .port_o_2_7 (sbox_AES_BoyarPeralta_18_port_o_2_7), //o
    .port_o_3_0 (sbox_AES_BoyarPeralta_18_port_o_3_0), //o
    .port_o_3_1 (sbox_AES_BoyarPeralta_18_port_o_3_1), //o
    .port_o_3_2 (sbox_AES_BoyarPeralta_18_port_o_3_2), //o
    .port_o_3_3 (sbox_AES_BoyarPeralta_18_port_o_3_3), //o
    .port_o_3_4 (sbox_AES_BoyarPeralta_18_port_o_3_4), //o
    .port_o_3_5 (sbox_AES_BoyarPeralta_18_port_o_3_5), //o
    .port_o_3_6 (sbox_AES_BoyarPeralta_18_port_o_3_6), //o
    .port_o_3_7 (sbox_AES_BoyarPeralta_18_port_o_3_7), //o
    .clk        (clk                                ), //i
    .reset      (reset                              )  //i
  );
  Sbox_AES_BoyarPeralta sbox_AES_BoyarPeralta_19 (
    .port_i_0_0 (keyAdd_port_state_out_3_0_0        ), //i
    .port_i_0_1 (keyAdd_port_state_out_3_0_1        ), //i
    .port_i_0_2 (keyAdd_port_state_out_3_0_2        ), //i
    .port_i_0_3 (keyAdd_port_state_out_3_0_3        ), //i
    .port_i_0_4 (keyAdd_port_state_out_3_0_4        ), //i
    .port_i_0_5 (keyAdd_port_state_out_3_0_5        ), //i
    .port_i_0_6 (keyAdd_port_state_out_3_0_6        ), //i
    .port_i_0_7 (keyAdd_port_state_out_3_0_7        ), //i
    .port_i_1_0 (keyAdd_port_state_out_3_1_0        ), //i
    .port_i_1_1 (keyAdd_port_state_out_3_1_1        ), //i
    .port_i_1_2 (keyAdd_port_state_out_3_1_2        ), //i
    .port_i_1_3 (keyAdd_port_state_out_3_1_3        ), //i
    .port_i_1_4 (keyAdd_port_state_out_3_1_4        ), //i
    .port_i_1_5 (keyAdd_port_state_out_3_1_5        ), //i
    .port_i_1_6 (keyAdd_port_state_out_3_1_6        ), //i
    .port_i_1_7 (keyAdd_port_state_out_3_1_7        ), //i
    .port_i_2_0 (keyAdd_port_state_out_3_2_0        ), //i
    .port_i_2_1 (keyAdd_port_state_out_3_2_1        ), //i
    .port_i_2_2 (keyAdd_port_state_out_3_2_2        ), //i
    .port_i_2_3 (keyAdd_port_state_out_3_2_3        ), //i
    .port_i_2_4 (keyAdd_port_state_out_3_2_4        ), //i
    .port_i_2_5 (keyAdd_port_state_out_3_2_5        ), //i
    .port_i_2_6 (keyAdd_port_state_out_3_2_6        ), //i
    .port_i_2_7 (keyAdd_port_state_out_3_2_7        ), //i
    .port_i_3_0 (keyAdd_port_state_out_3_3_0        ), //i
    .port_i_3_1 (keyAdd_port_state_out_3_3_1        ), //i
    .port_i_3_2 (keyAdd_port_state_out_3_3_2        ), //i
    .port_i_3_3 (keyAdd_port_state_out_3_3_3        ), //i
    .port_i_3_4 (keyAdd_port_state_out_3_3_4        ), //i
    .port_i_3_5 (keyAdd_port_state_out_3_3_5        ), //i
    .port_i_3_6 (keyAdd_port_state_out_3_3_6        ), //i
    .port_i_3_7 (keyAdd_port_state_out_3_3_7        ), //i
    .port_o_0_0 (sbox_AES_BoyarPeralta_19_port_o_0_0), //o
    .port_o_0_1 (sbox_AES_BoyarPeralta_19_port_o_0_1), //o
    .port_o_0_2 (sbox_AES_BoyarPeralta_19_port_o_0_2), //o
    .port_o_0_3 (sbox_AES_BoyarPeralta_19_port_o_0_3), //o
    .port_o_0_4 (sbox_AES_BoyarPeralta_19_port_o_0_4), //o
    .port_o_0_5 (sbox_AES_BoyarPeralta_19_port_o_0_5), //o
    .port_o_0_6 (sbox_AES_BoyarPeralta_19_port_o_0_6), //o
    .port_o_0_7 (sbox_AES_BoyarPeralta_19_port_o_0_7), //o
    .port_o_1_0 (sbox_AES_BoyarPeralta_19_port_o_1_0), //o
    .port_o_1_1 (sbox_AES_BoyarPeralta_19_port_o_1_1), //o
    .port_o_1_2 (sbox_AES_BoyarPeralta_19_port_o_1_2), //o
    .port_o_1_3 (sbox_AES_BoyarPeralta_19_port_o_1_3), //o
    .port_o_1_4 (sbox_AES_BoyarPeralta_19_port_o_1_4), //o
    .port_o_1_5 (sbox_AES_BoyarPeralta_19_port_o_1_5), //o
    .port_o_1_6 (sbox_AES_BoyarPeralta_19_port_o_1_6), //o
    .port_o_1_7 (sbox_AES_BoyarPeralta_19_port_o_1_7), //o
    .port_o_2_0 (sbox_AES_BoyarPeralta_19_port_o_2_0), //o
    .port_o_2_1 (sbox_AES_BoyarPeralta_19_port_o_2_1), //o
    .port_o_2_2 (sbox_AES_BoyarPeralta_19_port_o_2_2), //o
    .port_o_2_3 (sbox_AES_BoyarPeralta_19_port_o_2_3), //o
    .port_o_2_4 (sbox_AES_BoyarPeralta_19_port_o_2_4), //o
    .port_o_2_5 (sbox_AES_BoyarPeralta_19_port_o_2_5), //o
    .port_o_2_6 (sbox_AES_BoyarPeralta_19_port_o_2_6), //o
    .port_o_2_7 (sbox_AES_BoyarPeralta_19_port_o_2_7), //o
    .port_o_3_0 (sbox_AES_BoyarPeralta_19_port_o_3_0), //o
    .port_o_3_1 (sbox_AES_BoyarPeralta_19_port_o_3_1), //o
    .port_o_3_2 (sbox_AES_BoyarPeralta_19_port_o_3_2), //o
    .port_o_3_3 (sbox_AES_BoyarPeralta_19_port_o_3_3), //o
    .port_o_3_4 (sbox_AES_BoyarPeralta_19_port_o_3_4), //o
    .port_o_3_5 (sbox_AES_BoyarPeralta_19_port_o_3_5), //o
    .port_o_3_6 (sbox_AES_BoyarPeralta_19_port_o_3_6), //o
    .port_o_3_7 (sbox_AES_BoyarPeralta_19_port_o_3_7), //o
    .clk        (clk                                ), //i
    .reset      (reset                              )  //i
  );
  Sbox_AES_BoyarPeralta sbox_AES_BoyarPeralta_20 (
    .port_i_0_0 (keyAdd_port_state_out_4_0_0        ), //i
    .port_i_0_1 (keyAdd_port_state_out_4_0_1        ), //i
    .port_i_0_2 (keyAdd_port_state_out_4_0_2        ), //i
    .port_i_0_3 (keyAdd_port_state_out_4_0_3        ), //i
    .port_i_0_4 (keyAdd_port_state_out_4_0_4        ), //i
    .port_i_0_5 (keyAdd_port_state_out_4_0_5        ), //i
    .port_i_0_6 (keyAdd_port_state_out_4_0_6        ), //i
    .port_i_0_7 (keyAdd_port_state_out_4_0_7        ), //i
    .port_i_1_0 (keyAdd_port_state_out_4_1_0        ), //i
    .port_i_1_1 (keyAdd_port_state_out_4_1_1        ), //i
    .port_i_1_2 (keyAdd_port_state_out_4_1_2        ), //i
    .port_i_1_3 (keyAdd_port_state_out_4_1_3        ), //i
    .port_i_1_4 (keyAdd_port_state_out_4_1_4        ), //i
    .port_i_1_5 (keyAdd_port_state_out_4_1_5        ), //i
    .port_i_1_6 (keyAdd_port_state_out_4_1_6        ), //i
    .port_i_1_7 (keyAdd_port_state_out_4_1_7        ), //i
    .port_i_2_0 (keyAdd_port_state_out_4_2_0        ), //i
    .port_i_2_1 (keyAdd_port_state_out_4_2_1        ), //i
    .port_i_2_2 (keyAdd_port_state_out_4_2_2        ), //i
    .port_i_2_3 (keyAdd_port_state_out_4_2_3        ), //i
    .port_i_2_4 (keyAdd_port_state_out_4_2_4        ), //i
    .port_i_2_5 (keyAdd_port_state_out_4_2_5        ), //i
    .port_i_2_6 (keyAdd_port_state_out_4_2_6        ), //i
    .port_i_2_7 (keyAdd_port_state_out_4_2_7        ), //i
    .port_i_3_0 (keyAdd_port_state_out_4_3_0        ), //i
    .port_i_3_1 (keyAdd_port_state_out_4_3_1        ), //i
    .port_i_3_2 (keyAdd_port_state_out_4_3_2        ), //i
    .port_i_3_3 (keyAdd_port_state_out_4_3_3        ), //i
    .port_i_3_4 (keyAdd_port_state_out_4_3_4        ), //i
    .port_i_3_5 (keyAdd_port_state_out_4_3_5        ), //i
    .port_i_3_6 (keyAdd_port_state_out_4_3_6        ), //i
    .port_i_3_7 (keyAdd_port_state_out_4_3_7        ), //i
    .port_o_0_0 (sbox_AES_BoyarPeralta_20_port_o_0_0), //o
    .port_o_0_1 (sbox_AES_BoyarPeralta_20_port_o_0_1), //o
    .port_o_0_2 (sbox_AES_BoyarPeralta_20_port_o_0_2), //o
    .port_o_0_3 (sbox_AES_BoyarPeralta_20_port_o_0_3), //o
    .port_o_0_4 (sbox_AES_BoyarPeralta_20_port_o_0_4), //o
    .port_o_0_5 (sbox_AES_BoyarPeralta_20_port_o_0_5), //o
    .port_o_0_6 (sbox_AES_BoyarPeralta_20_port_o_0_6), //o
    .port_o_0_7 (sbox_AES_BoyarPeralta_20_port_o_0_7), //o
    .port_o_1_0 (sbox_AES_BoyarPeralta_20_port_o_1_0), //o
    .port_o_1_1 (sbox_AES_BoyarPeralta_20_port_o_1_1), //o
    .port_o_1_2 (sbox_AES_BoyarPeralta_20_port_o_1_2), //o
    .port_o_1_3 (sbox_AES_BoyarPeralta_20_port_o_1_3), //o
    .port_o_1_4 (sbox_AES_BoyarPeralta_20_port_o_1_4), //o
    .port_o_1_5 (sbox_AES_BoyarPeralta_20_port_o_1_5), //o
    .port_o_1_6 (sbox_AES_BoyarPeralta_20_port_o_1_6), //o
    .port_o_1_7 (sbox_AES_BoyarPeralta_20_port_o_1_7), //o
    .port_o_2_0 (sbox_AES_BoyarPeralta_20_port_o_2_0), //o
    .port_o_2_1 (sbox_AES_BoyarPeralta_20_port_o_2_1), //o
    .port_o_2_2 (sbox_AES_BoyarPeralta_20_port_o_2_2), //o
    .port_o_2_3 (sbox_AES_BoyarPeralta_20_port_o_2_3), //o
    .port_o_2_4 (sbox_AES_BoyarPeralta_20_port_o_2_4), //o
    .port_o_2_5 (sbox_AES_BoyarPeralta_20_port_o_2_5), //o
    .port_o_2_6 (sbox_AES_BoyarPeralta_20_port_o_2_6), //o
    .port_o_2_7 (sbox_AES_BoyarPeralta_20_port_o_2_7), //o
    .port_o_3_0 (sbox_AES_BoyarPeralta_20_port_o_3_0), //o
    .port_o_3_1 (sbox_AES_BoyarPeralta_20_port_o_3_1), //o
    .port_o_3_2 (sbox_AES_BoyarPeralta_20_port_o_3_2), //o
    .port_o_3_3 (sbox_AES_BoyarPeralta_20_port_o_3_3), //o
    .port_o_3_4 (sbox_AES_BoyarPeralta_20_port_o_3_4), //o
    .port_o_3_5 (sbox_AES_BoyarPeralta_20_port_o_3_5), //o
    .port_o_3_6 (sbox_AES_BoyarPeralta_20_port_o_3_6), //o
    .port_o_3_7 (sbox_AES_BoyarPeralta_20_port_o_3_7), //o
    .clk        (clk                                ), //i
    .reset      (reset                              )  //i
  );
  Sbox_AES_BoyarPeralta sbox_AES_BoyarPeralta_21 (
    .port_i_0_0 (keyAdd_port_state_out_5_0_0        ), //i
    .port_i_0_1 (keyAdd_port_state_out_5_0_1        ), //i
    .port_i_0_2 (keyAdd_port_state_out_5_0_2        ), //i
    .port_i_0_3 (keyAdd_port_state_out_5_0_3        ), //i
    .port_i_0_4 (keyAdd_port_state_out_5_0_4        ), //i
    .port_i_0_5 (keyAdd_port_state_out_5_0_5        ), //i
    .port_i_0_6 (keyAdd_port_state_out_5_0_6        ), //i
    .port_i_0_7 (keyAdd_port_state_out_5_0_7        ), //i
    .port_i_1_0 (keyAdd_port_state_out_5_1_0        ), //i
    .port_i_1_1 (keyAdd_port_state_out_5_1_1        ), //i
    .port_i_1_2 (keyAdd_port_state_out_5_1_2        ), //i
    .port_i_1_3 (keyAdd_port_state_out_5_1_3        ), //i
    .port_i_1_4 (keyAdd_port_state_out_5_1_4        ), //i
    .port_i_1_5 (keyAdd_port_state_out_5_1_5        ), //i
    .port_i_1_6 (keyAdd_port_state_out_5_1_6        ), //i
    .port_i_1_7 (keyAdd_port_state_out_5_1_7        ), //i
    .port_i_2_0 (keyAdd_port_state_out_5_2_0        ), //i
    .port_i_2_1 (keyAdd_port_state_out_5_2_1        ), //i
    .port_i_2_2 (keyAdd_port_state_out_5_2_2        ), //i
    .port_i_2_3 (keyAdd_port_state_out_5_2_3        ), //i
    .port_i_2_4 (keyAdd_port_state_out_5_2_4        ), //i
    .port_i_2_5 (keyAdd_port_state_out_5_2_5        ), //i
    .port_i_2_6 (keyAdd_port_state_out_5_2_6        ), //i
    .port_i_2_7 (keyAdd_port_state_out_5_2_7        ), //i
    .port_i_3_0 (keyAdd_port_state_out_5_3_0        ), //i
    .port_i_3_1 (keyAdd_port_state_out_5_3_1        ), //i
    .port_i_3_2 (keyAdd_port_state_out_5_3_2        ), //i
    .port_i_3_3 (keyAdd_port_state_out_5_3_3        ), //i
    .port_i_3_4 (keyAdd_port_state_out_5_3_4        ), //i
    .port_i_3_5 (keyAdd_port_state_out_5_3_5        ), //i
    .port_i_3_6 (keyAdd_port_state_out_5_3_6        ), //i
    .port_i_3_7 (keyAdd_port_state_out_5_3_7        ), //i
    .port_o_0_0 (sbox_AES_BoyarPeralta_21_port_o_0_0), //o
    .port_o_0_1 (sbox_AES_BoyarPeralta_21_port_o_0_1), //o
    .port_o_0_2 (sbox_AES_BoyarPeralta_21_port_o_0_2), //o
    .port_o_0_3 (sbox_AES_BoyarPeralta_21_port_o_0_3), //o
    .port_o_0_4 (sbox_AES_BoyarPeralta_21_port_o_0_4), //o
    .port_o_0_5 (sbox_AES_BoyarPeralta_21_port_o_0_5), //o
    .port_o_0_6 (sbox_AES_BoyarPeralta_21_port_o_0_6), //o
    .port_o_0_7 (sbox_AES_BoyarPeralta_21_port_o_0_7), //o
    .port_o_1_0 (sbox_AES_BoyarPeralta_21_port_o_1_0), //o
    .port_o_1_1 (sbox_AES_BoyarPeralta_21_port_o_1_1), //o
    .port_o_1_2 (sbox_AES_BoyarPeralta_21_port_o_1_2), //o
    .port_o_1_3 (sbox_AES_BoyarPeralta_21_port_o_1_3), //o
    .port_o_1_4 (sbox_AES_BoyarPeralta_21_port_o_1_4), //o
    .port_o_1_5 (sbox_AES_BoyarPeralta_21_port_o_1_5), //o
    .port_o_1_6 (sbox_AES_BoyarPeralta_21_port_o_1_6), //o
    .port_o_1_7 (sbox_AES_BoyarPeralta_21_port_o_1_7), //o
    .port_o_2_0 (sbox_AES_BoyarPeralta_21_port_o_2_0), //o
    .port_o_2_1 (sbox_AES_BoyarPeralta_21_port_o_2_1), //o
    .port_o_2_2 (sbox_AES_BoyarPeralta_21_port_o_2_2), //o
    .port_o_2_3 (sbox_AES_BoyarPeralta_21_port_o_2_3), //o
    .port_o_2_4 (sbox_AES_BoyarPeralta_21_port_o_2_4), //o
    .port_o_2_5 (sbox_AES_BoyarPeralta_21_port_o_2_5), //o
    .port_o_2_6 (sbox_AES_BoyarPeralta_21_port_o_2_6), //o
    .port_o_2_7 (sbox_AES_BoyarPeralta_21_port_o_2_7), //o
    .port_o_3_0 (sbox_AES_BoyarPeralta_21_port_o_3_0), //o
    .port_o_3_1 (sbox_AES_BoyarPeralta_21_port_o_3_1), //o
    .port_o_3_2 (sbox_AES_BoyarPeralta_21_port_o_3_2), //o
    .port_o_3_3 (sbox_AES_BoyarPeralta_21_port_o_3_3), //o
    .port_o_3_4 (sbox_AES_BoyarPeralta_21_port_o_3_4), //o
    .port_o_3_5 (sbox_AES_BoyarPeralta_21_port_o_3_5), //o
    .port_o_3_6 (sbox_AES_BoyarPeralta_21_port_o_3_6), //o
    .port_o_3_7 (sbox_AES_BoyarPeralta_21_port_o_3_7), //o
    .clk        (clk                                ), //i
    .reset      (reset                              )  //i
  );
  Sbox_AES_BoyarPeralta sbox_AES_BoyarPeralta_22 (
    .port_i_0_0 (keyAdd_port_state_out_6_0_0        ), //i
    .port_i_0_1 (keyAdd_port_state_out_6_0_1        ), //i
    .port_i_0_2 (keyAdd_port_state_out_6_0_2        ), //i
    .port_i_0_3 (keyAdd_port_state_out_6_0_3        ), //i
    .port_i_0_4 (keyAdd_port_state_out_6_0_4        ), //i
    .port_i_0_5 (keyAdd_port_state_out_6_0_5        ), //i
    .port_i_0_6 (keyAdd_port_state_out_6_0_6        ), //i
    .port_i_0_7 (keyAdd_port_state_out_6_0_7        ), //i
    .port_i_1_0 (keyAdd_port_state_out_6_1_0        ), //i
    .port_i_1_1 (keyAdd_port_state_out_6_1_1        ), //i
    .port_i_1_2 (keyAdd_port_state_out_6_1_2        ), //i
    .port_i_1_3 (keyAdd_port_state_out_6_1_3        ), //i
    .port_i_1_4 (keyAdd_port_state_out_6_1_4        ), //i
    .port_i_1_5 (keyAdd_port_state_out_6_1_5        ), //i
    .port_i_1_6 (keyAdd_port_state_out_6_1_6        ), //i
    .port_i_1_7 (keyAdd_port_state_out_6_1_7        ), //i
    .port_i_2_0 (keyAdd_port_state_out_6_2_0        ), //i
    .port_i_2_1 (keyAdd_port_state_out_6_2_1        ), //i
    .port_i_2_2 (keyAdd_port_state_out_6_2_2        ), //i
    .port_i_2_3 (keyAdd_port_state_out_6_2_3        ), //i
    .port_i_2_4 (keyAdd_port_state_out_6_2_4        ), //i
    .port_i_2_5 (keyAdd_port_state_out_6_2_5        ), //i
    .port_i_2_6 (keyAdd_port_state_out_6_2_6        ), //i
    .port_i_2_7 (keyAdd_port_state_out_6_2_7        ), //i
    .port_i_3_0 (keyAdd_port_state_out_6_3_0        ), //i
    .port_i_3_1 (keyAdd_port_state_out_6_3_1        ), //i
    .port_i_3_2 (keyAdd_port_state_out_6_3_2        ), //i
    .port_i_3_3 (keyAdd_port_state_out_6_3_3        ), //i
    .port_i_3_4 (keyAdd_port_state_out_6_3_4        ), //i
    .port_i_3_5 (keyAdd_port_state_out_6_3_5        ), //i
    .port_i_3_6 (keyAdd_port_state_out_6_3_6        ), //i
    .port_i_3_7 (keyAdd_port_state_out_6_3_7        ), //i
    .port_o_0_0 (sbox_AES_BoyarPeralta_22_port_o_0_0), //o
    .port_o_0_1 (sbox_AES_BoyarPeralta_22_port_o_0_1), //o
    .port_o_0_2 (sbox_AES_BoyarPeralta_22_port_o_0_2), //o
    .port_o_0_3 (sbox_AES_BoyarPeralta_22_port_o_0_3), //o
    .port_o_0_4 (sbox_AES_BoyarPeralta_22_port_o_0_4), //o
    .port_o_0_5 (sbox_AES_BoyarPeralta_22_port_o_0_5), //o
    .port_o_0_6 (sbox_AES_BoyarPeralta_22_port_o_0_6), //o
    .port_o_0_7 (sbox_AES_BoyarPeralta_22_port_o_0_7), //o
    .port_o_1_0 (sbox_AES_BoyarPeralta_22_port_o_1_0), //o
    .port_o_1_1 (sbox_AES_BoyarPeralta_22_port_o_1_1), //o
    .port_o_1_2 (sbox_AES_BoyarPeralta_22_port_o_1_2), //o
    .port_o_1_3 (sbox_AES_BoyarPeralta_22_port_o_1_3), //o
    .port_o_1_4 (sbox_AES_BoyarPeralta_22_port_o_1_4), //o
    .port_o_1_5 (sbox_AES_BoyarPeralta_22_port_o_1_5), //o
    .port_o_1_6 (sbox_AES_BoyarPeralta_22_port_o_1_6), //o
    .port_o_1_7 (sbox_AES_BoyarPeralta_22_port_o_1_7), //o
    .port_o_2_0 (sbox_AES_BoyarPeralta_22_port_o_2_0), //o
    .port_o_2_1 (sbox_AES_BoyarPeralta_22_port_o_2_1), //o
    .port_o_2_2 (sbox_AES_BoyarPeralta_22_port_o_2_2), //o
    .port_o_2_3 (sbox_AES_BoyarPeralta_22_port_o_2_3), //o
    .port_o_2_4 (sbox_AES_BoyarPeralta_22_port_o_2_4), //o
    .port_o_2_5 (sbox_AES_BoyarPeralta_22_port_o_2_5), //o
    .port_o_2_6 (sbox_AES_BoyarPeralta_22_port_o_2_6), //o
    .port_o_2_7 (sbox_AES_BoyarPeralta_22_port_o_2_7), //o
    .port_o_3_0 (sbox_AES_BoyarPeralta_22_port_o_3_0), //o
    .port_o_3_1 (sbox_AES_BoyarPeralta_22_port_o_3_1), //o
    .port_o_3_2 (sbox_AES_BoyarPeralta_22_port_o_3_2), //o
    .port_o_3_3 (sbox_AES_BoyarPeralta_22_port_o_3_3), //o
    .port_o_3_4 (sbox_AES_BoyarPeralta_22_port_o_3_4), //o
    .port_o_3_5 (sbox_AES_BoyarPeralta_22_port_o_3_5), //o
    .port_o_3_6 (sbox_AES_BoyarPeralta_22_port_o_3_6), //o
    .port_o_3_7 (sbox_AES_BoyarPeralta_22_port_o_3_7), //o
    .clk        (clk                                ), //i
    .reset      (reset                              )  //i
  );
  Sbox_AES_BoyarPeralta sbox_AES_BoyarPeralta_23 (
    .port_i_0_0 (keyAdd_port_state_out_7_0_0        ), //i
    .port_i_0_1 (keyAdd_port_state_out_7_0_1        ), //i
    .port_i_0_2 (keyAdd_port_state_out_7_0_2        ), //i
    .port_i_0_3 (keyAdd_port_state_out_7_0_3        ), //i
    .port_i_0_4 (keyAdd_port_state_out_7_0_4        ), //i
    .port_i_0_5 (keyAdd_port_state_out_7_0_5        ), //i
    .port_i_0_6 (keyAdd_port_state_out_7_0_6        ), //i
    .port_i_0_7 (keyAdd_port_state_out_7_0_7        ), //i
    .port_i_1_0 (keyAdd_port_state_out_7_1_0        ), //i
    .port_i_1_1 (keyAdd_port_state_out_7_1_1        ), //i
    .port_i_1_2 (keyAdd_port_state_out_7_1_2        ), //i
    .port_i_1_3 (keyAdd_port_state_out_7_1_3        ), //i
    .port_i_1_4 (keyAdd_port_state_out_7_1_4        ), //i
    .port_i_1_5 (keyAdd_port_state_out_7_1_5        ), //i
    .port_i_1_6 (keyAdd_port_state_out_7_1_6        ), //i
    .port_i_1_7 (keyAdd_port_state_out_7_1_7        ), //i
    .port_i_2_0 (keyAdd_port_state_out_7_2_0        ), //i
    .port_i_2_1 (keyAdd_port_state_out_7_2_1        ), //i
    .port_i_2_2 (keyAdd_port_state_out_7_2_2        ), //i
    .port_i_2_3 (keyAdd_port_state_out_7_2_3        ), //i
    .port_i_2_4 (keyAdd_port_state_out_7_2_4        ), //i
    .port_i_2_5 (keyAdd_port_state_out_7_2_5        ), //i
    .port_i_2_6 (keyAdd_port_state_out_7_2_6        ), //i
    .port_i_2_7 (keyAdd_port_state_out_7_2_7        ), //i
    .port_i_3_0 (keyAdd_port_state_out_7_3_0        ), //i
    .port_i_3_1 (keyAdd_port_state_out_7_3_1        ), //i
    .port_i_3_2 (keyAdd_port_state_out_7_3_2        ), //i
    .port_i_3_3 (keyAdd_port_state_out_7_3_3        ), //i
    .port_i_3_4 (keyAdd_port_state_out_7_3_4        ), //i
    .port_i_3_5 (keyAdd_port_state_out_7_3_5        ), //i
    .port_i_3_6 (keyAdd_port_state_out_7_3_6        ), //i
    .port_i_3_7 (keyAdd_port_state_out_7_3_7        ), //i
    .port_o_0_0 (sbox_AES_BoyarPeralta_23_port_o_0_0), //o
    .port_o_0_1 (sbox_AES_BoyarPeralta_23_port_o_0_1), //o
    .port_o_0_2 (sbox_AES_BoyarPeralta_23_port_o_0_2), //o
    .port_o_0_3 (sbox_AES_BoyarPeralta_23_port_o_0_3), //o
    .port_o_0_4 (sbox_AES_BoyarPeralta_23_port_o_0_4), //o
    .port_o_0_5 (sbox_AES_BoyarPeralta_23_port_o_0_5), //o
    .port_o_0_6 (sbox_AES_BoyarPeralta_23_port_o_0_6), //o
    .port_o_0_7 (sbox_AES_BoyarPeralta_23_port_o_0_7), //o
    .port_o_1_0 (sbox_AES_BoyarPeralta_23_port_o_1_0), //o
    .port_o_1_1 (sbox_AES_BoyarPeralta_23_port_o_1_1), //o
    .port_o_1_2 (sbox_AES_BoyarPeralta_23_port_o_1_2), //o
    .port_o_1_3 (sbox_AES_BoyarPeralta_23_port_o_1_3), //o
    .port_o_1_4 (sbox_AES_BoyarPeralta_23_port_o_1_4), //o
    .port_o_1_5 (sbox_AES_BoyarPeralta_23_port_o_1_5), //o
    .port_o_1_6 (sbox_AES_BoyarPeralta_23_port_o_1_6), //o
    .port_o_1_7 (sbox_AES_BoyarPeralta_23_port_o_1_7), //o
    .port_o_2_0 (sbox_AES_BoyarPeralta_23_port_o_2_0), //o
    .port_o_2_1 (sbox_AES_BoyarPeralta_23_port_o_2_1), //o
    .port_o_2_2 (sbox_AES_BoyarPeralta_23_port_o_2_2), //o
    .port_o_2_3 (sbox_AES_BoyarPeralta_23_port_o_2_3), //o
    .port_o_2_4 (sbox_AES_BoyarPeralta_23_port_o_2_4), //o
    .port_o_2_5 (sbox_AES_BoyarPeralta_23_port_o_2_5), //o
    .port_o_2_6 (sbox_AES_BoyarPeralta_23_port_o_2_6), //o
    .port_o_2_7 (sbox_AES_BoyarPeralta_23_port_o_2_7), //o
    .port_o_3_0 (sbox_AES_BoyarPeralta_23_port_o_3_0), //o
    .port_o_3_1 (sbox_AES_BoyarPeralta_23_port_o_3_1), //o
    .port_o_3_2 (sbox_AES_BoyarPeralta_23_port_o_3_2), //o
    .port_o_3_3 (sbox_AES_BoyarPeralta_23_port_o_3_3), //o
    .port_o_3_4 (sbox_AES_BoyarPeralta_23_port_o_3_4), //o
    .port_o_3_5 (sbox_AES_BoyarPeralta_23_port_o_3_5), //o
    .port_o_3_6 (sbox_AES_BoyarPeralta_23_port_o_3_6), //o
    .port_o_3_7 (sbox_AES_BoyarPeralta_23_port_o_3_7), //o
    .clk        (clk                                ), //i
    .reset      (reset                              )  //i
  );
  Sbox_AES_BoyarPeralta sbox_AES_BoyarPeralta_24 (
    .port_i_0_0 (keyAdd_port_state_out_8_0_0        ), //i
    .port_i_0_1 (keyAdd_port_state_out_8_0_1        ), //i
    .port_i_0_2 (keyAdd_port_state_out_8_0_2        ), //i
    .port_i_0_3 (keyAdd_port_state_out_8_0_3        ), //i
    .port_i_0_4 (keyAdd_port_state_out_8_0_4        ), //i
    .port_i_0_5 (keyAdd_port_state_out_8_0_5        ), //i
    .port_i_0_6 (keyAdd_port_state_out_8_0_6        ), //i
    .port_i_0_7 (keyAdd_port_state_out_8_0_7        ), //i
    .port_i_1_0 (keyAdd_port_state_out_8_1_0        ), //i
    .port_i_1_1 (keyAdd_port_state_out_8_1_1        ), //i
    .port_i_1_2 (keyAdd_port_state_out_8_1_2        ), //i
    .port_i_1_3 (keyAdd_port_state_out_8_1_3        ), //i
    .port_i_1_4 (keyAdd_port_state_out_8_1_4        ), //i
    .port_i_1_5 (keyAdd_port_state_out_8_1_5        ), //i
    .port_i_1_6 (keyAdd_port_state_out_8_1_6        ), //i
    .port_i_1_7 (keyAdd_port_state_out_8_1_7        ), //i
    .port_i_2_0 (keyAdd_port_state_out_8_2_0        ), //i
    .port_i_2_1 (keyAdd_port_state_out_8_2_1        ), //i
    .port_i_2_2 (keyAdd_port_state_out_8_2_2        ), //i
    .port_i_2_3 (keyAdd_port_state_out_8_2_3        ), //i
    .port_i_2_4 (keyAdd_port_state_out_8_2_4        ), //i
    .port_i_2_5 (keyAdd_port_state_out_8_2_5        ), //i
    .port_i_2_6 (keyAdd_port_state_out_8_2_6        ), //i
    .port_i_2_7 (keyAdd_port_state_out_8_2_7        ), //i
    .port_i_3_0 (keyAdd_port_state_out_8_3_0        ), //i
    .port_i_3_1 (keyAdd_port_state_out_8_3_1        ), //i
    .port_i_3_2 (keyAdd_port_state_out_8_3_2        ), //i
    .port_i_3_3 (keyAdd_port_state_out_8_3_3        ), //i
    .port_i_3_4 (keyAdd_port_state_out_8_3_4        ), //i
    .port_i_3_5 (keyAdd_port_state_out_8_3_5        ), //i
    .port_i_3_6 (keyAdd_port_state_out_8_3_6        ), //i
    .port_i_3_7 (keyAdd_port_state_out_8_3_7        ), //i
    .port_o_0_0 (sbox_AES_BoyarPeralta_24_port_o_0_0), //o
    .port_o_0_1 (sbox_AES_BoyarPeralta_24_port_o_0_1), //o
    .port_o_0_2 (sbox_AES_BoyarPeralta_24_port_o_0_2), //o
    .port_o_0_3 (sbox_AES_BoyarPeralta_24_port_o_0_3), //o
    .port_o_0_4 (sbox_AES_BoyarPeralta_24_port_o_0_4), //o
    .port_o_0_5 (sbox_AES_BoyarPeralta_24_port_o_0_5), //o
    .port_o_0_6 (sbox_AES_BoyarPeralta_24_port_o_0_6), //o
    .port_o_0_7 (sbox_AES_BoyarPeralta_24_port_o_0_7), //o
    .port_o_1_0 (sbox_AES_BoyarPeralta_24_port_o_1_0), //o
    .port_o_1_1 (sbox_AES_BoyarPeralta_24_port_o_1_1), //o
    .port_o_1_2 (sbox_AES_BoyarPeralta_24_port_o_1_2), //o
    .port_o_1_3 (sbox_AES_BoyarPeralta_24_port_o_1_3), //o
    .port_o_1_4 (sbox_AES_BoyarPeralta_24_port_o_1_4), //o
    .port_o_1_5 (sbox_AES_BoyarPeralta_24_port_o_1_5), //o
    .port_o_1_6 (sbox_AES_BoyarPeralta_24_port_o_1_6), //o
    .port_o_1_7 (sbox_AES_BoyarPeralta_24_port_o_1_7), //o
    .port_o_2_0 (sbox_AES_BoyarPeralta_24_port_o_2_0), //o
    .port_o_2_1 (sbox_AES_BoyarPeralta_24_port_o_2_1), //o
    .port_o_2_2 (sbox_AES_BoyarPeralta_24_port_o_2_2), //o
    .port_o_2_3 (sbox_AES_BoyarPeralta_24_port_o_2_3), //o
    .port_o_2_4 (sbox_AES_BoyarPeralta_24_port_o_2_4), //o
    .port_o_2_5 (sbox_AES_BoyarPeralta_24_port_o_2_5), //o
    .port_o_2_6 (sbox_AES_BoyarPeralta_24_port_o_2_6), //o
    .port_o_2_7 (sbox_AES_BoyarPeralta_24_port_o_2_7), //o
    .port_o_3_0 (sbox_AES_BoyarPeralta_24_port_o_3_0), //o
    .port_o_3_1 (sbox_AES_BoyarPeralta_24_port_o_3_1), //o
    .port_o_3_2 (sbox_AES_BoyarPeralta_24_port_o_3_2), //o
    .port_o_3_3 (sbox_AES_BoyarPeralta_24_port_o_3_3), //o
    .port_o_3_4 (sbox_AES_BoyarPeralta_24_port_o_3_4), //o
    .port_o_3_5 (sbox_AES_BoyarPeralta_24_port_o_3_5), //o
    .port_o_3_6 (sbox_AES_BoyarPeralta_24_port_o_3_6), //o
    .port_o_3_7 (sbox_AES_BoyarPeralta_24_port_o_3_7), //o
    .clk        (clk                                ), //i
    .reset      (reset                              )  //i
  );
  Sbox_AES_BoyarPeralta sbox_AES_BoyarPeralta_25 (
    .port_i_0_0 (keyAdd_port_state_out_9_0_0        ), //i
    .port_i_0_1 (keyAdd_port_state_out_9_0_1        ), //i
    .port_i_0_2 (keyAdd_port_state_out_9_0_2        ), //i
    .port_i_0_3 (keyAdd_port_state_out_9_0_3        ), //i
    .port_i_0_4 (keyAdd_port_state_out_9_0_4        ), //i
    .port_i_0_5 (keyAdd_port_state_out_9_0_5        ), //i
    .port_i_0_6 (keyAdd_port_state_out_9_0_6        ), //i
    .port_i_0_7 (keyAdd_port_state_out_9_0_7        ), //i
    .port_i_1_0 (keyAdd_port_state_out_9_1_0        ), //i
    .port_i_1_1 (keyAdd_port_state_out_9_1_1        ), //i
    .port_i_1_2 (keyAdd_port_state_out_9_1_2        ), //i
    .port_i_1_3 (keyAdd_port_state_out_9_1_3        ), //i
    .port_i_1_4 (keyAdd_port_state_out_9_1_4        ), //i
    .port_i_1_5 (keyAdd_port_state_out_9_1_5        ), //i
    .port_i_1_6 (keyAdd_port_state_out_9_1_6        ), //i
    .port_i_1_7 (keyAdd_port_state_out_9_1_7        ), //i
    .port_i_2_0 (keyAdd_port_state_out_9_2_0        ), //i
    .port_i_2_1 (keyAdd_port_state_out_9_2_1        ), //i
    .port_i_2_2 (keyAdd_port_state_out_9_2_2        ), //i
    .port_i_2_3 (keyAdd_port_state_out_9_2_3        ), //i
    .port_i_2_4 (keyAdd_port_state_out_9_2_4        ), //i
    .port_i_2_5 (keyAdd_port_state_out_9_2_5        ), //i
    .port_i_2_6 (keyAdd_port_state_out_9_2_6        ), //i
    .port_i_2_7 (keyAdd_port_state_out_9_2_7        ), //i
    .port_i_3_0 (keyAdd_port_state_out_9_3_0        ), //i
    .port_i_3_1 (keyAdd_port_state_out_9_3_1        ), //i
    .port_i_3_2 (keyAdd_port_state_out_9_3_2        ), //i
    .port_i_3_3 (keyAdd_port_state_out_9_3_3        ), //i
    .port_i_3_4 (keyAdd_port_state_out_9_3_4        ), //i
    .port_i_3_5 (keyAdd_port_state_out_9_3_5        ), //i
    .port_i_3_6 (keyAdd_port_state_out_9_3_6        ), //i
    .port_i_3_7 (keyAdd_port_state_out_9_3_7        ), //i
    .port_o_0_0 (sbox_AES_BoyarPeralta_25_port_o_0_0), //o
    .port_o_0_1 (sbox_AES_BoyarPeralta_25_port_o_0_1), //o
    .port_o_0_2 (sbox_AES_BoyarPeralta_25_port_o_0_2), //o
    .port_o_0_3 (sbox_AES_BoyarPeralta_25_port_o_0_3), //o
    .port_o_0_4 (sbox_AES_BoyarPeralta_25_port_o_0_4), //o
    .port_o_0_5 (sbox_AES_BoyarPeralta_25_port_o_0_5), //o
    .port_o_0_6 (sbox_AES_BoyarPeralta_25_port_o_0_6), //o
    .port_o_0_7 (sbox_AES_BoyarPeralta_25_port_o_0_7), //o
    .port_o_1_0 (sbox_AES_BoyarPeralta_25_port_o_1_0), //o
    .port_o_1_1 (sbox_AES_BoyarPeralta_25_port_o_1_1), //o
    .port_o_1_2 (sbox_AES_BoyarPeralta_25_port_o_1_2), //o
    .port_o_1_3 (sbox_AES_BoyarPeralta_25_port_o_1_3), //o
    .port_o_1_4 (sbox_AES_BoyarPeralta_25_port_o_1_4), //o
    .port_o_1_5 (sbox_AES_BoyarPeralta_25_port_o_1_5), //o
    .port_o_1_6 (sbox_AES_BoyarPeralta_25_port_o_1_6), //o
    .port_o_1_7 (sbox_AES_BoyarPeralta_25_port_o_1_7), //o
    .port_o_2_0 (sbox_AES_BoyarPeralta_25_port_o_2_0), //o
    .port_o_2_1 (sbox_AES_BoyarPeralta_25_port_o_2_1), //o
    .port_o_2_2 (sbox_AES_BoyarPeralta_25_port_o_2_2), //o
    .port_o_2_3 (sbox_AES_BoyarPeralta_25_port_o_2_3), //o
    .port_o_2_4 (sbox_AES_BoyarPeralta_25_port_o_2_4), //o
    .port_o_2_5 (sbox_AES_BoyarPeralta_25_port_o_2_5), //o
    .port_o_2_6 (sbox_AES_BoyarPeralta_25_port_o_2_6), //o
    .port_o_2_7 (sbox_AES_BoyarPeralta_25_port_o_2_7), //o
    .port_o_3_0 (sbox_AES_BoyarPeralta_25_port_o_3_0), //o
    .port_o_3_1 (sbox_AES_BoyarPeralta_25_port_o_3_1), //o
    .port_o_3_2 (sbox_AES_BoyarPeralta_25_port_o_3_2), //o
    .port_o_3_3 (sbox_AES_BoyarPeralta_25_port_o_3_3), //o
    .port_o_3_4 (sbox_AES_BoyarPeralta_25_port_o_3_4), //o
    .port_o_3_5 (sbox_AES_BoyarPeralta_25_port_o_3_5), //o
    .port_o_3_6 (sbox_AES_BoyarPeralta_25_port_o_3_6), //o
    .port_o_3_7 (sbox_AES_BoyarPeralta_25_port_o_3_7), //o
    .clk        (clk                                ), //i
    .reset      (reset                              )  //i
  );
  Sbox_AES_BoyarPeralta sbox_AES_BoyarPeralta_26 (
    .port_i_0_0 (keyAdd_port_state_out_10_0_0       ), //i
    .port_i_0_1 (keyAdd_port_state_out_10_0_1       ), //i
    .port_i_0_2 (keyAdd_port_state_out_10_0_2       ), //i
    .port_i_0_3 (keyAdd_port_state_out_10_0_3       ), //i
    .port_i_0_4 (keyAdd_port_state_out_10_0_4       ), //i
    .port_i_0_5 (keyAdd_port_state_out_10_0_5       ), //i
    .port_i_0_6 (keyAdd_port_state_out_10_0_6       ), //i
    .port_i_0_7 (keyAdd_port_state_out_10_0_7       ), //i
    .port_i_1_0 (keyAdd_port_state_out_10_1_0       ), //i
    .port_i_1_1 (keyAdd_port_state_out_10_1_1       ), //i
    .port_i_1_2 (keyAdd_port_state_out_10_1_2       ), //i
    .port_i_1_3 (keyAdd_port_state_out_10_1_3       ), //i
    .port_i_1_4 (keyAdd_port_state_out_10_1_4       ), //i
    .port_i_1_5 (keyAdd_port_state_out_10_1_5       ), //i
    .port_i_1_6 (keyAdd_port_state_out_10_1_6       ), //i
    .port_i_1_7 (keyAdd_port_state_out_10_1_7       ), //i
    .port_i_2_0 (keyAdd_port_state_out_10_2_0       ), //i
    .port_i_2_1 (keyAdd_port_state_out_10_2_1       ), //i
    .port_i_2_2 (keyAdd_port_state_out_10_2_2       ), //i
    .port_i_2_3 (keyAdd_port_state_out_10_2_3       ), //i
    .port_i_2_4 (keyAdd_port_state_out_10_2_4       ), //i
    .port_i_2_5 (keyAdd_port_state_out_10_2_5       ), //i
    .port_i_2_6 (keyAdd_port_state_out_10_2_6       ), //i
    .port_i_2_7 (keyAdd_port_state_out_10_2_7       ), //i
    .port_i_3_0 (keyAdd_port_state_out_10_3_0       ), //i
    .port_i_3_1 (keyAdd_port_state_out_10_3_1       ), //i
    .port_i_3_2 (keyAdd_port_state_out_10_3_2       ), //i
    .port_i_3_3 (keyAdd_port_state_out_10_3_3       ), //i
    .port_i_3_4 (keyAdd_port_state_out_10_3_4       ), //i
    .port_i_3_5 (keyAdd_port_state_out_10_3_5       ), //i
    .port_i_3_6 (keyAdd_port_state_out_10_3_6       ), //i
    .port_i_3_7 (keyAdd_port_state_out_10_3_7       ), //i
    .port_o_0_0 (sbox_AES_BoyarPeralta_26_port_o_0_0), //o
    .port_o_0_1 (sbox_AES_BoyarPeralta_26_port_o_0_1), //o
    .port_o_0_2 (sbox_AES_BoyarPeralta_26_port_o_0_2), //o
    .port_o_0_3 (sbox_AES_BoyarPeralta_26_port_o_0_3), //o
    .port_o_0_4 (sbox_AES_BoyarPeralta_26_port_o_0_4), //o
    .port_o_0_5 (sbox_AES_BoyarPeralta_26_port_o_0_5), //o
    .port_o_0_6 (sbox_AES_BoyarPeralta_26_port_o_0_6), //o
    .port_o_0_7 (sbox_AES_BoyarPeralta_26_port_o_0_7), //o
    .port_o_1_0 (sbox_AES_BoyarPeralta_26_port_o_1_0), //o
    .port_o_1_1 (sbox_AES_BoyarPeralta_26_port_o_1_1), //o
    .port_o_1_2 (sbox_AES_BoyarPeralta_26_port_o_1_2), //o
    .port_o_1_3 (sbox_AES_BoyarPeralta_26_port_o_1_3), //o
    .port_o_1_4 (sbox_AES_BoyarPeralta_26_port_o_1_4), //o
    .port_o_1_5 (sbox_AES_BoyarPeralta_26_port_o_1_5), //o
    .port_o_1_6 (sbox_AES_BoyarPeralta_26_port_o_1_6), //o
    .port_o_1_7 (sbox_AES_BoyarPeralta_26_port_o_1_7), //o
    .port_o_2_0 (sbox_AES_BoyarPeralta_26_port_o_2_0), //o
    .port_o_2_1 (sbox_AES_BoyarPeralta_26_port_o_2_1), //o
    .port_o_2_2 (sbox_AES_BoyarPeralta_26_port_o_2_2), //o
    .port_o_2_3 (sbox_AES_BoyarPeralta_26_port_o_2_3), //o
    .port_o_2_4 (sbox_AES_BoyarPeralta_26_port_o_2_4), //o
    .port_o_2_5 (sbox_AES_BoyarPeralta_26_port_o_2_5), //o
    .port_o_2_6 (sbox_AES_BoyarPeralta_26_port_o_2_6), //o
    .port_o_2_7 (sbox_AES_BoyarPeralta_26_port_o_2_7), //o
    .port_o_3_0 (sbox_AES_BoyarPeralta_26_port_o_3_0), //o
    .port_o_3_1 (sbox_AES_BoyarPeralta_26_port_o_3_1), //o
    .port_o_3_2 (sbox_AES_BoyarPeralta_26_port_o_3_2), //o
    .port_o_3_3 (sbox_AES_BoyarPeralta_26_port_o_3_3), //o
    .port_o_3_4 (sbox_AES_BoyarPeralta_26_port_o_3_4), //o
    .port_o_3_5 (sbox_AES_BoyarPeralta_26_port_o_3_5), //o
    .port_o_3_6 (sbox_AES_BoyarPeralta_26_port_o_3_6), //o
    .port_o_3_7 (sbox_AES_BoyarPeralta_26_port_o_3_7), //o
    .clk        (clk                                ), //i
    .reset      (reset                              )  //i
  );
  Sbox_AES_BoyarPeralta sbox_AES_BoyarPeralta_27 (
    .port_i_0_0 (keyAdd_port_state_out_11_0_0       ), //i
    .port_i_0_1 (keyAdd_port_state_out_11_0_1       ), //i
    .port_i_0_2 (keyAdd_port_state_out_11_0_2       ), //i
    .port_i_0_3 (keyAdd_port_state_out_11_0_3       ), //i
    .port_i_0_4 (keyAdd_port_state_out_11_0_4       ), //i
    .port_i_0_5 (keyAdd_port_state_out_11_0_5       ), //i
    .port_i_0_6 (keyAdd_port_state_out_11_0_6       ), //i
    .port_i_0_7 (keyAdd_port_state_out_11_0_7       ), //i
    .port_i_1_0 (keyAdd_port_state_out_11_1_0       ), //i
    .port_i_1_1 (keyAdd_port_state_out_11_1_1       ), //i
    .port_i_1_2 (keyAdd_port_state_out_11_1_2       ), //i
    .port_i_1_3 (keyAdd_port_state_out_11_1_3       ), //i
    .port_i_1_4 (keyAdd_port_state_out_11_1_4       ), //i
    .port_i_1_5 (keyAdd_port_state_out_11_1_5       ), //i
    .port_i_1_6 (keyAdd_port_state_out_11_1_6       ), //i
    .port_i_1_7 (keyAdd_port_state_out_11_1_7       ), //i
    .port_i_2_0 (keyAdd_port_state_out_11_2_0       ), //i
    .port_i_2_1 (keyAdd_port_state_out_11_2_1       ), //i
    .port_i_2_2 (keyAdd_port_state_out_11_2_2       ), //i
    .port_i_2_3 (keyAdd_port_state_out_11_2_3       ), //i
    .port_i_2_4 (keyAdd_port_state_out_11_2_4       ), //i
    .port_i_2_5 (keyAdd_port_state_out_11_2_5       ), //i
    .port_i_2_6 (keyAdd_port_state_out_11_2_6       ), //i
    .port_i_2_7 (keyAdd_port_state_out_11_2_7       ), //i
    .port_i_3_0 (keyAdd_port_state_out_11_3_0       ), //i
    .port_i_3_1 (keyAdd_port_state_out_11_3_1       ), //i
    .port_i_3_2 (keyAdd_port_state_out_11_3_2       ), //i
    .port_i_3_3 (keyAdd_port_state_out_11_3_3       ), //i
    .port_i_3_4 (keyAdd_port_state_out_11_3_4       ), //i
    .port_i_3_5 (keyAdd_port_state_out_11_3_5       ), //i
    .port_i_3_6 (keyAdd_port_state_out_11_3_6       ), //i
    .port_i_3_7 (keyAdd_port_state_out_11_3_7       ), //i
    .port_o_0_0 (sbox_AES_BoyarPeralta_27_port_o_0_0), //o
    .port_o_0_1 (sbox_AES_BoyarPeralta_27_port_o_0_1), //o
    .port_o_0_2 (sbox_AES_BoyarPeralta_27_port_o_0_2), //o
    .port_o_0_3 (sbox_AES_BoyarPeralta_27_port_o_0_3), //o
    .port_o_0_4 (sbox_AES_BoyarPeralta_27_port_o_0_4), //o
    .port_o_0_5 (sbox_AES_BoyarPeralta_27_port_o_0_5), //o
    .port_o_0_6 (sbox_AES_BoyarPeralta_27_port_o_0_6), //o
    .port_o_0_7 (sbox_AES_BoyarPeralta_27_port_o_0_7), //o
    .port_o_1_0 (sbox_AES_BoyarPeralta_27_port_o_1_0), //o
    .port_o_1_1 (sbox_AES_BoyarPeralta_27_port_o_1_1), //o
    .port_o_1_2 (sbox_AES_BoyarPeralta_27_port_o_1_2), //o
    .port_o_1_3 (sbox_AES_BoyarPeralta_27_port_o_1_3), //o
    .port_o_1_4 (sbox_AES_BoyarPeralta_27_port_o_1_4), //o
    .port_o_1_5 (sbox_AES_BoyarPeralta_27_port_o_1_5), //o
    .port_o_1_6 (sbox_AES_BoyarPeralta_27_port_o_1_6), //o
    .port_o_1_7 (sbox_AES_BoyarPeralta_27_port_o_1_7), //o
    .port_o_2_0 (sbox_AES_BoyarPeralta_27_port_o_2_0), //o
    .port_o_2_1 (sbox_AES_BoyarPeralta_27_port_o_2_1), //o
    .port_o_2_2 (sbox_AES_BoyarPeralta_27_port_o_2_2), //o
    .port_o_2_3 (sbox_AES_BoyarPeralta_27_port_o_2_3), //o
    .port_o_2_4 (sbox_AES_BoyarPeralta_27_port_o_2_4), //o
    .port_o_2_5 (sbox_AES_BoyarPeralta_27_port_o_2_5), //o
    .port_o_2_6 (sbox_AES_BoyarPeralta_27_port_o_2_6), //o
    .port_o_2_7 (sbox_AES_BoyarPeralta_27_port_o_2_7), //o
    .port_o_3_0 (sbox_AES_BoyarPeralta_27_port_o_3_0), //o
    .port_o_3_1 (sbox_AES_BoyarPeralta_27_port_o_3_1), //o
    .port_o_3_2 (sbox_AES_BoyarPeralta_27_port_o_3_2), //o
    .port_o_3_3 (sbox_AES_BoyarPeralta_27_port_o_3_3), //o
    .port_o_3_4 (sbox_AES_BoyarPeralta_27_port_o_3_4), //o
    .port_o_3_5 (sbox_AES_BoyarPeralta_27_port_o_3_5), //o
    .port_o_3_6 (sbox_AES_BoyarPeralta_27_port_o_3_6), //o
    .port_o_3_7 (sbox_AES_BoyarPeralta_27_port_o_3_7), //o
    .clk        (clk                                ), //i
    .reset      (reset                              )  //i
  );
  Sbox_AES_BoyarPeralta sbox_AES_BoyarPeralta_28 (
    .port_i_0_0 (keyAdd_port_state_out_12_0_0       ), //i
    .port_i_0_1 (keyAdd_port_state_out_12_0_1       ), //i
    .port_i_0_2 (keyAdd_port_state_out_12_0_2       ), //i
    .port_i_0_3 (keyAdd_port_state_out_12_0_3       ), //i
    .port_i_0_4 (keyAdd_port_state_out_12_0_4       ), //i
    .port_i_0_5 (keyAdd_port_state_out_12_0_5       ), //i
    .port_i_0_6 (keyAdd_port_state_out_12_0_6       ), //i
    .port_i_0_7 (keyAdd_port_state_out_12_0_7       ), //i
    .port_i_1_0 (keyAdd_port_state_out_12_1_0       ), //i
    .port_i_1_1 (keyAdd_port_state_out_12_1_1       ), //i
    .port_i_1_2 (keyAdd_port_state_out_12_1_2       ), //i
    .port_i_1_3 (keyAdd_port_state_out_12_1_3       ), //i
    .port_i_1_4 (keyAdd_port_state_out_12_1_4       ), //i
    .port_i_1_5 (keyAdd_port_state_out_12_1_5       ), //i
    .port_i_1_6 (keyAdd_port_state_out_12_1_6       ), //i
    .port_i_1_7 (keyAdd_port_state_out_12_1_7       ), //i
    .port_i_2_0 (keyAdd_port_state_out_12_2_0       ), //i
    .port_i_2_1 (keyAdd_port_state_out_12_2_1       ), //i
    .port_i_2_2 (keyAdd_port_state_out_12_2_2       ), //i
    .port_i_2_3 (keyAdd_port_state_out_12_2_3       ), //i
    .port_i_2_4 (keyAdd_port_state_out_12_2_4       ), //i
    .port_i_2_5 (keyAdd_port_state_out_12_2_5       ), //i
    .port_i_2_6 (keyAdd_port_state_out_12_2_6       ), //i
    .port_i_2_7 (keyAdd_port_state_out_12_2_7       ), //i
    .port_i_3_0 (keyAdd_port_state_out_12_3_0       ), //i
    .port_i_3_1 (keyAdd_port_state_out_12_3_1       ), //i
    .port_i_3_2 (keyAdd_port_state_out_12_3_2       ), //i
    .port_i_3_3 (keyAdd_port_state_out_12_3_3       ), //i
    .port_i_3_4 (keyAdd_port_state_out_12_3_4       ), //i
    .port_i_3_5 (keyAdd_port_state_out_12_3_5       ), //i
    .port_i_3_6 (keyAdd_port_state_out_12_3_6       ), //i
    .port_i_3_7 (keyAdd_port_state_out_12_3_7       ), //i
    .port_o_0_0 (sbox_AES_BoyarPeralta_28_port_o_0_0), //o
    .port_o_0_1 (sbox_AES_BoyarPeralta_28_port_o_0_1), //o
    .port_o_0_2 (sbox_AES_BoyarPeralta_28_port_o_0_2), //o
    .port_o_0_3 (sbox_AES_BoyarPeralta_28_port_o_0_3), //o
    .port_o_0_4 (sbox_AES_BoyarPeralta_28_port_o_0_4), //o
    .port_o_0_5 (sbox_AES_BoyarPeralta_28_port_o_0_5), //o
    .port_o_0_6 (sbox_AES_BoyarPeralta_28_port_o_0_6), //o
    .port_o_0_7 (sbox_AES_BoyarPeralta_28_port_o_0_7), //o
    .port_o_1_0 (sbox_AES_BoyarPeralta_28_port_o_1_0), //o
    .port_o_1_1 (sbox_AES_BoyarPeralta_28_port_o_1_1), //o
    .port_o_1_2 (sbox_AES_BoyarPeralta_28_port_o_1_2), //o
    .port_o_1_3 (sbox_AES_BoyarPeralta_28_port_o_1_3), //o
    .port_o_1_4 (sbox_AES_BoyarPeralta_28_port_o_1_4), //o
    .port_o_1_5 (sbox_AES_BoyarPeralta_28_port_o_1_5), //o
    .port_o_1_6 (sbox_AES_BoyarPeralta_28_port_o_1_6), //o
    .port_o_1_7 (sbox_AES_BoyarPeralta_28_port_o_1_7), //o
    .port_o_2_0 (sbox_AES_BoyarPeralta_28_port_o_2_0), //o
    .port_o_2_1 (sbox_AES_BoyarPeralta_28_port_o_2_1), //o
    .port_o_2_2 (sbox_AES_BoyarPeralta_28_port_o_2_2), //o
    .port_o_2_3 (sbox_AES_BoyarPeralta_28_port_o_2_3), //o
    .port_o_2_4 (sbox_AES_BoyarPeralta_28_port_o_2_4), //o
    .port_o_2_5 (sbox_AES_BoyarPeralta_28_port_o_2_5), //o
    .port_o_2_6 (sbox_AES_BoyarPeralta_28_port_o_2_6), //o
    .port_o_2_7 (sbox_AES_BoyarPeralta_28_port_o_2_7), //o
    .port_o_3_0 (sbox_AES_BoyarPeralta_28_port_o_3_0), //o
    .port_o_3_1 (sbox_AES_BoyarPeralta_28_port_o_3_1), //o
    .port_o_3_2 (sbox_AES_BoyarPeralta_28_port_o_3_2), //o
    .port_o_3_3 (sbox_AES_BoyarPeralta_28_port_o_3_3), //o
    .port_o_3_4 (sbox_AES_BoyarPeralta_28_port_o_3_4), //o
    .port_o_3_5 (sbox_AES_BoyarPeralta_28_port_o_3_5), //o
    .port_o_3_6 (sbox_AES_BoyarPeralta_28_port_o_3_6), //o
    .port_o_3_7 (sbox_AES_BoyarPeralta_28_port_o_3_7), //o
    .clk        (clk                                ), //i
    .reset      (reset                              )  //i
  );
  Sbox_AES_BoyarPeralta sbox_AES_BoyarPeralta_29 (
    .port_i_0_0 (keyAdd_port_state_out_13_0_0       ), //i
    .port_i_0_1 (keyAdd_port_state_out_13_0_1       ), //i
    .port_i_0_2 (keyAdd_port_state_out_13_0_2       ), //i
    .port_i_0_3 (keyAdd_port_state_out_13_0_3       ), //i
    .port_i_0_4 (keyAdd_port_state_out_13_0_4       ), //i
    .port_i_0_5 (keyAdd_port_state_out_13_0_5       ), //i
    .port_i_0_6 (keyAdd_port_state_out_13_0_6       ), //i
    .port_i_0_7 (keyAdd_port_state_out_13_0_7       ), //i
    .port_i_1_0 (keyAdd_port_state_out_13_1_0       ), //i
    .port_i_1_1 (keyAdd_port_state_out_13_1_1       ), //i
    .port_i_1_2 (keyAdd_port_state_out_13_1_2       ), //i
    .port_i_1_3 (keyAdd_port_state_out_13_1_3       ), //i
    .port_i_1_4 (keyAdd_port_state_out_13_1_4       ), //i
    .port_i_1_5 (keyAdd_port_state_out_13_1_5       ), //i
    .port_i_1_6 (keyAdd_port_state_out_13_1_6       ), //i
    .port_i_1_7 (keyAdd_port_state_out_13_1_7       ), //i
    .port_i_2_0 (keyAdd_port_state_out_13_2_0       ), //i
    .port_i_2_1 (keyAdd_port_state_out_13_2_1       ), //i
    .port_i_2_2 (keyAdd_port_state_out_13_2_2       ), //i
    .port_i_2_3 (keyAdd_port_state_out_13_2_3       ), //i
    .port_i_2_4 (keyAdd_port_state_out_13_2_4       ), //i
    .port_i_2_5 (keyAdd_port_state_out_13_2_5       ), //i
    .port_i_2_6 (keyAdd_port_state_out_13_2_6       ), //i
    .port_i_2_7 (keyAdd_port_state_out_13_2_7       ), //i
    .port_i_3_0 (keyAdd_port_state_out_13_3_0       ), //i
    .port_i_3_1 (keyAdd_port_state_out_13_3_1       ), //i
    .port_i_3_2 (keyAdd_port_state_out_13_3_2       ), //i
    .port_i_3_3 (keyAdd_port_state_out_13_3_3       ), //i
    .port_i_3_4 (keyAdd_port_state_out_13_3_4       ), //i
    .port_i_3_5 (keyAdd_port_state_out_13_3_5       ), //i
    .port_i_3_6 (keyAdd_port_state_out_13_3_6       ), //i
    .port_i_3_7 (keyAdd_port_state_out_13_3_7       ), //i
    .port_o_0_0 (sbox_AES_BoyarPeralta_29_port_o_0_0), //o
    .port_o_0_1 (sbox_AES_BoyarPeralta_29_port_o_0_1), //o
    .port_o_0_2 (sbox_AES_BoyarPeralta_29_port_o_0_2), //o
    .port_o_0_3 (sbox_AES_BoyarPeralta_29_port_o_0_3), //o
    .port_o_0_4 (sbox_AES_BoyarPeralta_29_port_o_0_4), //o
    .port_o_0_5 (sbox_AES_BoyarPeralta_29_port_o_0_5), //o
    .port_o_0_6 (sbox_AES_BoyarPeralta_29_port_o_0_6), //o
    .port_o_0_7 (sbox_AES_BoyarPeralta_29_port_o_0_7), //o
    .port_o_1_0 (sbox_AES_BoyarPeralta_29_port_o_1_0), //o
    .port_o_1_1 (sbox_AES_BoyarPeralta_29_port_o_1_1), //o
    .port_o_1_2 (sbox_AES_BoyarPeralta_29_port_o_1_2), //o
    .port_o_1_3 (sbox_AES_BoyarPeralta_29_port_o_1_3), //o
    .port_o_1_4 (sbox_AES_BoyarPeralta_29_port_o_1_4), //o
    .port_o_1_5 (sbox_AES_BoyarPeralta_29_port_o_1_5), //o
    .port_o_1_6 (sbox_AES_BoyarPeralta_29_port_o_1_6), //o
    .port_o_1_7 (sbox_AES_BoyarPeralta_29_port_o_1_7), //o
    .port_o_2_0 (sbox_AES_BoyarPeralta_29_port_o_2_0), //o
    .port_o_2_1 (sbox_AES_BoyarPeralta_29_port_o_2_1), //o
    .port_o_2_2 (sbox_AES_BoyarPeralta_29_port_o_2_2), //o
    .port_o_2_3 (sbox_AES_BoyarPeralta_29_port_o_2_3), //o
    .port_o_2_4 (sbox_AES_BoyarPeralta_29_port_o_2_4), //o
    .port_o_2_5 (sbox_AES_BoyarPeralta_29_port_o_2_5), //o
    .port_o_2_6 (sbox_AES_BoyarPeralta_29_port_o_2_6), //o
    .port_o_2_7 (sbox_AES_BoyarPeralta_29_port_o_2_7), //o
    .port_o_3_0 (sbox_AES_BoyarPeralta_29_port_o_3_0), //o
    .port_o_3_1 (sbox_AES_BoyarPeralta_29_port_o_3_1), //o
    .port_o_3_2 (sbox_AES_BoyarPeralta_29_port_o_3_2), //o
    .port_o_3_3 (sbox_AES_BoyarPeralta_29_port_o_3_3), //o
    .port_o_3_4 (sbox_AES_BoyarPeralta_29_port_o_3_4), //o
    .port_o_3_5 (sbox_AES_BoyarPeralta_29_port_o_3_5), //o
    .port_o_3_6 (sbox_AES_BoyarPeralta_29_port_o_3_6), //o
    .port_o_3_7 (sbox_AES_BoyarPeralta_29_port_o_3_7), //o
    .clk        (clk                                ), //i
    .reset      (reset                              )  //i
  );
  Sbox_AES_BoyarPeralta sbox_AES_BoyarPeralta_30 (
    .port_i_0_0 (keyAdd_port_state_out_14_0_0       ), //i
    .port_i_0_1 (keyAdd_port_state_out_14_0_1       ), //i
    .port_i_0_2 (keyAdd_port_state_out_14_0_2       ), //i
    .port_i_0_3 (keyAdd_port_state_out_14_0_3       ), //i
    .port_i_0_4 (keyAdd_port_state_out_14_0_4       ), //i
    .port_i_0_5 (keyAdd_port_state_out_14_0_5       ), //i
    .port_i_0_6 (keyAdd_port_state_out_14_0_6       ), //i
    .port_i_0_7 (keyAdd_port_state_out_14_0_7       ), //i
    .port_i_1_0 (keyAdd_port_state_out_14_1_0       ), //i
    .port_i_1_1 (keyAdd_port_state_out_14_1_1       ), //i
    .port_i_1_2 (keyAdd_port_state_out_14_1_2       ), //i
    .port_i_1_3 (keyAdd_port_state_out_14_1_3       ), //i
    .port_i_1_4 (keyAdd_port_state_out_14_1_4       ), //i
    .port_i_1_5 (keyAdd_port_state_out_14_1_5       ), //i
    .port_i_1_6 (keyAdd_port_state_out_14_1_6       ), //i
    .port_i_1_7 (keyAdd_port_state_out_14_1_7       ), //i
    .port_i_2_0 (keyAdd_port_state_out_14_2_0       ), //i
    .port_i_2_1 (keyAdd_port_state_out_14_2_1       ), //i
    .port_i_2_2 (keyAdd_port_state_out_14_2_2       ), //i
    .port_i_2_3 (keyAdd_port_state_out_14_2_3       ), //i
    .port_i_2_4 (keyAdd_port_state_out_14_2_4       ), //i
    .port_i_2_5 (keyAdd_port_state_out_14_2_5       ), //i
    .port_i_2_6 (keyAdd_port_state_out_14_2_6       ), //i
    .port_i_2_7 (keyAdd_port_state_out_14_2_7       ), //i
    .port_i_3_0 (keyAdd_port_state_out_14_3_0       ), //i
    .port_i_3_1 (keyAdd_port_state_out_14_3_1       ), //i
    .port_i_3_2 (keyAdd_port_state_out_14_3_2       ), //i
    .port_i_3_3 (keyAdd_port_state_out_14_3_3       ), //i
    .port_i_3_4 (keyAdd_port_state_out_14_3_4       ), //i
    .port_i_3_5 (keyAdd_port_state_out_14_3_5       ), //i
    .port_i_3_6 (keyAdd_port_state_out_14_3_6       ), //i
    .port_i_3_7 (keyAdd_port_state_out_14_3_7       ), //i
    .port_o_0_0 (sbox_AES_BoyarPeralta_30_port_o_0_0), //o
    .port_o_0_1 (sbox_AES_BoyarPeralta_30_port_o_0_1), //o
    .port_o_0_2 (sbox_AES_BoyarPeralta_30_port_o_0_2), //o
    .port_o_0_3 (sbox_AES_BoyarPeralta_30_port_o_0_3), //o
    .port_o_0_4 (sbox_AES_BoyarPeralta_30_port_o_0_4), //o
    .port_o_0_5 (sbox_AES_BoyarPeralta_30_port_o_0_5), //o
    .port_o_0_6 (sbox_AES_BoyarPeralta_30_port_o_0_6), //o
    .port_o_0_7 (sbox_AES_BoyarPeralta_30_port_o_0_7), //o
    .port_o_1_0 (sbox_AES_BoyarPeralta_30_port_o_1_0), //o
    .port_o_1_1 (sbox_AES_BoyarPeralta_30_port_o_1_1), //o
    .port_o_1_2 (sbox_AES_BoyarPeralta_30_port_o_1_2), //o
    .port_o_1_3 (sbox_AES_BoyarPeralta_30_port_o_1_3), //o
    .port_o_1_4 (sbox_AES_BoyarPeralta_30_port_o_1_4), //o
    .port_o_1_5 (sbox_AES_BoyarPeralta_30_port_o_1_5), //o
    .port_o_1_6 (sbox_AES_BoyarPeralta_30_port_o_1_6), //o
    .port_o_1_7 (sbox_AES_BoyarPeralta_30_port_o_1_7), //o
    .port_o_2_0 (sbox_AES_BoyarPeralta_30_port_o_2_0), //o
    .port_o_2_1 (sbox_AES_BoyarPeralta_30_port_o_2_1), //o
    .port_o_2_2 (sbox_AES_BoyarPeralta_30_port_o_2_2), //o
    .port_o_2_3 (sbox_AES_BoyarPeralta_30_port_o_2_3), //o
    .port_o_2_4 (sbox_AES_BoyarPeralta_30_port_o_2_4), //o
    .port_o_2_5 (sbox_AES_BoyarPeralta_30_port_o_2_5), //o
    .port_o_2_6 (sbox_AES_BoyarPeralta_30_port_o_2_6), //o
    .port_o_2_7 (sbox_AES_BoyarPeralta_30_port_o_2_7), //o
    .port_o_3_0 (sbox_AES_BoyarPeralta_30_port_o_3_0), //o
    .port_o_3_1 (sbox_AES_BoyarPeralta_30_port_o_3_1), //o
    .port_o_3_2 (sbox_AES_BoyarPeralta_30_port_o_3_2), //o
    .port_o_3_3 (sbox_AES_BoyarPeralta_30_port_o_3_3), //o
    .port_o_3_4 (sbox_AES_BoyarPeralta_30_port_o_3_4), //o
    .port_o_3_5 (sbox_AES_BoyarPeralta_30_port_o_3_5), //o
    .port_o_3_6 (sbox_AES_BoyarPeralta_30_port_o_3_6), //o
    .port_o_3_7 (sbox_AES_BoyarPeralta_30_port_o_3_7), //o
    .clk        (clk                                ), //i
    .reset      (reset                              )  //i
  );
  Sbox_AES_BoyarPeralta sbox_AES_BoyarPeralta_31 (
    .port_i_0_0 (keyAdd_port_state_out_15_0_0       ), //i
    .port_i_0_1 (keyAdd_port_state_out_15_0_1       ), //i
    .port_i_0_2 (keyAdd_port_state_out_15_0_2       ), //i
    .port_i_0_3 (keyAdd_port_state_out_15_0_3       ), //i
    .port_i_0_4 (keyAdd_port_state_out_15_0_4       ), //i
    .port_i_0_5 (keyAdd_port_state_out_15_0_5       ), //i
    .port_i_0_6 (keyAdd_port_state_out_15_0_6       ), //i
    .port_i_0_7 (keyAdd_port_state_out_15_0_7       ), //i
    .port_i_1_0 (keyAdd_port_state_out_15_1_0       ), //i
    .port_i_1_1 (keyAdd_port_state_out_15_1_1       ), //i
    .port_i_1_2 (keyAdd_port_state_out_15_1_2       ), //i
    .port_i_1_3 (keyAdd_port_state_out_15_1_3       ), //i
    .port_i_1_4 (keyAdd_port_state_out_15_1_4       ), //i
    .port_i_1_5 (keyAdd_port_state_out_15_1_5       ), //i
    .port_i_1_6 (keyAdd_port_state_out_15_1_6       ), //i
    .port_i_1_7 (keyAdd_port_state_out_15_1_7       ), //i
    .port_i_2_0 (keyAdd_port_state_out_15_2_0       ), //i
    .port_i_2_1 (keyAdd_port_state_out_15_2_1       ), //i
    .port_i_2_2 (keyAdd_port_state_out_15_2_2       ), //i
    .port_i_2_3 (keyAdd_port_state_out_15_2_3       ), //i
    .port_i_2_4 (keyAdd_port_state_out_15_2_4       ), //i
    .port_i_2_5 (keyAdd_port_state_out_15_2_5       ), //i
    .port_i_2_6 (keyAdd_port_state_out_15_2_6       ), //i
    .port_i_2_7 (keyAdd_port_state_out_15_2_7       ), //i
    .port_i_3_0 (keyAdd_port_state_out_15_3_0       ), //i
    .port_i_3_1 (keyAdd_port_state_out_15_3_1       ), //i
    .port_i_3_2 (keyAdd_port_state_out_15_3_2       ), //i
    .port_i_3_3 (keyAdd_port_state_out_15_3_3       ), //i
    .port_i_3_4 (keyAdd_port_state_out_15_3_4       ), //i
    .port_i_3_5 (keyAdd_port_state_out_15_3_5       ), //i
    .port_i_3_6 (keyAdd_port_state_out_15_3_6       ), //i
    .port_i_3_7 (keyAdd_port_state_out_15_3_7       ), //i
    .port_o_0_0 (sbox_AES_BoyarPeralta_31_port_o_0_0), //o
    .port_o_0_1 (sbox_AES_BoyarPeralta_31_port_o_0_1), //o
    .port_o_0_2 (sbox_AES_BoyarPeralta_31_port_o_0_2), //o
    .port_o_0_3 (sbox_AES_BoyarPeralta_31_port_o_0_3), //o
    .port_o_0_4 (sbox_AES_BoyarPeralta_31_port_o_0_4), //o
    .port_o_0_5 (sbox_AES_BoyarPeralta_31_port_o_0_5), //o
    .port_o_0_6 (sbox_AES_BoyarPeralta_31_port_o_0_6), //o
    .port_o_0_7 (sbox_AES_BoyarPeralta_31_port_o_0_7), //o
    .port_o_1_0 (sbox_AES_BoyarPeralta_31_port_o_1_0), //o
    .port_o_1_1 (sbox_AES_BoyarPeralta_31_port_o_1_1), //o
    .port_o_1_2 (sbox_AES_BoyarPeralta_31_port_o_1_2), //o
    .port_o_1_3 (sbox_AES_BoyarPeralta_31_port_o_1_3), //o
    .port_o_1_4 (sbox_AES_BoyarPeralta_31_port_o_1_4), //o
    .port_o_1_5 (sbox_AES_BoyarPeralta_31_port_o_1_5), //o
    .port_o_1_6 (sbox_AES_BoyarPeralta_31_port_o_1_6), //o
    .port_o_1_7 (sbox_AES_BoyarPeralta_31_port_o_1_7), //o
    .port_o_2_0 (sbox_AES_BoyarPeralta_31_port_o_2_0), //o
    .port_o_2_1 (sbox_AES_BoyarPeralta_31_port_o_2_1), //o
    .port_o_2_2 (sbox_AES_BoyarPeralta_31_port_o_2_2), //o
    .port_o_2_3 (sbox_AES_BoyarPeralta_31_port_o_2_3), //o
    .port_o_2_4 (sbox_AES_BoyarPeralta_31_port_o_2_4), //o
    .port_o_2_5 (sbox_AES_BoyarPeralta_31_port_o_2_5), //o
    .port_o_2_6 (sbox_AES_BoyarPeralta_31_port_o_2_6), //o
    .port_o_2_7 (sbox_AES_BoyarPeralta_31_port_o_2_7), //o
    .port_o_3_0 (sbox_AES_BoyarPeralta_31_port_o_3_0), //o
    .port_o_3_1 (sbox_AES_BoyarPeralta_31_port_o_3_1), //o
    .port_o_3_2 (sbox_AES_BoyarPeralta_31_port_o_3_2), //o
    .port_o_3_3 (sbox_AES_BoyarPeralta_31_port_o_3_3), //o
    .port_o_3_4 (sbox_AES_BoyarPeralta_31_port_o_3_4), //o
    .port_o_3_5 (sbox_AES_BoyarPeralta_31_port_o_3_5), //o
    .port_o_3_6 (sbox_AES_BoyarPeralta_31_port_o_3_6), //o
    .port_o_3_7 (sbox_AES_BoyarPeralta_31_port_o_3_7), //o
    .clk        (clk                                ), //i
    .reset      (reset                              )  //i
  );
  AES_ShiftRows shiftRows (
    .port_state_in_0_0_0   (subBytes_out_0_0_0             ), //i
    .port_state_in_0_0_1   (subBytes_out_0_0_1             ), //i
    .port_state_in_0_0_2   (subBytes_out_0_0_2             ), //i
    .port_state_in_0_0_3   (subBytes_out_0_0_3             ), //i
    .port_state_in_0_0_4   (subBytes_out_0_0_4             ), //i
    .port_state_in_0_0_5   (subBytes_out_0_0_5             ), //i
    .port_state_in_0_0_6   (subBytes_out_0_0_6             ), //i
    .port_state_in_0_0_7   (subBytes_out_0_0_7             ), //i
    .port_state_in_0_1_0   (subBytes_out_0_1_0             ), //i
    .port_state_in_0_1_1   (subBytes_out_0_1_1             ), //i
    .port_state_in_0_1_2   (subBytes_out_0_1_2             ), //i
    .port_state_in_0_1_3   (subBytes_out_0_1_3             ), //i
    .port_state_in_0_1_4   (subBytes_out_0_1_4             ), //i
    .port_state_in_0_1_5   (subBytes_out_0_1_5             ), //i
    .port_state_in_0_1_6   (subBytes_out_0_1_6             ), //i
    .port_state_in_0_1_7   (subBytes_out_0_1_7             ), //i
    .port_state_in_0_2_0   (subBytes_out_0_2_0             ), //i
    .port_state_in_0_2_1   (subBytes_out_0_2_1             ), //i
    .port_state_in_0_2_2   (subBytes_out_0_2_2             ), //i
    .port_state_in_0_2_3   (subBytes_out_0_2_3             ), //i
    .port_state_in_0_2_4   (subBytes_out_0_2_4             ), //i
    .port_state_in_0_2_5   (subBytes_out_0_2_5             ), //i
    .port_state_in_0_2_6   (subBytes_out_0_2_6             ), //i
    .port_state_in_0_2_7   (subBytes_out_0_2_7             ), //i
    .port_state_in_0_3_0   (subBytes_out_0_3_0             ), //i
    .port_state_in_0_3_1   (subBytes_out_0_3_1             ), //i
    .port_state_in_0_3_2   (subBytes_out_0_3_2             ), //i
    .port_state_in_0_3_3   (subBytes_out_0_3_3             ), //i
    .port_state_in_0_3_4   (subBytes_out_0_3_4             ), //i
    .port_state_in_0_3_5   (subBytes_out_0_3_5             ), //i
    .port_state_in_0_3_6   (subBytes_out_0_3_6             ), //i
    .port_state_in_0_3_7   (subBytes_out_0_3_7             ), //i
    .port_state_in_1_0_0   (subBytes_out_1_0_0             ), //i
    .port_state_in_1_0_1   (subBytes_out_1_0_1             ), //i
    .port_state_in_1_0_2   (subBytes_out_1_0_2             ), //i
    .port_state_in_1_0_3   (subBytes_out_1_0_3             ), //i
    .port_state_in_1_0_4   (subBytes_out_1_0_4             ), //i
    .port_state_in_1_0_5   (subBytes_out_1_0_5             ), //i
    .port_state_in_1_0_6   (subBytes_out_1_0_6             ), //i
    .port_state_in_1_0_7   (subBytes_out_1_0_7             ), //i
    .port_state_in_1_1_0   (subBytes_out_1_1_0             ), //i
    .port_state_in_1_1_1   (subBytes_out_1_1_1             ), //i
    .port_state_in_1_1_2   (subBytes_out_1_1_2             ), //i
    .port_state_in_1_1_3   (subBytes_out_1_1_3             ), //i
    .port_state_in_1_1_4   (subBytes_out_1_1_4             ), //i
    .port_state_in_1_1_5   (subBytes_out_1_1_5             ), //i
    .port_state_in_1_1_6   (subBytes_out_1_1_6             ), //i
    .port_state_in_1_1_7   (subBytes_out_1_1_7             ), //i
    .port_state_in_1_2_0   (subBytes_out_1_2_0             ), //i
    .port_state_in_1_2_1   (subBytes_out_1_2_1             ), //i
    .port_state_in_1_2_2   (subBytes_out_1_2_2             ), //i
    .port_state_in_1_2_3   (subBytes_out_1_2_3             ), //i
    .port_state_in_1_2_4   (subBytes_out_1_2_4             ), //i
    .port_state_in_1_2_5   (subBytes_out_1_2_5             ), //i
    .port_state_in_1_2_6   (subBytes_out_1_2_6             ), //i
    .port_state_in_1_2_7   (subBytes_out_1_2_7             ), //i
    .port_state_in_1_3_0   (subBytes_out_1_3_0             ), //i
    .port_state_in_1_3_1   (subBytes_out_1_3_1             ), //i
    .port_state_in_1_3_2   (subBytes_out_1_3_2             ), //i
    .port_state_in_1_3_3   (subBytes_out_1_3_3             ), //i
    .port_state_in_1_3_4   (subBytes_out_1_3_4             ), //i
    .port_state_in_1_3_5   (subBytes_out_1_3_5             ), //i
    .port_state_in_1_3_6   (subBytes_out_1_3_6             ), //i
    .port_state_in_1_3_7   (subBytes_out_1_3_7             ), //i
    .port_state_in_2_0_0   (subBytes_out_2_0_0             ), //i
    .port_state_in_2_0_1   (subBytes_out_2_0_1             ), //i
    .port_state_in_2_0_2   (subBytes_out_2_0_2             ), //i
    .port_state_in_2_0_3   (subBytes_out_2_0_3             ), //i
    .port_state_in_2_0_4   (subBytes_out_2_0_4             ), //i
    .port_state_in_2_0_5   (subBytes_out_2_0_5             ), //i
    .port_state_in_2_0_6   (subBytes_out_2_0_6             ), //i
    .port_state_in_2_0_7   (subBytes_out_2_0_7             ), //i
    .port_state_in_2_1_0   (subBytes_out_2_1_0             ), //i
    .port_state_in_2_1_1   (subBytes_out_2_1_1             ), //i
    .port_state_in_2_1_2   (subBytes_out_2_1_2             ), //i
    .port_state_in_2_1_3   (subBytes_out_2_1_3             ), //i
    .port_state_in_2_1_4   (subBytes_out_2_1_4             ), //i
    .port_state_in_2_1_5   (subBytes_out_2_1_5             ), //i
    .port_state_in_2_1_6   (subBytes_out_2_1_6             ), //i
    .port_state_in_2_1_7   (subBytes_out_2_1_7             ), //i
    .port_state_in_2_2_0   (subBytes_out_2_2_0             ), //i
    .port_state_in_2_2_1   (subBytes_out_2_2_1             ), //i
    .port_state_in_2_2_2   (subBytes_out_2_2_2             ), //i
    .port_state_in_2_2_3   (subBytes_out_2_2_3             ), //i
    .port_state_in_2_2_4   (subBytes_out_2_2_4             ), //i
    .port_state_in_2_2_5   (subBytes_out_2_2_5             ), //i
    .port_state_in_2_2_6   (subBytes_out_2_2_6             ), //i
    .port_state_in_2_2_7   (subBytes_out_2_2_7             ), //i
    .port_state_in_2_3_0   (subBytes_out_2_3_0             ), //i
    .port_state_in_2_3_1   (subBytes_out_2_3_1             ), //i
    .port_state_in_2_3_2   (subBytes_out_2_3_2             ), //i
    .port_state_in_2_3_3   (subBytes_out_2_3_3             ), //i
    .port_state_in_2_3_4   (subBytes_out_2_3_4             ), //i
    .port_state_in_2_3_5   (subBytes_out_2_3_5             ), //i
    .port_state_in_2_3_6   (subBytes_out_2_3_6             ), //i
    .port_state_in_2_3_7   (subBytes_out_2_3_7             ), //i
    .port_state_in_3_0_0   (subBytes_out_3_0_0             ), //i
    .port_state_in_3_0_1   (subBytes_out_3_0_1             ), //i
    .port_state_in_3_0_2   (subBytes_out_3_0_2             ), //i
    .port_state_in_3_0_3   (subBytes_out_3_0_3             ), //i
    .port_state_in_3_0_4   (subBytes_out_3_0_4             ), //i
    .port_state_in_3_0_5   (subBytes_out_3_0_5             ), //i
    .port_state_in_3_0_6   (subBytes_out_3_0_6             ), //i
    .port_state_in_3_0_7   (subBytes_out_3_0_7             ), //i
    .port_state_in_3_1_0   (subBytes_out_3_1_0             ), //i
    .port_state_in_3_1_1   (subBytes_out_3_1_1             ), //i
    .port_state_in_3_1_2   (subBytes_out_3_1_2             ), //i
    .port_state_in_3_1_3   (subBytes_out_3_1_3             ), //i
    .port_state_in_3_1_4   (subBytes_out_3_1_4             ), //i
    .port_state_in_3_1_5   (subBytes_out_3_1_5             ), //i
    .port_state_in_3_1_6   (subBytes_out_3_1_6             ), //i
    .port_state_in_3_1_7   (subBytes_out_3_1_7             ), //i
    .port_state_in_3_2_0   (subBytes_out_3_2_0             ), //i
    .port_state_in_3_2_1   (subBytes_out_3_2_1             ), //i
    .port_state_in_3_2_2   (subBytes_out_3_2_2             ), //i
    .port_state_in_3_2_3   (subBytes_out_3_2_3             ), //i
    .port_state_in_3_2_4   (subBytes_out_3_2_4             ), //i
    .port_state_in_3_2_5   (subBytes_out_3_2_5             ), //i
    .port_state_in_3_2_6   (subBytes_out_3_2_6             ), //i
    .port_state_in_3_2_7   (subBytes_out_3_2_7             ), //i
    .port_state_in_3_3_0   (subBytes_out_3_3_0             ), //i
    .port_state_in_3_3_1   (subBytes_out_3_3_1             ), //i
    .port_state_in_3_3_2   (subBytes_out_3_3_2             ), //i
    .port_state_in_3_3_3   (subBytes_out_3_3_3             ), //i
    .port_state_in_3_3_4   (subBytes_out_3_3_4             ), //i
    .port_state_in_3_3_5   (subBytes_out_3_3_5             ), //i
    .port_state_in_3_3_6   (subBytes_out_3_3_6             ), //i
    .port_state_in_3_3_7   (subBytes_out_3_3_7             ), //i
    .port_state_in_4_0_0   (subBytes_out_4_0_0             ), //i
    .port_state_in_4_0_1   (subBytes_out_4_0_1             ), //i
    .port_state_in_4_0_2   (subBytes_out_4_0_2             ), //i
    .port_state_in_4_0_3   (subBytes_out_4_0_3             ), //i
    .port_state_in_4_0_4   (subBytes_out_4_0_4             ), //i
    .port_state_in_4_0_5   (subBytes_out_4_0_5             ), //i
    .port_state_in_4_0_6   (subBytes_out_4_0_6             ), //i
    .port_state_in_4_0_7   (subBytes_out_4_0_7             ), //i
    .port_state_in_4_1_0   (subBytes_out_4_1_0             ), //i
    .port_state_in_4_1_1   (subBytes_out_4_1_1             ), //i
    .port_state_in_4_1_2   (subBytes_out_4_1_2             ), //i
    .port_state_in_4_1_3   (subBytes_out_4_1_3             ), //i
    .port_state_in_4_1_4   (subBytes_out_4_1_4             ), //i
    .port_state_in_4_1_5   (subBytes_out_4_1_5             ), //i
    .port_state_in_4_1_6   (subBytes_out_4_1_6             ), //i
    .port_state_in_4_1_7   (subBytes_out_4_1_7             ), //i
    .port_state_in_4_2_0   (subBytes_out_4_2_0             ), //i
    .port_state_in_4_2_1   (subBytes_out_4_2_1             ), //i
    .port_state_in_4_2_2   (subBytes_out_4_2_2             ), //i
    .port_state_in_4_2_3   (subBytes_out_4_2_3             ), //i
    .port_state_in_4_2_4   (subBytes_out_4_2_4             ), //i
    .port_state_in_4_2_5   (subBytes_out_4_2_5             ), //i
    .port_state_in_4_2_6   (subBytes_out_4_2_6             ), //i
    .port_state_in_4_2_7   (subBytes_out_4_2_7             ), //i
    .port_state_in_4_3_0   (subBytes_out_4_3_0             ), //i
    .port_state_in_4_3_1   (subBytes_out_4_3_1             ), //i
    .port_state_in_4_3_2   (subBytes_out_4_3_2             ), //i
    .port_state_in_4_3_3   (subBytes_out_4_3_3             ), //i
    .port_state_in_4_3_4   (subBytes_out_4_3_4             ), //i
    .port_state_in_4_3_5   (subBytes_out_4_3_5             ), //i
    .port_state_in_4_3_6   (subBytes_out_4_3_6             ), //i
    .port_state_in_4_3_7   (subBytes_out_4_3_7             ), //i
    .port_state_in_5_0_0   (subBytes_out_5_0_0             ), //i
    .port_state_in_5_0_1   (subBytes_out_5_0_1             ), //i
    .port_state_in_5_0_2   (subBytes_out_5_0_2             ), //i
    .port_state_in_5_0_3   (subBytes_out_5_0_3             ), //i
    .port_state_in_5_0_4   (subBytes_out_5_0_4             ), //i
    .port_state_in_5_0_5   (subBytes_out_5_0_5             ), //i
    .port_state_in_5_0_6   (subBytes_out_5_0_6             ), //i
    .port_state_in_5_0_7   (subBytes_out_5_0_7             ), //i
    .port_state_in_5_1_0   (subBytes_out_5_1_0             ), //i
    .port_state_in_5_1_1   (subBytes_out_5_1_1             ), //i
    .port_state_in_5_1_2   (subBytes_out_5_1_2             ), //i
    .port_state_in_5_1_3   (subBytes_out_5_1_3             ), //i
    .port_state_in_5_1_4   (subBytes_out_5_1_4             ), //i
    .port_state_in_5_1_5   (subBytes_out_5_1_5             ), //i
    .port_state_in_5_1_6   (subBytes_out_5_1_6             ), //i
    .port_state_in_5_1_7   (subBytes_out_5_1_7             ), //i
    .port_state_in_5_2_0   (subBytes_out_5_2_0             ), //i
    .port_state_in_5_2_1   (subBytes_out_5_2_1             ), //i
    .port_state_in_5_2_2   (subBytes_out_5_2_2             ), //i
    .port_state_in_5_2_3   (subBytes_out_5_2_3             ), //i
    .port_state_in_5_2_4   (subBytes_out_5_2_4             ), //i
    .port_state_in_5_2_5   (subBytes_out_5_2_5             ), //i
    .port_state_in_5_2_6   (subBytes_out_5_2_6             ), //i
    .port_state_in_5_2_7   (subBytes_out_5_2_7             ), //i
    .port_state_in_5_3_0   (subBytes_out_5_3_0             ), //i
    .port_state_in_5_3_1   (subBytes_out_5_3_1             ), //i
    .port_state_in_5_3_2   (subBytes_out_5_3_2             ), //i
    .port_state_in_5_3_3   (subBytes_out_5_3_3             ), //i
    .port_state_in_5_3_4   (subBytes_out_5_3_4             ), //i
    .port_state_in_5_3_5   (subBytes_out_5_3_5             ), //i
    .port_state_in_5_3_6   (subBytes_out_5_3_6             ), //i
    .port_state_in_5_3_7   (subBytes_out_5_3_7             ), //i
    .port_state_in_6_0_0   (subBytes_out_6_0_0             ), //i
    .port_state_in_6_0_1   (subBytes_out_6_0_1             ), //i
    .port_state_in_6_0_2   (subBytes_out_6_0_2             ), //i
    .port_state_in_6_0_3   (subBytes_out_6_0_3             ), //i
    .port_state_in_6_0_4   (subBytes_out_6_0_4             ), //i
    .port_state_in_6_0_5   (subBytes_out_6_0_5             ), //i
    .port_state_in_6_0_6   (subBytes_out_6_0_6             ), //i
    .port_state_in_6_0_7   (subBytes_out_6_0_7             ), //i
    .port_state_in_6_1_0   (subBytes_out_6_1_0             ), //i
    .port_state_in_6_1_1   (subBytes_out_6_1_1             ), //i
    .port_state_in_6_1_2   (subBytes_out_6_1_2             ), //i
    .port_state_in_6_1_3   (subBytes_out_6_1_3             ), //i
    .port_state_in_6_1_4   (subBytes_out_6_1_4             ), //i
    .port_state_in_6_1_5   (subBytes_out_6_1_5             ), //i
    .port_state_in_6_1_6   (subBytes_out_6_1_6             ), //i
    .port_state_in_6_1_7   (subBytes_out_6_1_7             ), //i
    .port_state_in_6_2_0   (subBytes_out_6_2_0             ), //i
    .port_state_in_6_2_1   (subBytes_out_6_2_1             ), //i
    .port_state_in_6_2_2   (subBytes_out_6_2_2             ), //i
    .port_state_in_6_2_3   (subBytes_out_6_2_3             ), //i
    .port_state_in_6_2_4   (subBytes_out_6_2_4             ), //i
    .port_state_in_6_2_5   (subBytes_out_6_2_5             ), //i
    .port_state_in_6_2_6   (subBytes_out_6_2_6             ), //i
    .port_state_in_6_2_7   (subBytes_out_6_2_7             ), //i
    .port_state_in_6_3_0   (subBytes_out_6_3_0             ), //i
    .port_state_in_6_3_1   (subBytes_out_6_3_1             ), //i
    .port_state_in_6_3_2   (subBytes_out_6_3_2             ), //i
    .port_state_in_6_3_3   (subBytes_out_6_3_3             ), //i
    .port_state_in_6_3_4   (subBytes_out_6_3_4             ), //i
    .port_state_in_6_3_5   (subBytes_out_6_3_5             ), //i
    .port_state_in_6_3_6   (subBytes_out_6_3_6             ), //i
    .port_state_in_6_3_7   (subBytes_out_6_3_7             ), //i
    .port_state_in_7_0_0   (subBytes_out_7_0_0             ), //i
    .port_state_in_7_0_1   (subBytes_out_7_0_1             ), //i
    .port_state_in_7_0_2   (subBytes_out_7_0_2             ), //i
    .port_state_in_7_0_3   (subBytes_out_7_0_3             ), //i
    .port_state_in_7_0_4   (subBytes_out_7_0_4             ), //i
    .port_state_in_7_0_5   (subBytes_out_7_0_5             ), //i
    .port_state_in_7_0_6   (subBytes_out_7_0_6             ), //i
    .port_state_in_7_0_7   (subBytes_out_7_0_7             ), //i
    .port_state_in_7_1_0   (subBytes_out_7_1_0             ), //i
    .port_state_in_7_1_1   (subBytes_out_7_1_1             ), //i
    .port_state_in_7_1_2   (subBytes_out_7_1_2             ), //i
    .port_state_in_7_1_3   (subBytes_out_7_1_3             ), //i
    .port_state_in_7_1_4   (subBytes_out_7_1_4             ), //i
    .port_state_in_7_1_5   (subBytes_out_7_1_5             ), //i
    .port_state_in_7_1_6   (subBytes_out_7_1_6             ), //i
    .port_state_in_7_1_7   (subBytes_out_7_1_7             ), //i
    .port_state_in_7_2_0   (subBytes_out_7_2_0             ), //i
    .port_state_in_7_2_1   (subBytes_out_7_2_1             ), //i
    .port_state_in_7_2_2   (subBytes_out_7_2_2             ), //i
    .port_state_in_7_2_3   (subBytes_out_7_2_3             ), //i
    .port_state_in_7_2_4   (subBytes_out_7_2_4             ), //i
    .port_state_in_7_2_5   (subBytes_out_7_2_5             ), //i
    .port_state_in_7_2_6   (subBytes_out_7_2_6             ), //i
    .port_state_in_7_2_7   (subBytes_out_7_2_7             ), //i
    .port_state_in_7_3_0   (subBytes_out_7_3_0             ), //i
    .port_state_in_7_3_1   (subBytes_out_7_3_1             ), //i
    .port_state_in_7_3_2   (subBytes_out_7_3_2             ), //i
    .port_state_in_7_3_3   (subBytes_out_7_3_3             ), //i
    .port_state_in_7_3_4   (subBytes_out_7_3_4             ), //i
    .port_state_in_7_3_5   (subBytes_out_7_3_5             ), //i
    .port_state_in_7_3_6   (subBytes_out_7_3_6             ), //i
    .port_state_in_7_3_7   (subBytes_out_7_3_7             ), //i
    .port_state_in_8_0_0   (subBytes_out_8_0_0             ), //i
    .port_state_in_8_0_1   (subBytes_out_8_0_1             ), //i
    .port_state_in_8_0_2   (subBytes_out_8_0_2             ), //i
    .port_state_in_8_0_3   (subBytes_out_8_0_3             ), //i
    .port_state_in_8_0_4   (subBytes_out_8_0_4             ), //i
    .port_state_in_8_0_5   (subBytes_out_8_0_5             ), //i
    .port_state_in_8_0_6   (subBytes_out_8_0_6             ), //i
    .port_state_in_8_0_7   (subBytes_out_8_0_7             ), //i
    .port_state_in_8_1_0   (subBytes_out_8_1_0             ), //i
    .port_state_in_8_1_1   (subBytes_out_8_1_1             ), //i
    .port_state_in_8_1_2   (subBytes_out_8_1_2             ), //i
    .port_state_in_8_1_3   (subBytes_out_8_1_3             ), //i
    .port_state_in_8_1_4   (subBytes_out_8_1_4             ), //i
    .port_state_in_8_1_5   (subBytes_out_8_1_5             ), //i
    .port_state_in_8_1_6   (subBytes_out_8_1_6             ), //i
    .port_state_in_8_1_7   (subBytes_out_8_1_7             ), //i
    .port_state_in_8_2_0   (subBytes_out_8_2_0             ), //i
    .port_state_in_8_2_1   (subBytes_out_8_2_1             ), //i
    .port_state_in_8_2_2   (subBytes_out_8_2_2             ), //i
    .port_state_in_8_2_3   (subBytes_out_8_2_3             ), //i
    .port_state_in_8_2_4   (subBytes_out_8_2_4             ), //i
    .port_state_in_8_2_5   (subBytes_out_8_2_5             ), //i
    .port_state_in_8_2_6   (subBytes_out_8_2_6             ), //i
    .port_state_in_8_2_7   (subBytes_out_8_2_7             ), //i
    .port_state_in_8_3_0   (subBytes_out_8_3_0             ), //i
    .port_state_in_8_3_1   (subBytes_out_8_3_1             ), //i
    .port_state_in_8_3_2   (subBytes_out_8_3_2             ), //i
    .port_state_in_8_3_3   (subBytes_out_8_3_3             ), //i
    .port_state_in_8_3_4   (subBytes_out_8_3_4             ), //i
    .port_state_in_8_3_5   (subBytes_out_8_3_5             ), //i
    .port_state_in_8_3_6   (subBytes_out_8_3_6             ), //i
    .port_state_in_8_3_7   (subBytes_out_8_3_7             ), //i
    .port_state_in_9_0_0   (subBytes_out_9_0_0             ), //i
    .port_state_in_9_0_1   (subBytes_out_9_0_1             ), //i
    .port_state_in_9_0_2   (subBytes_out_9_0_2             ), //i
    .port_state_in_9_0_3   (subBytes_out_9_0_3             ), //i
    .port_state_in_9_0_4   (subBytes_out_9_0_4             ), //i
    .port_state_in_9_0_5   (subBytes_out_9_0_5             ), //i
    .port_state_in_9_0_6   (subBytes_out_9_0_6             ), //i
    .port_state_in_9_0_7   (subBytes_out_9_0_7             ), //i
    .port_state_in_9_1_0   (subBytes_out_9_1_0             ), //i
    .port_state_in_9_1_1   (subBytes_out_9_1_1             ), //i
    .port_state_in_9_1_2   (subBytes_out_9_1_2             ), //i
    .port_state_in_9_1_3   (subBytes_out_9_1_3             ), //i
    .port_state_in_9_1_4   (subBytes_out_9_1_4             ), //i
    .port_state_in_9_1_5   (subBytes_out_9_1_5             ), //i
    .port_state_in_9_1_6   (subBytes_out_9_1_6             ), //i
    .port_state_in_9_1_7   (subBytes_out_9_1_7             ), //i
    .port_state_in_9_2_0   (subBytes_out_9_2_0             ), //i
    .port_state_in_9_2_1   (subBytes_out_9_2_1             ), //i
    .port_state_in_9_2_2   (subBytes_out_9_2_2             ), //i
    .port_state_in_9_2_3   (subBytes_out_9_2_3             ), //i
    .port_state_in_9_2_4   (subBytes_out_9_2_4             ), //i
    .port_state_in_9_2_5   (subBytes_out_9_2_5             ), //i
    .port_state_in_9_2_6   (subBytes_out_9_2_6             ), //i
    .port_state_in_9_2_7   (subBytes_out_9_2_7             ), //i
    .port_state_in_9_3_0   (subBytes_out_9_3_0             ), //i
    .port_state_in_9_3_1   (subBytes_out_9_3_1             ), //i
    .port_state_in_9_3_2   (subBytes_out_9_3_2             ), //i
    .port_state_in_9_3_3   (subBytes_out_9_3_3             ), //i
    .port_state_in_9_3_4   (subBytes_out_9_3_4             ), //i
    .port_state_in_9_3_5   (subBytes_out_9_3_5             ), //i
    .port_state_in_9_3_6   (subBytes_out_9_3_6             ), //i
    .port_state_in_9_3_7   (subBytes_out_9_3_7             ), //i
    .port_state_in_10_0_0  (subBytes_out_10_0_0            ), //i
    .port_state_in_10_0_1  (subBytes_out_10_0_1            ), //i
    .port_state_in_10_0_2  (subBytes_out_10_0_2            ), //i
    .port_state_in_10_0_3  (subBytes_out_10_0_3            ), //i
    .port_state_in_10_0_4  (subBytes_out_10_0_4            ), //i
    .port_state_in_10_0_5  (subBytes_out_10_0_5            ), //i
    .port_state_in_10_0_6  (subBytes_out_10_0_6            ), //i
    .port_state_in_10_0_7  (subBytes_out_10_0_7            ), //i
    .port_state_in_10_1_0  (subBytes_out_10_1_0            ), //i
    .port_state_in_10_1_1  (subBytes_out_10_1_1            ), //i
    .port_state_in_10_1_2  (subBytes_out_10_1_2            ), //i
    .port_state_in_10_1_3  (subBytes_out_10_1_3            ), //i
    .port_state_in_10_1_4  (subBytes_out_10_1_4            ), //i
    .port_state_in_10_1_5  (subBytes_out_10_1_5            ), //i
    .port_state_in_10_1_6  (subBytes_out_10_1_6            ), //i
    .port_state_in_10_1_7  (subBytes_out_10_1_7            ), //i
    .port_state_in_10_2_0  (subBytes_out_10_2_0            ), //i
    .port_state_in_10_2_1  (subBytes_out_10_2_1            ), //i
    .port_state_in_10_2_2  (subBytes_out_10_2_2            ), //i
    .port_state_in_10_2_3  (subBytes_out_10_2_3            ), //i
    .port_state_in_10_2_4  (subBytes_out_10_2_4            ), //i
    .port_state_in_10_2_5  (subBytes_out_10_2_5            ), //i
    .port_state_in_10_2_6  (subBytes_out_10_2_6            ), //i
    .port_state_in_10_2_7  (subBytes_out_10_2_7            ), //i
    .port_state_in_10_3_0  (subBytes_out_10_3_0            ), //i
    .port_state_in_10_3_1  (subBytes_out_10_3_1            ), //i
    .port_state_in_10_3_2  (subBytes_out_10_3_2            ), //i
    .port_state_in_10_3_3  (subBytes_out_10_3_3            ), //i
    .port_state_in_10_3_4  (subBytes_out_10_3_4            ), //i
    .port_state_in_10_3_5  (subBytes_out_10_3_5            ), //i
    .port_state_in_10_3_6  (subBytes_out_10_3_6            ), //i
    .port_state_in_10_3_7  (subBytes_out_10_3_7            ), //i
    .port_state_in_11_0_0  (subBytes_out_11_0_0            ), //i
    .port_state_in_11_0_1  (subBytes_out_11_0_1            ), //i
    .port_state_in_11_0_2  (subBytes_out_11_0_2            ), //i
    .port_state_in_11_0_3  (subBytes_out_11_0_3            ), //i
    .port_state_in_11_0_4  (subBytes_out_11_0_4            ), //i
    .port_state_in_11_0_5  (subBytes_out_11_0_5            ), //i
    .port_state_in_11_0_6  (subBytes_out_11_0_6            ), //i
    .port_state_in_11_0_7  (subBytes_out_11_0_7            ), //i
    .port_state_in_11_1_0  (subBytes_out_11_1_0            ), //i
    .port_state_in_11_1_1  (subBytes_out_11_1_1            ), //i
    .port_state_in_11_1_2  (subBytes_out_11_1_2            ), //i
    .port_state_in_11_1_3  (subBytes_out_11_1_3            ), //i
    .port_state_in_11_1_4  (subBytes_out_11_1_4            ), //i
    .port_state_in_11_1_5  (subBytes_out_11_1_5            ), //i
    .port_state_in_11_1_6  (subBytes_out_11_1_6            ), //i
    .port_state_in_11_1_7  (subBytes_out_11_1_7            ), //i
    .port_state_in_11_2_0  (subBytes_out_11_2_0            ), //i
    .port_state_in_11_2_1  (subBytes_out_11_2_1            ), //i
    .port_state_in_11_2_2  (subBytes_out_11_2_2            ), //i
    .port_state_in_11_2_3  (subBytes_out_11_2_3            ), //i
    .port_state_in_11_2_4  (subBytes_out_11_2_4            ), //i
    .port_state_in_11_2_5  (subBytes_out_11_2_5            ), //i
    .port_state_in_11_2_6  (subBytes_out_11_2_6            ), //i
    .port_state_in_11_2_7  (subBytes_out_11_2_7            ), //i
    .port_state_in_11_3_0  (subBytes_out_11_3_0            ), //i
    .port_state_in_11_3_1  (subBytes_out_11_3_1            ), //i
    .port_state_in_11_3_2  (subBytes_out_11_3_2            ), //i
    .port_state_in_11_3_3  (subBytes_out_11_3_3            ), //i
    .port_state_in_11_3_4  (subBytes_out_11_3_4            ), //i
    .port_state_in_11_3_5  (subBytes_out_11_3_5            ), //i
    .port_state_in_11_3_6  (subBytes_out_11_3_6            ), //i
    .port_state_in_11_3_7  (subBytes_out_11_3_7            ), //i
    .port_state_in_12_0_0  (subBytes_out_12_0_0            ), //i
    .port_state_in_12_0_1  (subBytes_out_12_0_1            ), //i
    .port_state_in_12_0_2  (subBytes_out_12_0_2            ), //i
    .port_state_in_12_0_3  (subBytes_out_12_0_3            ), //i
    .port_state_in_12_0_4  (subBytes_out_12_0_4            ), //i
    .port_state_in_12_0_5  (subBytes_out_12_0_5            ), //i
    .port_state_in_12_0_6  (subBytes_out_12_0_6            ), //i
    .port_state_in_12_0_7  (subBytes_out_12_0_7            ), //i
    .port_state_in_12_1_0  (subBytes_out_12_1_0            ), //i
    .port_state_in_12_1_1  (subBytes_out_12_1_1            ), //i
    .port_state_in_12_1_2  (subBytes_out_12_1_2            ), //i
    .port_state_in_12_1_3  (subBytes_out_12_1_3            ), //i
    .port_state_in_12_1_4  (subBytes_out_12_1_4            ), //i
    .port_state_in_12_1_5  (subBytes_out_12_1_5            ), //i
    .port_state_in_12_1_6  (subBytes_out_12_1_6            ), //i
    .port_state_in_12_1_7  (subBytes_out_12_1_7            ), //i
    .port_state_in_12_2_0  (subBytes_out_12_2_0            ), //i
    .port_state_in_12_2_1  (subBytes_out_12_2_1            ), //i
    .port_state_in_12_2_2  (subBytes_out_12_2_2            ), //i
    .port_state_in_12_2_3  (subBytes_out_12_2_3            ), //i
    .port_state_in_12_2_4  (subBytes_out_12_2_4            ), //i
    .port_state_in_12_2_5  (subBytes_out_12_2_5            ), //i
    .port_state_in_12_2_6  (subBytes_out_12_2_6            ), //i
    .port_state_in_12_2_7  (subBytes_out_12_2_7            ), //i
    .port_state_in_12_3_0  (subBytes_out_12_3_0            ), //i
    .port_state_in_12_3_1  (subBytes_out_12_3_1            ), //i
    .port_state_in_12_3_2  (subBytes_out_12_3_2            ), //i
    .port_state_in_12_3_3  (subBytes_out_12_3_3            ), //i
    .port_state_in_12_3_4  (subBytes_out_12_3_4            ), //i
    .port_state_in_12_3_5  (subBytes_out_12_3_5            ), //i
    .port_state_in_12_3_6  (subBytes_out_12_3_6            ), //i
    .port_state_in_12_3_7  (subBytes_out_12_3_7            ), //i
    .port_state_in_13_0_0  (subBytes_out_13_0_0            ), //i
    .port_state_in_13_0_1  (subBytes_out_13_0_1            ), //i
    .port_state_in_13_0_2  (subBytes_out_13_0_2            ), //i
    .port_state_in_13_0_3  (subBytes_out_13_0_3            ), //i
    .port_state_in_13_0_4  (subBytes_out_13_0_4            ), //i
    .port_state_in_13_0_5  (subBytes_out_13_0_5            ), //i
    .port_state_in_13_0_6  (subBytes_out_13_0_6            ), //i
    .port_state_in_13_0_7  (subBytes_out_13_0_7            ), //i
    .port_state_in_13_1_0  (subBytes_out_13_1_0            ), //i
    .port_state_in_13_1_1  (subBytes_out_13_1_1            ), //i
    .port_state_in_13_1_2  (subBytes_out_13_1_2            ), //i
    .port_state_in_13_1_3  (subBytes_out_13_1_3            ), //i
    .port_state_in_13_1_4  (subBytes_out_13_1_4            ), //i
    .port_state_in_13_1_5  (subBytes_out_13_1_5            ), //i
    .port_state_in_13_1_6  (subBytes_out_13_1_6            ), //i
    .port_state_in_13_1_7  (subBytes_out_13_1_7            ), //i
    .port_state_in_13_2_0  (subBytes_out_13_2_0            ), //i
    .port_state_in_13_2_1  (subBytes_out_13_2_1            ), //i
    .port_state_in_13_2_2  (subBytes_out_13_2_2            ), //i
    .port_state_in_13_2_3  (subBytes_out_13_2_3            ), //i
    .port_state_in_13_2_4  (subBytes_out_13_2_4            ), //i
    .port_state_in_13_2_5  (subBytes_out_13_2_5            ), //i
    .port_state_in_13_2_6  (subBytes_out_13_2_6            ), //i
    .port_state_in_13_2_7  (subBytes_out_13_2_7            ), //i
    .port_state_in_13_3_0  (subBytes_out_13_3_0            ), //i
    .port_state_in_13_3_1  (subBytes_out_13_3_1            ), //i
    .port_state_in_13_3_2  (subBytes_out_13_3_2            ), //i
    .port_state_in_13_3_3  (subBytes_out_13_3_3            ), //i
    .port_state_in_13_3_4  (subBytes_out_13_3_4            ), //i
    .port_state_in_13_3_5  (subBytes_out_13_3_5            ), //i
    .port_state_in_13_3_6  (subBytes_out_13_3_6            ), //i
    .port_state_in_13_3_7  (subBytes_out_13_3_7            ), //i
    .port_state_in_14_0_0  (subBytes_out_14_0_0            ), //i
    .port_state_in_14_0_1  (subBytes_out_14_0_1            ), //i
    .port_state_in_14_0_2  (subBytes_out_14_0_2            ), //i
    .port_state_in_14_0_3  (subBytes_out_14_0_3            ), //i
    .port_state_in_14_0_4  (subBytes_out_14_0_4            ), //i
    .port_state_in_14_0_5  (subBytes_out_14_0_5            ), //i
    .port_state_in_14_0_6  (subBytes_out_14_0_6            ), //i
    .port_state_in_14_0_7  (subBytes_out_14_0_7            ), //i
    .port_state_in_14_1_0  (subBytes_out_14_1_0            ), //i
    .port_state_in_14_1_1  (subBytes_out_14_1_1            ), //i
    .port_state_in_14_1_2  (subBytes_out_14_1_2            ), //i
    .port_state_in_14_1_3  (subBytes_out_14_1_3            ), //i
    .port_state_in_14_1_4  (subBytes_out_14_1_4            ), //i
    .port_state_in_14_1_5  (subBytes_out_14_1_5            ), //i
    .port_state_in_14_1_6  (subBytes_out_14_1_6            ), //i
    .port_state_in_14_1_7  (subBytes_out_14_1_7            ), //i
    .port_state_in_14_2_0  (subBytes_out_14_2_0            ), //i
    .port_state_in_14_2_1  (subBytes_out_14_2_1            ), //i
    .port_state_in_14_2_2  (subBytes_out_14_2_2            ), //i
    .port_state_in_14_2_3  (subBytes_out_14_2_3            ), //i
    .port_state_in_14_2_4  (subBytes_out_14_2_4            ), //i
    .port_state_in_14_2_5  (subBytes_out_14_2_5            ), //i
    .port_state_in_14_2_6  (subBytes_out_14_2_6            ), //i
    .port_state_in_14_2_7  (subBytes_out_14_2_7            ), //i
    .port_state_in_14_3_0  (subBytes_out_14_3_0            ), //i
    .port_state_in_14_3_1  (subBytes_out_14_3_1            ), //i
    .port_state_in_14_3_2  (subBytes_out_14_3_2            ), //i
    .port_state_in_14_3_3  (subBytes_out_14_3_3            ), //i
    .port_state_in_14_3_4  (subBytes_out_14_3_4            ), //i
    .port_state_in_14_3_5  (subBytes_out_14_3_5            ), //i
    .port_state_in_14_3_6  (subBytes_out_14_3_6            ), //i
    .port_state_in_14_3_7  (subBytes_out_14_3_7            ), //i
    .port_state_in_15_0_0  (subBytes_out_15_0_0            ), //i
    .port_state_in_15_0_1  (subBytes_out_15_0_1            ), //i
    .port_state_in_15_0_2  (subBytes_out_15_0_2            ), //i
    .port_state_in_15_0_3  (subBytes_out_15_0_3            ), //i
    .port_state_in_15_0_4  (subBytes_out_15_0_4            ), //i
    .port_state_in_15_0_5  (subBytes_out_15_0_5            ), //i
    .port_state_in_15_0_6  (subBytes_out_15_0_6            ), //i
    .port_state_in_15_0_7  (subBytes_out_15_0_7            ), //i
    .port_state_in_15_1_0  (subBytes_out_15_1_0            ), //i
    .port_state_in_15_1_1  (subBytes_out_15_1_1            ), //i
    .port_state_in_15_1_2  (subBytes_out_15_1_2            ), //i
    .port_state_in_15_1_3  (subBytes_out_15_1_3            ), //i
    .port_state_in_15_1_4  (subBytes_out_15_1_4            ), //i
    .port_state_in_15_1_5  (subBytes_out_15_1_5            ), //i
    .port_state_in_15_1_6  (subBytes_out_15_1_6            ), //i
    .port_state_in_15_1_7  (subBytes_out_15_1_7            ), //i
    .port_state_in_15_2_0  (subBytes_out_15_2_0            ), //i
    .port_state_in_15_2_1  (subBytes_out_15_2_1            ), //i
    .port_state_in_15_2_2  (subBytes_out_15_2_2            ), //i
    .port_state_in_15_2_3  (subBytes_out_15_2_3            ), //i
    .port_state_in_15_2_4  (subBytes_out_15_2_4            ), //i
    .port_state_in_15_2_5  (subBytes_out_15_2_5            ), //i
    .port_state_in_15_2_6  (subBytes_out_15_2_6            ), //i
    .port_state_in_15_2_7  (subBytes_out_15_2_7            ), //i
    .port_state_in_15_3_0  (subBytes_out_15_3_0            ), //i
    .port_state_in_15_3_1  (subBytes_out_15_3_1            ), //i
    .port_state_in_15_3_2  (subBytes_out_15_3_2            ), //i
    .port_state_in_15_3_3  (subBytes_out_15_3_3            ), //i
    .port_state_in_15_3_4  (subBytes_out_15_3_4            ), //i
    .port_state_in_15_3_5  (subBytes_out_15_3_5            ), //i
    .port_state_in_15_3_6  (subBytes_out_15_3_6            ), //i
    .port_state_in_15_3_7  (subBytes_out_15_3_7            ), //i
    .port_state_out_0_0_0  (shiftRows_port_state_out_0_0_0 ), //o
    .port_state_out_0_0_1  (shiftRows_port_state_out_0_0_1 ), //o
    .port_state_out_0_0_2  (shiftRows_port_state_out_0_0_2 ), //o
    .port_state_out_0_0_3  (shiftRows_port_state_out_0_0_3 ), //o
    .port_state_out_0_0_4  (shiftRows_port_state_out_0_0_4 ), //o
    .port_state_out_0_0_5  (shiftRows_port_state_out_0_0_5 ), //o
    .port_state_out_0_0_6  (shiftRows_port_state_out_0_0_6 ), //o
    .port_state_out_0_0_7  (shiftRows_port_state_out_0_0_7 ), //o
    .port_state_out_0_1_0  (shiftRows_port_state_out_0_1_0 ), //o
    .port_state_out_0_1_1  (shiftRows_port_state_out_0_1_1 ), //o
    .port_state_out_0_1_2  (shiftRows_port_state_out_0_1_2 ), //o
    .port_state_out_0_1_3  (shiftRows_port_state_out_0_1_3 ), //o
    .port_state_out_0_1_4  (shiftRows_port_state_out_0_1_4 ), //o
    .port_state_out_0_1_5  (shiftRows_port_state_out_0_1_5 ), //o
    .port_state_out_0_1_6  (shiftRows_port_state_out_0_1_6 ), //o
    .port_state_out_0_1_7  (shiftRows_port_state_out_0_1_7 ), //o
    .port_state_out_0_2_0  (shiftRows_port_state_out_0_2_0 ), //o
    .port_state_out_0_2_1  (shiftRows_port_state_out_0_2_1 ), //o
    .port_state_out_0_2_2  (shiftRows_port_state_out_0_2_2 ), //o
    .port_state_out_0_2_3  (shiftRows_port_state_out_0_2_3 ), //o
    .port_state_out_0_2_4  (shiftRows_port_state_out_0_2_4 ), //o
    .port_state_out_0_2_5  (shiftRows_port_state_out_0_2_5 ), //o
    .port_state_out_0_2_6  (shiftRows_port_state_out_0_2_6 ), //o
    .port_state_out_0_2_7  (shiftRows_port_state_out_0_2_7 ), //o
    .port_state_out_0_3_0  (shiftRows_port_state_out_0_3_0 ), //o
    .port_state_out_0_3_1  (shiftRows_port_state_out_0_3_1 ), //o
    .port_state_out_0_3_2  (shiftRows_port_state_out_0_3_2 ), //o
    .port_state_out_0_3_3  (shiftRows_port_state_out_0_3_3 ), //o
    .port_state_out_0_3_4  (shiftRows_port_state_out_0_3_4 ), //o
    .port_state_out_0_3_5  (shiftRows_port_state_out_0_3_5 ), //o
    .port_state_out_0_3_6  (shiftRows_port_state_out_0_3_6 ), //o
    .port_state_out_0_3_7  (shiftRows_port_state_out_0_3_7 ), //o
    .port_state_out_1_0_0  (shiftRows_port_state_out_1_0_0 ), //o
    .port_state_out_1_0_1  (shiftRows_port_state_out_1_0_1 ), //o
    .port_state_out_1_0_2  (shiftRows_port_state_out_1_0_2 ), //o
    .port_state_out_1_0_3  (shiftRows_port_state_out_1_0_3 ), //o
    .port_state_out_1_0_4  (shiftRows_port_state_out_1_0_4 ), //o
    .port_state_out_1_0_5  (shiftRows_port_state_out_1_0_5 ), //o
    .port_state_out_1_0_6  (shiftRows_port_state_out_1_0_6 ), //o
    .port_state_out_1_0_7  (shiftRows_port_state_out_1_0_7 ), //o
    .port_state_out_1_1_0  (shiftRows_port_state_out_1_1_0 ), //o
    .port_state_out_1_1_1  (shiftRows_port_state_out_1_1_1 ), //o
    .port_state_out_1_1_2  (shiftRows_port_state_out_1_1_2 ), //o
    .port_state_out_1_1_3  (shiftRows_port_state_out_1_1_3 ), //o
    .port_state_out_1_1_4  (shiftRows_port_state_out_1_1_4 ), //o
    .port_state_out_1_1_5  (shiftRows_port_state_out_1_1_5 ), //o
    .port_state_out_1_1_6  (shiftRows_port_state_out_1_1_6 ), //o
    .port_state_out_1_1_7  (shiftRows_port_state_out_1_1_7 ), //o
    .port_state_out_1_2_0  (shiftRows_port_state_out_1_2_0 ), //o
    .port_state_out_1_2_1  (shiftRows_port_state_out_1_2_1 ), //o
    .port_state_out_1_2_2  (shiftRows_port_state_out_1_2_2 ), //o
    .port_state_out_1_2_3  (shiftRows_port_state_out_1_2_3 ), //o
    .port_state_out_1_2_4  (shiftRows_port_state_out_1_2_4 ), //o
    .port_state_out_1_2_5  (shiftRows_port_state_out_1_2_5 ), //o
    .port_state_out_1_2_6  (shiftRows_port_state_out_1_2_6 ), //o
    .port_state_out_1_2_7  (shiftRows_port_state_out_1_2_7 ), //o
    .port_state_out_1_3_0  (shiftRows_port_state_out_1_3_0 ), //o
    .port_state_out_1_3_1  (shiftRows_port_state_out_1_3_1 ), //o
    .port_state_out_1_3_2  (shiftRows_port_state_out_1_3_2 ), //o
    .port_state_out_1_3_3  (shiftRows_port_state_out_1_3_3 ), //o
    .port_state_out_1_3_4  (shiftRows_port_state_out_1_3_4 ), //o
    .port_state_out_1_3_5  (shiftRows_port_state_out_1_3_5 ), //o
    .port_state_out_1_3_6  (shiftRows_port_state_out_1_3_6 ), //o
    .port_state_out_1_3_7  (shiftRows_port_state_out_1_3_7 ), //o
    .port_state_out_2_0_0  (shiftRows_port_state_out_2_0_0 ), //o
    .port_state_out_2_0_1  (shiftRows_port_state_out_2_0_1 ), //o
    .port_state_out_2_0_2  (shiftRows_port_state_out_2_0_2 ), //o
    .port_state_out_2_0_3  (shiftRows_port_state_out_2_0_3 ), //o
    .port_state_out_2_0_4  (shiftRows_port_state_out_2_0_4 ), //o
    .port_state_out_2_0_5  (shiftRows_port_state_out_2_0_5 ), //o
    .port_state_out_2_0_6  (shiftRows_port_state_out_2_0_6 ), //o
    .port_state_out_2_0_7  (shiftRows_port_state_out_2_0_7 ), //o
    .port_state_out_2_1_0  (shiftRows_port_state_out_2_1_0 ), //o
    .port_state_out_2_1_1  (shiftRows_port_state_out_2_1_1 ), //o
    .port_state_out_2_1_2  (shiftRows_port_state_out_2_1_2 ), //o
    .port_state_out_2_1_3  (shiftRows_port_state_out_2_1_3 ), //o
    .port_state_out_2_1_4  (shiftRows_port_state_out_2_1_4 ), //o
    .port_state_out_2_1_5  (shiftRows_port_state_out_2_1_5 ), //o
    .port_state_out_2_1_6  (shiftRows_port_state_out_2_1_6 ), //o
    .port_state_out_2_1_7  (shiftRows_port_state_out_2_1_7 ), //o
    .port_state_out_2_2_0  (shiftRows_port_state_out_2_2_0 ), //o
    .port_state_out_2_2_1  (shiftRows_port_state_out_2_2_1 ), //o
    .port_state_out_2_2_2  (shiftRows_port_state_out_2_2_2 ), //o
    .port_state_out_2_2_3  (shiftRows_port_state_out_2_2_3 ), //o
    .port_state_out_2_2_4  (shiftRows_port_state_out_2_2_4 ), //o
    .port_state_out_2_2_5  (shiftRows_port_state_out_2_2_5 ), //o
    .port_state_out_2_2_6  (shiftRows_port_state_out_2_2_6 ), //o
    .port_state_out_2_2_7  (shiftRows_port_state_out_2_2_7 ), //o
    .port_state_out_2_3_0  (shiftRows_port_state_out_2_3_0 ), //o
    .port_state_out_2_3_1  (shiftRows_port_state_out_2_3_1 ), //o
    .port_state_out_2_3_2  (shiftRows_port_state_out_2_3_2 ), //o
    .port_state_out_2_3_3  (shiftRows_port_state_out_2_3_3 ), //o
    .port_state_out_2_3_4  (shiftRows_port_state_out_2_3_4 ), //o
    .port_state_out_2_3_5  (shiftRows_port_state_out_2_3_5 ), //o
    .port_state_out_2_3_6  (shiftRows_port_state_out_2_3_6 ), //o
    .port_state_out_2_3_7  (shiftRows_port_state_out_2_3_7 ), //o
    .port_state_out_3_0_0  (shiftRows_port_state_out_3_0_0 ), //o
    .port_state_out_3_0_1  (shiftRows_port_state_out_3_0_1 ), //o
    .port_state_out_3_0_2  (shiftRows_port_state_out_3_0_2 ), //o
    .port_state_out_3_0_3  (shiftRows_port_state_out_3_0_3 ), //o
    .port_state_out_3_0_4  (shiftRows_port_state_out_3_0_4 ), //o
    .port_state_out_3_0_5  (shiftRows_port_state_out_3_0_5 ), //o
    .port_state_out_3_0_6  (shiftRows_port_state_out_3_0_6 ), //o
    .port_state_out_3_0_7  (shiftRows_port_state_out_3_0_7 ), //o
    .port_state_out_3_1_0  (shiftRows_port_state_out_3_1_0 ), //o
    .port_state_out_3_1_1  (shiftRows_port_state_out_3_1_1 ), //o
    .port_state_out_3_1_2  (shiftRows_port_state_out_3_1_2 ), //o
    .port_state_out_3_1_3  (shiftRows_port_state_out_3_1_3 ), //o
    .port_state_out_3_1_4  (shiftRows_port_state_out_3_1_4 ), //o
    .port_state_out_3_1_5  (shiftRows_port_state_out_3_1_5 ), //o
    .port_state_out_3_1_6  (shiftRows_port_state_out_3_1_6 ), //o
    .port_state_out_3_1_7  (shiftRows_port_state_out_3_1_7 ), //o
    .port_state_out_3_2_0  (shiftRows_port_state_out_3_2_0 ), //o
    .port_state_out_3_2_1  (shiftRows_port_state_out_3_2_1 ), //o
    .port_state_out_3_2_2  (shiftRows_port_state_out_3_2_2 ), //o
    .port_state_out_3_2_3  (shiftRows_port_state_out_3_2_3 ), //o
    .port_state_out_3_2_4  (shiftRows_port_state_out_3_2_4 ), //o
    .port_state_out_3_2_5  (shiftRows_port_state_out_3_2_5 ), //o
    .port_state_out_3_2_6  (shiftRows_port_state_out_3_2_6 ), //o
    .port_state_out_3_2_7  (shiftRows_port_state_out_3_2_7 ), //o
    .port_state_out_3_3_0  (shiftRows_port_state_out_3_3_0 ), //o
    .port_state_out_3_3_1  (shiftRows_port_state_out_3_3_1 ), //o
    .port_state_out_3_3_2  (shiftRows_port_state_out_3_3_2 ), //o
    .port_state_out_3_3_3  (shiftRows_port_state_out_3_3_3 ), //o
    .port_state_out_3_3_4  (shiftRows_port_state_out_3_3_4 ), //o
    .port_state_out_3_3_5  (shiftRows_port_state_out_3_3_5 ), //o
    .port_state_out_3_3_6  (shiftRows_port_state_out_3_3_6 ), //o
    .port_state_out_3_3_7  (shiftRows_port_state_out_3_3_7 ), //o
    .port_state_out_4_0_0  (shiftRows_port_state_out_4_0_0 ), //o
    .port_state_out_4_0_1  (shiftRows_port_state_out_4_0_1 ), //o
    .port_state_out_4_0_2  (shiftRows_port_state_out_4_0_2 ), //o
    .port_state_out_4_0_3  (shiftRows_port_state_out_4_0_3 ), //o
    .port_state_out_4_0_4  (shiftRows_port_state_out_4_0_4 ), //o
    .port_state_out_4_0_5  (shiftRows_port_state_out_4_0_5 ), //o
    .port_state_out_4_0_6  (shiftRows_port_state_out_4_0_6 ), //o
    .port_state_out_4_0_7  (shiftRows_port_state_out_4_0_7 ), //o
    .port_state_out_4_1_0  (shiftRows_port_state_out_4_1_0 ), //o
    .port_state_out_4_1_1  (shiftRows_port_state_out_4_1_1 ), //o
    .port_state_out_4_1_2  (shiftRows_port_state_out_4_1_2 ), //o
    .port_state_out_4_1_3  (shiftRows_port_state_out_4_1_3 ), //o
    .port_state_out_4_1_4  (shiftRows_port_state_out_4_1_4 ), //o
    .port_state_out_4_1_5  (shiftRows_port_state_out_4_1_5 ), //o
    .port_state_out_4_1_6  (shiftRows_port_state_out_4_1_6 ), //o
    .port_state_out_4_1_7  (shiftRows_port_state_out_4_1_7 ), //o
    .port_state_out_4_2_0  (shiftRows_port_state_out_4_2_0 ), //o
    .port_state_out_4_2_1  (shiftRows_port_state_out_4_2_1 ), //o
    .port_state_out_4_2_2  (shiftRows_port_state_out_4_2_2 ), //o
    .port_state_out_4_2_3  (shiftRows_port_state_out_4_2_3 ), //o
    .port_state_out_4_2_4  (shiftRows_port_state_out_4_2_4 ), //o
    .port_state_out_4_2_5  (shiftRows_port_state_out_4_2_5 ), //o
    .port_state_out_4_2_6  (shiftRows_port_state_out_4_2_6 ), //o
    .port_state_out_4_2_7  (shiftRows_port_state_out_4_2_7 ), //o
    .port_state_out_4_3_0  (shiftRows_port_state_out_4_3_0 ), //o
    .port_state_out_4_3_1  (shiftRows_port_state_out_4_3_1 ), //o
    .port_state_out_4_3_2  (shiftRows_port_state_out_4_3_2 ), //o
    .port_state_out_4_3_3  (shiftRows_port_state_out_4_3_3 ), //o
    .port_state_out_4_3_4  (shiftRows_port_state_out_4_3_4 ), //o
    .port_state_out_4_3_5  (shiftRows_port_state_out_4_3_5 ), //o
    .port_state_out_4_3_6  (shiftRows_port_state_out_4_3_6 ), //o
    .port_state_out_4_3_7  (shiftRows_port_state_out_4_3_7 ), //o
    .port_state_out_5_0_0  (shiftRows_port_state_out_5_0_0 ), //o
    .port_state_out_5_0_1  (shiftRows_port_state_out_5_0_1 ), //o
    .port_state_out_5_0_2  (shiftRows_port_state_out_5_0_2 ), //o
    .port_state_out_5_0_3  (shiftRows_port_state_out_5_0_3 ), //o
    .port_state_out_5_0_4  (shiftRows_port_state_out_5_0_4 ), //o
    .port_state_out_5_0_5  (shiftRows_port_state_out_5_0_5 ), //o
    .port_state_out_5_0_6  (shiftRows_port_state_out_5_0_6 ), //o
    .port_state_out_5_0_7  (shiftRows_port_state_out_5_0_7 ), //o
    .port_state_out_5_1_0  (shiftRows_port_state_out_5_1_0 ), //o
    .port_state_out_5_1_1  (shiftRows_port_state_out_5_1_1 ), //o
    .port_state_out_5_1_2  (shiftRows_port_state_out_5_1_2 ), //o
    .port_state_out_5_1_3  (shiftRows_port_state_out_5_1_3 ), //o
    .port_state_out_5_1_4  (shiftRows_port_state_out_5_1_4 ), //o
    .port_state_out_5_1_5  (shiftRows_port_state_out_5_1_5 ), //o
    .port_state_out_5_1_6  (shiftRows_port_state_out_5_1_6 ), //o
    .port_state_out_5_1_7  (shiftRows_port_state_out_5_1_7 ), //o
    .port_state_out_5_2_0  (shiftRows_port_state_out_5_2_0 ), //o
    .port_state_out_5_2_1  (shiftRows_port_state_out_5_2_1 ), //o
    .port_state_out_5_2_2  (shiftRows_port_state_out_5_2_2 ), //o
    .port_state_out_5_2_3  (shiftRows_port_state_out_5_2_3 ), //o
    .port_state_out_5_2_4  (shiftRows_port_state_out_5_2_4 ), //o
    .port_state_out_5_2_5  (shiftRows_port_state_out_5_2_5 ), //o
    .port_state_out_5_2_6  (shiftRows_port_state_out_5_2_6 ), //o
    .port_state_out_5_2_7  (shiftRows_port_state_out_5_2_7 ), //o
    .port_state_out_5_3_0  (shiftRows_port_state_out_5_3_0 ), //o
    .port_state_out_5_3_1  (shiftRows_port_state_out_5_3_1 ), //o
    .port_state_out_5_3_2  (shiftRows_port_state_out_5_3_2 ), //o
    .port_state_out_5_3_3  (shiftRows_port_state_out_5_3_3 ), //o
    .port_state_out_5_3_4  (shiftRows_port_state_out_5_3_4 ), //o
    .port_state_out_5_3_5  (shiftRows_port_state_out_5_3_5 ), //o
    .port_state_out_5_3_6  (shiftRows_port_state_out_5_3_6 ), //o
    .port_state_out_5_3_7  (shiftRows_port_state_out_5_3_7 ), //o
    .port_state_out_6_0_0  (shiftRows_port_state_out_6_0_0 ), //o
    .port_state_out_6_0_1  (shiftRows_port_state_out_6_0_1 ), //o
    .port_state_out_6_0_2  (shiftRows_port_state_out_6_0_2 ), //o
    .port_state_out_6_0_3  (shiftRows_port_state_out_6_0_3 ), //o
    .port_state_out_6_0_4  (shiftRows_port_state_out_6_0_4 ), //o
    .port_state_out_6_0_5  (shiftRows_port_state_out_6_0_5 ), //o
    .port_state_out_6_0_6  (shiftRows_port_state_out_6_0_6 ), //o
    .port_state_out_6_0_7  (shiftRows_port_state_out_6_0_7 ), //o
    .port_state_out_6_1_0  (shiftRows_port_state_out_6_1_0 ), //o
    .port_state_out_6_1_1  (shiftRows_port_state_out_6_1_1 ), //o
    .port_state_out_6_1_2  (shiftRows_port_state_out_6_1_2 ), //o
    .port_state_out_6_1_3  (shiftRows_port_state_out_6_1_3 ), //o
    .port_state_out_6_1_4  (shiftRows_port_state_out_6_1_4 ), //o
    .port_state_out_6_1_5  (shiftRows_port_state_out_6_1_5 ), //o
    .port_state_out_6_1_6  (shiftRows_port_state_out_6_1_6 ), //o
    .port_state_out_6_1_7  (shiftRows_port_state_out_6_1_7 ), //o
    .port_state_out_6_2_0  (shiftRows_port_state_out_6_2_0 ), //o
    .port_state_out_6_2_1  (shiftRows_port_state_out_6_2_1 ), //o
    .port_state_out_6_2_2  (shiftRows_port_state_out_6_2_2 ), //o
    .port_state_out_6_2_3  (shiftRows_port_state_out_6_2_3 ), //o
    .port_state_out_6_2_4  (shiftRows_port_state_out_6_2_4 ), //o
    .port_state_out_6_2_5  (shiftRows_port_state_out_6_2_5 ), //o
    .port_state_out_6_2_6  (shiftRows_port_state_out_6_2_6 ), //o
    .port_state_out_6_2_7  (shiftRows_port_state_out_6_2_7 ), //o
    .port_state_out_6_3_0  (shiftRows_port_state_out_6_3_0 ), //o
    .port_state_out_6_3_1  (shiftRows_port_state_out_6_3_1 ), //o
    .port_state_out_6_3_2  (shiftRows_port_state_out_6_3_2 ), //o
    .port_state_out_6_3_3  (shiftRows_port_state_out_6_3_3 ), //o
    .port_state_out_6_3_4  (shiftRows_port_state_out_6_3_4 ), //o
    .port_state_out_6_3_5  (shiftRows_port_state_out_6_3_5 ), //o
    .port_state_out_6_3_6  (shiftRows_port_state_out_6_3_6 ), //o
    .port_state_out_6_3_7  (shiftRows_port_state_out_6_3_7 ), //o
    .port_state_out_7_0_0  (shiftRows_port_state_out_7_0_0 ), //o
    .port_state_out_7_0_1  (shiftRows_port_state_out_7_0_1 ), //o
    .port_state_out_7_0_2  (shiftRows_port_state_out_7_0_2 ), //o
    .port_state_out_7_0_3  (shiftRows_port_state_out_7_0_3 ), //o
    .port_state_out_7_0_4  (shiftRows_port_state_out_7_0_4 ), //o
    .port_state_out_7_0_5  (shiftRows_port_state_out_7_0_5 ), //o
    .port_state_out_7_0_6  (shiftRows_port_state_out_7_0_6 ), //o
    .port_state_out_7_0_7  (shiftRows_port_state_out_7_0_7 ), //o
    .port_state_out_7_1_0  (shiftRows_port_state_out_7_1_0 ), //o
    .port_state_out_7_1_1  (shiftRows_port_state_out_7_1_1 ), //o
    .port_state_out_7_1_2  (shiftRows_port_state_out_7_1_2 ), //o
    .port_state_out_7_1_3  (shiftRows_port_state_out_7_1_3 ), //o
    .port_state_out_7_1_4  (shiftRows_port_state_out_7_1_4 ), //o
    .port_state_out_7_1_5  (shiftRows_port_state_out_7_1_5 ), //o
    .port_state_out_7_1_6  (shiftRows_port_state_out_7_1_6 ), //o
    .port_state_out_7_1_7  (shiftRows_port_state_out_7_1_7 ), //o
    .port_state_out_7_2_0  (shiftRows_port_state_out_7_2_0 ), //o
    .port_state_out_7_2_1  (shiftRows_port_state_out_7_2_1 ), //o
    .port_state_out_7_2_2  (shiftRows_port_state_out_7_2_2 ), //o
    .port_state_out_7_2_3  (shiftRows_port_state_out_7_2_3 ), //o
    .port_state_out_7_2_4  (shiftRows_port_state_out_7_2_4 ), //o
    .port_state_out_7_2_5  (shiftRows_port_state_out_7_2_5 ), //o
    .port_state_out_7_2_6  (shiftRows_port_state_out_7_2_6 ), //o
    .port_state_out_7_2_7  (shiftRows_port_state_out_7_2_7 ), //o
    .port_state_out_7_3_0  (shiftRows_port_state_out_7_3_0 ), //o
    .port_state_out_7_3_1  (shiftRows_port_state_out_7_3_1 ), //o
    .port_state_out_7_3_2  (shiftRows_port_state_out_7_3_2 ), //o
    .port_state_out_7_3_3  (shiftRows_port_state_out_7_3_3 ), //o
    .port_state_out_7_3_4  (shiftRows_port_state_out_7_3_4 ), //o
    .port_state_out_7_3_5  (shiftRows_port_state_out_7_3_5 ), //o
    .port_state_out_7_3_6  (shiftRows_port_state_out_7_3_6 ), //o
    .port_state_out_7_3_7  (shiftRows_port_state_out_7_3_7 ), //o
    .port_state_out_8_0_0  (shiftRows_port_state_out_8_0_0 ), //o
    .port_state_out_8_0_1  (shiftRows_port_state_out_8_0_1 ), //o
    .port_state_out_8_0_2  (shiftRows_port_state_out_8_0_2 ), //o
    .port_state_out_8_0_3  (shiftRows_port_state_out_8_0_3 ), //o
    .port_state_out_8_0_4  (shiftRows_port_state_out_8_0_4 ), //o
    .port_state_out_8_0_5  (shiftRows_port_state_out_8_0_5 ), //o
    .port_state_out_8_0_6  (shiftRows_port_state_out_8_0_6 ), //o
    .port_state_out_8_0_7  (shiftRows_port_state_out_8_0_7 ), //o
    .port_state_out_8_1_0  (shiftRows_port_state_out_8_1_0 ), //o
    .port_state_out_8_1_1  (shiftRows_port_state_out_8_1_1 ), //o
    .port_state_out_8_1_2  (shiftRows_port_state_out_8_1_2 ), //o
    .port_state_out_8_1_3  (shiftRows_port_state_out_8_1_3 ), //o
    .port_state_out_8_1_4  (shiftRows_port_state_out_8_1_4 ), //o
    .port_state_out_8_1_5  (shiftRows_port_state_out_8_1_5 ), //o
    .port_state_out_8_1_6  (shiftRows_port_state_out_8_1_6 ), //o
    .port_state_out_8_1_7  (shiftRows_port_state_out_8_1_7 ), //o
    .port_state_out_8_2_0  (shiftRows_port_state_out_8_2_0 ), //o
    .port_state_out_8_2_1  (shiftRows_port_state_out_8_2_1 ), //o
    .port_state_out_8_2_2  (shiftRows_port_state_out_8_2_2 ), //o
    .port_state_out_8_2_3  (shiftRows_port_state_out_8_2_3 ), //o
    .port_state_out_8_2_4  (shiftRows_port_state_out_8_2_4 ), //o
    .port_state_out_8_2_5  (shiftRows_port_state_out_8_2_5 ), //o
    .port_state_out_8_2_6  (shiftRows_port_state_out_8_2_6 ), //o
    .port_state_out_8_2_7  (shiftRows_port_state_out_8_2_7 ), //o
    .port_state_out_8_3_0  (shiftRows_port_state_out_8_3_0 ), //o
    .port_state_out_8_3_1  (shiftRows_port_state_out_8_3_1 ), //o
    .port_state_out_8_3_2  (shiftRows_port_state_out_8_3_2 ), //o
    .port_state_out_8_3_3  (shiftRows_port_state_out_8_3_3 ), //o
    .port_state_out_8_3_4  (shiftRows_port_state_out_8_3_4 ), //o
    .port_state_out_8_3_5  (shiftRows_port_state_out_8_3_5 ), //o
    .port_state_out_8_3_6  (shiftRows_port_state_out_8_3_6 ), //o
    .port_state_out_8_3_7  (shiftRows_port_state_out_8_3_7 ), //o
    .port_state_out_9_0_0  (shiftRows_port_state_out_9_0_0 ), //o
    .port_state_out_9_0_1  (shiftRows_port_state_out_9_0_1 ), //o
    .port_state_out_9_0_2  (shiftRows_port_state_out_9_0_2 ), //o
    .port_state_out_9_0_3  (shiftRows_port_state_out_9_0_3 ), //o
    .port_state_out_9_0_4  (shiftRows_port_state_out_9_0_4 ), //o
    .port_state_out_9_0_5  (shiftRows_port_state_out_9_0_5 ), //o
    .port_state_out_9_0_6  (shiftRows_port_state_out_9_0_6 ), //o
    .port_state_out_9_0_7  (shiftRows_port_state_out_9_0_7 ), //o
    .port_state_out_9_1_0  (shiftRows_port_state_out_9_1_0 ), //o
    .port_state_out_9_1_1  (shiftRows_port_state_out_9_1_1 ), //o
    .port_state_out_9_1_2  (shiftRows_port_state_out_9_1_2 ), //o
    .port_state_out_9_1_3  (shiftRows_port_state_out_9_1_3 ), //o
    .port_state_out_9_1_4  (shiftRows_port_state_out_9_1_4 ), //o
    .port_state_out_9_1_5  (shiftRows_port_state_out_9_1_5 ), //o
    .port_state_out_9_1_6  (shiftRows_port_state_out_9_1_6 ), //o
    .port_state_out_9_1_7  (shiftRows_port_state_out_9_1_7 ), //o
    .port_state_out_9_2_0  (shiftRows_port_state_out_9_2_0 ), //o
    .port_state_out_9_2_1  (shiftRows_port_state_out_9_2_1 ), //o
    .port_state_out_9_2_2  (shiftRows_port_state_out_9_2_2 ), //o
    .port_state_out_9_2_3  (shiftRows_port_state_out_9_2_3 ), //o
    .port_state_out_9_2_4  (shiftRows_port_state_out_9_2_4 ), //o
    .port_state_out_9_2_5  (shiftRows_port_state_out_9_2_5 ), //o
    .port_state_out_9_2_6  (shiftRows_port_state_out_9_2_6 ), //o
    .port_state_out_9_2_7  (shiftRows_port_state_out_9_2_7 ), //o
    .port_state_out_9_3_0  (shiftRows_port_state_out_9_3_0 ), //o
    .port_state_out_9_3_1  (shiftRows_port_state_out_9_3_1 ), //o
    .port_state_out_9_3_2  (shiftRows_port_state_out_9_3_2 ), //o
    .port_state_out_9_3_3  (shiftRows_port_state_out_9_3_3 ), //o
    .port_state_out_9_3_4  (shiftRows_port_state_out_9_3_4 ), //o
    .port_state_out_9_3_5  (shiftRows_port_state_out_9_3_5 ), //o
    .port_state_out_9_3_6  (shiftRows_port_state_out_9_3_6 ), //o
    .port_state_out_9_3_7  (shiftRows_port_state_out_9_3_7 ), //o
    .port_state_out_10_0_0 (shiftRows_port_state_out_10_0_0), //o
    .port_state_out_10_0_1 (shiftRows_port_state_out_10_0_1), //o
    .port_state_out_10_0_2 (shiftRows_port_state_out_10_0_2), //o
    .port_state_out_10_0_3 (shiftRows_port_state_out_10_0_3), //o
    .port_state_out_10_0_4 (shiftRows_port_state_out_10_0_4), //o
    .port_state_out_10_0_5 (shiftRows_port_state_out_10_0_5), //o
    .port_state_out_10_0_6 (shiftRows_port_state_out_10_0_6), //o
    .port_state_out_10_0_7 (shiftRows_port_state_out_10_0_7), //o
    .port_state_out_10_1_0 (shiftRows_port_state_out_10_1_0), //o
    .port_state_out_10_1_1 (shiftRows_port_state_out_10_1_1), //o
    .port_state_out_10_1_2 (shiftRows_port_state_out_10_1_2), //o
    .port_state_out_10_1_3 (shiftRows_port_state_out_10_1_3), //o
    .port_state_out_10_1_4 (shiftRows_port_state_out_10_1_4), //o
    .port_state_out_10_1_5 (shiftRows_port_state_out_10_1_5), //o
    .port_state_out_10_1_6 (shiftRows_port_state_out_10_1_6), //o
    .port_state_out_10_1_7 (shiftRows_port_state_out_10_1_7), //o
    .port_state_out_10_2_0 (shiftRows_port_state_out_10_2_0), //o
    .port_state_out_10_2_1 (shiftRows_port_state_out_10_2_1), //o
    .port_state_out_10_2_2 (shiftRows_port_state_out_10_2_2), //o
    .port_state_out_10_2_3 (shiftRows_port_state_out_10_2_3), //o
    .port_state_out_10_2_4 (shiftRows_port_state_out_10_2_4), //o
    .port_state_out_10_2_5 (shiftRows_port_state_out_10_2_5), //o
    .port_state_out_10_2_6 (shiftRows_port_state_out_10_2_6), //o
    .port_state_out_10_2_7 (shiftRows_port_state_out_10_2_7), //o
    .port_state_out_10_3_0 (shiftRows_port_state_out_10_3_0), //o
    .port_state_out_10_3_1 (shiftRows_port_state_out_10_3_1), //o
    .port_state_out_10_3_2 (shiftRows_port_state_out_10_3_2), //o
    .port_state_out_10_3_3 (shiftRows_port_state_out_10_3_3), //o
    .port_state_out_10_3_4 (shiftRows_port_state_out_10_3_4), //o
    .port_state_out_10_3_5 (shiftRows_port_state_out_10_3_5), //o
    .port_state_out_10_3_6 (shiftRows_port_state_out_10_3_6), //o
    .port_state_out_10_3_7 (shiftRows_port_state_out_10_3_7), //o
    .port_state_out_11_0_0 (shiftRows_port_state_out_11_0_0), //o
    .port_state_out_11_0_1 (shiftRows_port_state_out_11_0_1), //o
    .port_state_out_11_0_2 (shiftRows_port_state_out_11_0_2), //o
    .port_state_out_11_0_3 (shiftRows_port_state_out_11_0_3), //o
    .port_state_out_11_0_4 (shiftRows_port_state_out_11_0_4), //o
    .port_state_out_11_0_5 (shiftRows_port_state_out_11_0_5), //o
    .port_state_out_11_0_6 (shiftRows_port_state_out_11_0_6), //o
    .port_state_out_11_0_7 (shiftRows_port_state_out_11_0_7), //o
    .port_state_out_11_1_0 (shiftRows_port_state_out_11_1_0), //o
    .port_state_out_11_1_1 (shiftRows_port_state_out_11_1_1), //o
    .port_state_out_11_1_2 (shiftRows_port_state_out_11_1_2), //o
    .port_state_out_11_1_3 (shiftRows_port_state_out_11_1_3), //o
    .port_state_out_11_1_4 (shiftRows_port_state_out_11_1_4), //o
    .port_state_out_11_1_5 (shiftRows_port_state_out_11_1_5), //o
    .port_state_out_11_1_6 (shiftRows_port_state_out_11_1_6), //o
    .port_state_out_11_1_7 (shiftRows_port_state_out_11_1_7), //o
    .port_state_out_11_2_0 (shiftRows_port_state_out_11_2_0), //o
    .port_state_out_11_2_1 (shiftRows_port_state_out_11_2_1), //o
    .port_state_out_11_2_2 (shiftRows_port_state_out_11_2_2), //o
    .port_state_out_11_2_3 (shiftRows_port_state_out_11_2_3), //o
    .port_state_out_11_2_4 (shiftRows_port_state_out_11_2_4), //o
    .port_state_out_11_2_5 (shiftRows_port_state_out_11_2_5), //o
    .port_state_out_11_2_6 (shiftRows_port_state_out_11_2_6), //o
    .port_state_out_11_2_7 (shiftRows_port_state_out_11_2_7), //o
    .port_state_out_11_3_0 (shiftRows_port_state_out_11_3_0), //o
    .port_state_out_11_3_1 (shiftRows_port_state_out_11_3_1), //o
    .port_state_out_11_3_2 (shiftRows_port_state_out_11_3_2), //o
    .port_state_out_11_3_3 (shiftRows_port_state_out_11_3_3), //o
    .port_state_out_11_3_4 (shiftRows_port_state_out_11_3_4), //o
    .port_state_out_11_3_5 (shiftRows_port_state_out_11_3_5), //o
    .port_state_out_11_3_6 (shiftRows_port_state_out_11_3_6), //o
    .port_state_out_11_3_7 (shiftRows_port_state_out_11_3_7), //o
    .port_state_out_12_0_0 (shiftRows_port_state_out_12_0_0), //o
    .port_state_out_12_0_1 (shiftRows_port_state_out_12_0_1), //o
    .port_state_out_12_0_2 (shiftRows_port_state_out_12_0_2), //o
    .port_state_out_12_0_3 (shiftRows_port_state_out_12_0_3), //o
    .port_state_out_12_0_4 (shiftRows_port_state_out_12_0_4), //o
    .port_state_out_12_0_5 (shiftRows_port_state_out_12_0_5), //o
    .port_state_out_12_0_6 (shiftRows_port_state_out_12_0_6), //o
    .port_state_out_12_0_7 (shiftRows_port_state_out_12_0_7), //o
    .port_state_out_12_1_0 (shiftRows_port_state_out_12_1_0), //o
    .port_state_out_12_1_1 (shiftRows_port_state_out_12_1_1), //o
    .port_state_out_12_1_2 (shiftRows_port_state_out_12_1_2), //o
    .port_state_out_12_1_3 (shiftRows_port_state_out_12_1_3), //o
    .port_state_out_12_1_4 (shiftRows_port_state_out_12_1_4), //o
    .port_state_out_12_1_5 (shiftRows_port_state_out_12_1_5), //o
    .port_state_out_12_1_6 (shiftRows_port_state_out_12_1_6), //o
    .port_state_out_12_1_7 (shiftRows_port_state_out_12_1_7), //o
    .port_state_out_12_2_0 (shiftRows_port_state_out_12_2_0), //o
    .port_state_out_12_2_1 (shiftRows_port_state_out_12_2_1), //o
    .port_state_out_12_2_2 (shiftRows_port_state_out_12_2_2), //o
    .port_state_out_12_2_3 (shiftRows_port_state_out_12_2_3), //o
    .port_state_out_12_2_4 (shiftRows_port_state_out_12_2_4), //o
    .port_state_out_12_2_5 (shiftRows_port_state_out_12_2_5), //o
    .port_state_out_12_2_6 (shiftRows_port_state_out_12_2_6), //o
    .port_state_out_12_2_7 (shiftRows_port_state_out_12_2_7), //o
    .port_state_out_12_3_0 (shiftRows_port_state_out_12_3_0), //o
    .port_state_out_12_3_1 (shiftRows_port_state_out_12_3_1), //o
    .port_state_out_12_3_2 (shiftRows_port_state_out_12_3_2), //o
    .port_state_out_12_3_3 (shiftRows_port_state_out_12_3_3), //o
    .port_state_out_12_3_4 (shiftRows_port_state_out_12_3_4), //o
    .port_state_out_12_3_5 (shiftRows_port_state_out_12_3_5), //o
    .port_state_out_12_3_6 (shiftRows_port_state_out_12_3_6), //o
    .port_state_out_12_3_7 (shiftRows_port_state_out_12_3_7), //o
    .port_state_out_13_0_0 (shiftRows_port_state_out_13_0_0), //o
    .port_state_out_13_0_1 (shiftRows_port_state_out_13_0_1), //o
    .port_state_out_13_0_2 (shiftRows_port_state_out_13_0_2), //o
    .port_state_out_13_0_3 (shiftRows_port_state_out_13_0_3), //o
    .port_state_out_13_0_4 (shiftRows_port_state_out_13_0_4), //o
    .port_state_out_13_0_5 (shiftRows_port_state_out_13_0_5), //o
    .port_state_out_13_0_6 (shiftRows_port_state_out_13_0_6), //o
    .port_state_out_13_0_7 (shiftRows_port_state_out_13_0_7), //o
    .port_state_out_13_1_0 (shiftRows_port_state_out_13_1_0), //o
    .port_state_out_13_1_1 (shiftRows_port_state_out_13_1_1), //o
    .port_state_out_13_1_2 (shiftRows_port_state_out_13_1_2), //o
    .port_state_out_13_1_3 (shiftRows_port_state_out_13_1_3), //o
    .port_state_out_13_1_4 (shiftRows_port_state_out_13_1_4), //o
    .port_state_out_13_1_5 (shiftRows_port_state_out_13_1_5), //o
    .port_state_out_13_1_6 (shiftRows_port_state_out_13_1_6), //o
    .port_state_out_13_1_7 (shiftRows_port_state_out_13_1_7), //o
    .port_state_out_13_2_0 (shiftRows_port_state_out_13_2_0), //o
    .port_state_out_13_2_1 (shiftRows_port_state_out_13_2_1), //o
    .port_state_out_13_2_2 (shiftRows_port_state_out_13_2_2), //o
    .port_state_out_13_2_3 (shiftRows_port_state_out_13_2_3), //o
    .port_state_out_13_2_4 (shiftRows_port_state_out_13_2_4), //o
    .port_state_out_13_2_5 (shiftRows_port_state_out_13_2_5), //o
    .port_state_out_13_2_6 (shiftRows_port_state_out_13_2_6), //o
    .port_state_out_13_2_7 (shiftRows_port_state_out_13_2_7), //o
    .port_state_out_13_3_0 (shiftRows_port_state_out_13_3_0), //o
    .port_state_out_13_3_1 (shiftRows_port_state_out_13_3_1), //o
    .port_state_out_13_3_2 (shiftRows_port_state_out_13_3_2), //o
    .port_state_out_13_3_3 (shiftRows_port_state_out_13_3_3), //o
    .port_state_out_13_3_4 (shiftRows_port_state_out_13_3_4), //o
    .port_state_out_13_3_5 (shiftRows_port_state_out_13_3_5), //o
    .port_state_out_13_3_6 (shiftRows_port_state_out_13_3_6), //o
    .port_state_out_13_3_7 (shiftRows_port_state_out_13_3_7), //o
    .port_state_out_14_0_0 (shiftRows_port_state_out_14_0_0), //o
    .port_state_out_14_0_1 (shiftRows_port_state_out_14_0_1), //o
    .port_state_out_14_0_2 (shiftRows_port_state_out_14_0_2), //o
    .port_state_out_14_0_3 (shiftRows_port_state_out_14_0_3), //o
    .port_state_out_14_0_4 (shiftRows_port_state_out_14_0_4), //o
    .port_state_out_14_0_5 (shiftRows_port_state_out_14_0_5), //o
    .port_state_out_14_0_6 (shiftRows_port_state_out_14_0_6), //o
    .port_state_out_14_0_7 (shiftRows_port_state_out_14_0_7), //o
    .port_state_out_14_1_0 (shiftRows_port_state_out_14_1_0), //o
    .port_state_out_14_1_1 (shiftRows_port_state_out_14_1_1), //o
    .port_state_out_14_1_2 (shiftRows_port_state_out_14_1_2), //o
    .port_state_out_14_1_3 (shiftRows_port_state_out_14_1_3), //o
    .port_state_out_14_1_4 (shiftRows_port_state_out_14_1_4), //o
    .port_state_out_14_1_5 (shiftRows_port_state_out_14_1_5), //o
    .port_state_out_14_1_6 (shiftRows_port_state_out_14_1_6), //o
    .port_state_out_14_1_7 (shiftRows_port_state_out_14_1_7), //o
    .port_state_out_14_2_0 (shiftRows_port_state_out_14_2_0), //o
    .port_state_out_14_2_1 (shiftRows_port_state_out_14_2_1), //o
    .port_state_out_14_2_2 (shiftRows_port_state_out_14_2_2), //o
    .port_state_out_14_2_3 (shiftRows_port_state_out_14_2_3), //o
    .port_state_out_14_2_4 (shiftRows_port_state_out_14_2_4), //o
    .port_state_out_14_2_5 (shiftRows_port_state_out_14_2_5), //o
    .port_state_out_14_2_6 (shiftRows_port_state_out_14_2_6), //o
    .port_state_out_14_2_7 (shiftRows_port_state_out_14_2_7), //o
    .port_state_out_14_3_0 (shiftRows_port_state_out_14_3_0), //o
    .port_state_out_14_3_1 (shiftRows_port_state_out_14_3_1), //o
    .port_state_out_14_3_2 (shiftRows_port_state_out_14_3_2), //o
    .port_state_out_14_3_3 (shiftRows_port_state_out_14_3_3), //o
    .port_state_out_14_3_4 (shiftRows_port_state_out_14_3_4), //o
    .port_state_out_14_3_5 (shiftRows_port_state_out_14_3_5), //o
    .port_state_out_14_3_6 (shiftRows_port_state_out_14_3_6), //o
    .port_state_out_14_3_7 (shiftRows_port_state_out_14_3_7), //o
    .port_state_out_15_0_0 (shiftRows_port_state_out_15_0_0), //o
    .port_state_out_15_0_1 (shiftRows_port_state_out_15_0_1), //o
    .port_state_out_15_0_2 (shiftRows_port_state_out_15_0_2), //o
    .port_state_out_15_0_3 (shiftRows_port_state_out_15_0_3), //o
    .port_state_out_15_0_4 (shiftRows_port_state_out_15_0_4), //o
    .port_state_out_15_0_5 (shiftRows_port_state_out_15_0_5), //o
    .port_state_out_15_0_6 (shiftRows_port_state_out_15_0_6), //o
    .port_state_out_15_0_7 (shiftRows_port_state_out_15_0_7), //o
    .port_state_out_15_1_0 (shiftRows_port_state_out_15_1_0), //o
    .port_state_out_15_1_1 (shiftRows_port_state_out_15_1_1), //o
    .port_state_out_15_1_2 (shiftRows_port_state_out_15_1_2), //o
    .port_state_out_15_1_3 (shiftRows_port_state_out_15_1_3), //o
    .port_state_out_15_1_4 (shiftRows_port_state_out_15_1_4), //o
    .port_state_out_15_1_5 (shiftRows_port_state_out_15_1_5), //o
    .port_state_out_15_1_6 (shiftRows_port_state_out_15_1_6), //o
    .port_state_out_15_1_7 (shiftRows_port_state_out_15_1_7), //o
    .port_state_out_15_2_0 (shiftRows_port_state_out_15_2_0), //o
    .port_state_out_15_2_1 (shiftRows_port_state_out_15_2_1), //o
    .port_state_out_15_2_2 (shiftRows_port_state_out_15_2_2), //o
    .port_state_out_15_2_3 (shiftRows_port_state_out_15_2_3), //o
    .port_state_out_15_2_4 (shiftRows_port_state_out_15_2_4), //o
    .port_state_out_15_2_5 (shiftRows_port_state_out_15_2_5), //o
    .port_state_out_15_2_6 (shiftRows_port_state_out_15_2_6), //o
    .port_state_out_15_2_7 (shiftRows_port_state_out_15_2_7), //o
    .port_state_out_15_3_0 (shiftRows_port_state_out_15_3_0), //o
    .port_state_out_15_3_1 (shiftRows_port_state_out_15_3_1), //o
    .port_state_out_15_3_2 (shiftRows_port_state_out_15_3_2), //o
    .port_state_out_15_3_3 (shiftRows_port_state_out_15_3_3), //o
    .port_state_out_15_3_4 (shiftRows_port_state_out_15_3_4), //o
    .port_state_out_15_3_5 (shiftRows_port_state_out_15_3_5), //o
    .port_state_out_15_3_6 (shiftRows_port_state_out_15_3_6), //o
    .port_state_out_15_3_7 (shiftRows_port_state_out_15_3_7)  //o
  );
  Aes_MixColumn mixColumns (
    .port_state_in_0_0_0   (shiftRows_port_state_out_0_0_0  ), //i
    .port_state_in_0_0_1   (shiftRows_port_state_out_0_0_1  ), //i
    .port_state_in_0_0_2   (shiftRows_port_state_out_0_0_2  ), //i
    .port_state_in_0_0_3   (shiftRows_port_state_out_0_0_3  ), //i
    .port_state_in_0_0_4   (shiftRows_port_state_out_0_0_4  ), //i
    .port_state_in_0_0_5   (shiftRows_port_state_out_0_0_5  ), //i
    .port_state_in_0_0_6   (shiftRows_port_state_out_0_0_6  ), //i
    .port_state_in_0_0_7   (shiftRows_port_state_out_0_0_7  ), //i
    .port_state_in_0_1_0   (shiftRows_port_state_out_0_1_0  ), //i
    .port_state_in_0_1_1   (shiftRows_port_state_out_0_1_1  ), //i
    .port_state_in_0_1_2   (shiftRows_port_state_out_0_1_2  ), //i
    .port_state_in_0_1_3   (shiftRows_port_state_out_0_1_3  ), //i
    .port_state_in_0_1_4   (shiftRows_port_state_out_0_1_4  ), //i
    .port_state_in_0_1_5   (shiftRows_port_state_out_0_1_5  ), //i
    .port_state_in_0_1_6   (shiftRows_port_state_out_0_1_6  ), //i
    .port_state_in_0_1_7   (shiftRows_port_state_out_0_1_7  ), //i
    .port_state_in_0_2_0   (shiftRows_port_state_out_0_2_0  ), //i
    .port_state_in_0_2_1   (shiftRows_port_state_out_0_2_1  ), //i
    .port_state_in_0_2_2   (shiftRows_port_state_out_0_2_2  ), //i
    .port_state_in_0_2_3   (shiftRows_port_state_out_0_2_3  ), //i
    .port_state_in_0_2_4   (shiftRows_port_state_out_0_2_4  ), //i
    .port_state_in_0_2_5   (shiftRows_port_state_out_0_2_5  ), //i
    .port_state_in_0_2_6   (shiftRows_port_state_out_0_2_6  ), //i
    .port_state_in_0_2_7   (shiftRows_port_state_out_0_2_7  ), //i
    .port_state_in_0_3_0   (shiftRows_port_state_out_0_3_0  ), //i
    .port_state_in_0_3_1   (shiftRows_port_state_out_0_3_1  ), //i
    .port_state_in_0_3_2   (shiftRows_port_state_out_0_3_2  ), //i
    .port_state_in_0_3_3   (shiftRows_port_state_out_0_3_3  ), //i
    .port_state_in_0_3_4   (shiftRows_port_state_out_0_3_4  ), //i
    .port_state_in_0_3_5   (shiftRows_port_state_out_0_3_5  ), //i
    .port_state_in_0_3_6   (shiftRows_port_state_out_0_3_6  ), //i
    .port_state_in_0_3_7   (shiftRows_port_state_out_0_3_7  ), //i
    .port_state_in_1_0_0   (shiftRows_port_state_out_1_0_0  ), //i
    .port_state_in_1_0_1   (shiftRows_port_state_out_1_0_1  ), //i
    .port_state_in_1_0_2   (shiftRows_port_state_out_1_0_2  ), //i
    .port_state_in_1_0_3   (shiftRows_port_state_out_1_0_3  ), //i
    .port_state_in_1_0_4   (shiftRows_port_state_out_1_0_4  ), //i
    .port_state_in_1_0_5   (shiftRows_port_state_out_1_0_5  ), //i
    .port_state_in_1_0_6   (shiftRows_port_state_out_1_0_6  ), //i
    .port_state_in_1_0_7   (shiftRows_port_state_out_1_0_7  ), //i
    .port_state_in_1_1_0   (shiftRows_port_state_out_1_1_0  ), //i
    .port_state_in_1_1_1   (shiftRows_port_state_out_1_1_1  ), //i
    .port_state_in_1_1_2   (shiftRows_port_state_out_1_1_2  ), //i
    .port_state_in_1_1_3   (shiftRows_port_state_out_1_1_3  ), //i
    .port_state_in_1_1_4   (shiftRows_port_state_out_1_1_4  ), //i
    .port_state_in_1_1_5   (shiftRows_port_state_out_1_1_5  ), //i
    .port_state_in_1_1_6   (shiftRows_port_state_out_1_1_6  ), //i
    .port_state_in_1_1_7   (shiftRows_port_state_out_1_1_7  ), //i
    .port_state_in_1_2_0   (shiftRows_port_state_out_1_2_0  ), //i
    .port_state_in_1_2_1   (shiftRows_port_state_out_1_2_1  ), //i
    .port_state_in_1_2_2   (shiftRows_port_state_out_1_2_2  ), //i
    .port_state_in_1_2_3   (shiftRows_port_state_out_1_2_3  ), //i
    .port_state_in_1_2_4   (shiftRows_port_state_out_1_2_4  ), //i
    .port_state_in_1_2_5   (shiftRows_port_state_out_1_2_5  ), //i
    .port_state_in_1_2_6   (shiftRows_port_state_out_1_2_6  ), //i
    .port_state_in_1_2_7   (shiftRows_port_state_out_1_2_7  ), //i
    .port_state_in_1_3_0   (shiftRows_port_state_out_1_3_0  ), //i
    .port_state_in_1_3_1   (shiftRows_port_state_out_1_3_1  ), //i
    .port_state_in_1_3_2   (shiftRows_port_state_out_1_3_2  ), //i
    .port_state_in_1_3_3   (shiftRows_port_state_out_1_3_3  ), //i
    .port_state_in_1_3_4   (shiftRows_port_state_out_1_3_4  ), //i
    .port_state_in_1_3_5   (shiftRows_port_state_out_1_3_5  ), //i
    .port_state_in_1_3_6   (shiftRows_port_state_out_1_3_6  ), //i
    .port_state_in_1_3_7   (shiftRows_port_state_out_1_3_7  ), //i
    .port_state_in_2_0_0   (shiftRows_port_state_out_2_0_0  ), //i
    .port_state_in_2_0_1   (shiftRows_port_state_out_2_0_1  ), //i
    .port_state_in_2_0_2   (shiftRows_port_state_out_2_0_2  ), //i
    .port_state_in_2_0_3   (shiftRows_port_state_out_2_0_3  ), //i
    .port_state_in_2_0_4   (shiftRows_port_state_out_2_0_4  ), //i
    .port_state_in_2_0_5   (shiftRows_port_state_out_2_0_5  ), //i
    .port_state_in_2_0_6   (shiftRows_port_state_out_2_0_6  ), //i
    .port_state_in_2_0_7   (shiftRows_port_state_out_2_0_7  ), //i
    .port_state_in_2_1_0   (shiftRows_port_state_out_2_1_0  ), //i
    .port_state_in_2_1_1   (shiftRows_port_state_out_2_1_1  ), //i
    .port_state_in_2_1_2   (shiftRows_port_state_out_2_1_2  ), //i
    .port_state_in_2_1_3   (shiftRows_port_state_out_2_1_3  ), //i
    .port_state_in_2_1_4   (shiftRows_port_state_out_2_1_4  ), //i
    .port_state_in_2_1_5   (shiftRows_port_state_out_2_1_5  ), //i
    .port_state_in_2_1_6   (shiftRows_port_state_out_2_1_6  ), //i
    .port_state_in_2_1_7   (shiftRows_port_state_out_2_1_7  ), //i
    .port_state_in_2_2_0   (shiftRows_port_state_out_2_2_0  ), //i
    .port_state_in_2_2_1   (shiftRows_port_state_out_2_2_1  ), //i
    .port_state_in_2_2_2   (shiftRows_port_state_out_2_2_2  ), //i
    .port_state_in_2_2_3   (shiftRows_port_state_out_2_2_3  ), //i
    .port_state_in_2_2_4   (shiftRows_port_state_out_2_2_4  ), //i
    .port_state_in_2_2_5   (shiftRows_port_state_out_2_2_5  ), //i
    .port_state_in_2_2_6   (shiftRows_port_state_out_2_2_6  ), //i
    .port_state_in_2_2_7   (shiftRows_port_state_out_2_2_7  ), //i
    .port_state_in_2_3_0   (shiftRows_port_state_out_2_3_0  ), //i
    .port_state_in_2_3_1   (shiftRows_port_state_out_2_3_1  ), //i
    .port_state_in_2_3_2   (shiftRows_port_state_out_2_3_2  ), //i
    .port_state_in_2_3_3   (shiftRows_port_state_out_2_3_3  ), //i
    .port_state_in_2_3_4   (shiftRows_port_state_out_2_3_4  ), //i
    .port_state_in_2_3_5   (shiftRows_port_state_out_2_3_5  ), //i
    .port_state_in_2_3_6   (shiftRows_port_state_out_2_3_6  ), //i
    .port_state_in_2_3_7   (shiftRows_port_state_out_2_3_7  ), //i
    .port_state_in_3_0_0   (shiftRows_port_state_out_3_0_0  ), //i
    .port_state_in_3_0_1   (shiftRows_port_state_out_3_0_1  ), //i
    .port_state_in_3_0_2   (shiftRows_port_state_out_3_0_2  ), //i
    .port_state_in_3_0_3   (shiftRows_port_state_out_3_0_3  ), //i
    .port_state_in_3_0_4   (shiftRows_port_state_out_3_0_4  ), //i
    .port_state_in_3_0_5   (shiftRows_port_state_out_3_0_5  ), //i
    .port_state_in_3_0_6   (shiftRows_port_state_out_3_0_6  ), //i
    .port_state_in_3_0_7   (shiftRows_port_state_out_3_0_7  ), //i
    .port_state_in_3_1_0   (shiftRows_port_state_out_3_1_0  ), //i
    .port_state_in_3_1_1   (shiftRows_port_state_out_3_1_1  ), //i
    .port_state_in_3_1_2   (shiftRows_port_state_out_3_1_2  ), //i
    .port_state_in_3_1_3   (shiftRows_port_state_out_3_1_3  ), //i
    .port_state_in_3_1_4   (shiftRows_port_state_out_3_1_4  ), //i
    .port_state_in_3_1_5   (shiftRows_port_state_out_3_1_5  ), //i
    .port_state_in_3_1_6   (shiftRows_port_state_out_3_1_6  ), //i
    .port_state_in_3_1_7   (shiftRows_port_state_out_3_1_7  ), //i
    .port_state_in_3_2_0   (shiftRows_port_state_out_3_2_0  ), //i
    .port_state_in_3_2_1   (shiftRows_port_state_out_3_2_1  ), //i
    .port_state_in_3_2_2   (shiftRows_port_state_out_3_2_2  ), //i
    .port_state_in_3_2_3   (shiftRows_port_state_out_3_2_3  ), //i
    .port_state_in_3_2_4   (shiftRows_port_state_out_3_2_4  ), //i
    .port_state_in_3_2_5   (shiftRows_port_state_out_3_2_5  ), //i
    .port_state_in_3_2_6   (shiftRows_port_state_out_3_2_6  ), //i
    .port_state_in_3_2_7   (shiftRows_port_state_out_3_2_7  ), //i
    .port_state_in_3_3_0   (shiftRows_port_state_out_3_3_0  ), //i
    .port_state_in_3_3_1   (shiftRows_port_state_out_3_3_1  ), //i
    .port_state_in_3_3_2   (shiftRows_port_state_out_3_3_2  ), //i
    .port_state_in_3_3_3   (shiftRows_port_state_out_3_3_3  ), //i
    .port_state_in_3_3_4   (shiftRows_port_state_out_3_3_4  ), //i
    .port_state_in_3_3_5   (shiftRows_port_state_out_3_3_5  ), //i
    .port_state_in_3_3_6   (shiftRows_port_state_out_3_3_6  ), //i
    .port_state_in_3_3_7   (shiftRows_port_state_out_3_3_7  ), //i
    .port_state_in_4_0_0   (shiftRows_port_state_out_4_0_0  ), //i
    .port_state_in_4_0_1   (shiftRows_port_state_out_4_0_1  ), //i
    .port_state_in_4_0_2   (shiftRows_port_state_out_4_0_2  ), //i
    .port_state_in_4_0_3   (shiftRows_port_state_out_4_0_3  ), //i
    .port_state_in_4_0_4   (shiftRows_port_state_out_4_0_4  ), //i
    .port_state_in_4_0_5   (shiftRows_port_state_out_4_0_5  ), //i
    .port_state_in_4_0_6   (shiftRows_port_state_out_4_0_6  ), //i
    .port_state_in_4_0_7   (shiftRows_port_state_out_4_0_7  ), //i
    .port_state_in_4_1_0   (shiftRows_port_state_out_4_1_0  ), //i
    .port_state_in_4_1_1   (shiftRows_port_state_out_4_1_1  ), //i
    .port_state_in_4_1_2   (shiftRows_port_state_out_4_1_2  ), //i
    .port_state_in_4_1_3   (shiftRows_port_state_out_4_1_3  ), //i
    .port_state_in_4_1_4   (shiftRows_port_state_out_4_1_4  ), //i
    .port_state_in_4_1_5   (shiftRows_port_state_out_4_1_5  ), //i
    .port_state_in_4_1_6   (shiftRows_port_state_out_4_1_6  ), //i
    .port_state_in_4_1_7   (shiftRows_port_state_out_4_1_7  ), //i
    .port_state_in_4_2_0   (shiftRows_port_state_out_4_2_0  ), //i
    .port_state_in_4_2_1   (shiftRows_port_state_out_4_2_1  ), //i
    .port_state_in_4_2_2   (shiftRows_port_state_out_4_2_2  ), //i
    .port_state_in_4_2_3   (shiftRows_port_state_out_4_2_3  ), //i
    .port_state_in_4_2_4   (shiftRows_port_state_out_4_2_4  ), //i
    .port_state_in_4_2_5   (shiftRows_port_state_out_4_2_5  ), //i
    .port_state_in_4_2_6   (shiftRows_port_state_out_4_2_6  ), //i
    .port_state_in_4_2_7   (shiftRows_port_state_out_4_2_7  ), //i
    .port_state_in_4_3_0   (shiftRows_port_state_out_4_3_0  ), //i
    .port_state_in_4_3_1   (shiftRows_port_state_out_4_3_1  ), //i
    .port_state_in_4_3_2   (shiftRows_port_state_out_4_3_2  ), //i
    .port_state_in_4_3_3   (shiftRows_port_state_out_4_3_3  ), //i
    .port_state_in_4_3_4   (shiftRows_port_state_out_4_3_4  ), //i
    .port_state_in_4_3_5   (shiftRows_port_state_out_4_3_5  ), //i
    .port_state_in_4_3_6   (shiftRows_port_state_out_4_3_6  ), //i
    .port_state_in_4_3_7   (shiftRows_port_state_out_4_3_7  ), //i
    .port_state_in_5_0_0   (shiftRows_port_state_out_5_0_0  ), //i
    .port_state_in_5_0_1   (shiftRows_port_state_out_5_0_1  ), //i
    .port_state_in_5_0_2   (shiftRows_port_state_out_5_0_2  ), //i
    .port_state_in_5_0_3   (shiftRows_port_state_out_5_0_3  ), //i
    .port_state_in_5_0_4   (shiftRows_port_state_out_5_0_4  ), //i
    .port_state_in_5_0_5   (shiftRows_port_state_out_5_0_5  ), //i
    .port_state_in_5_0_6   (shiftRows_port_state_out_5_0_6  ), //i
    .port_state_in_5_0_7   (shiftRows_port_state_out_5_0_7  ), //i
    .port_state_in_5_1_0   (shiftRows_port_state_out_5_1_0  ), //i
    .port_state_in_5_1_1   (shiftRows_port_state_out_5_1_1  ), //i
    .port_state_in_5_1_2   (shiftRows_port_state_out_5_1_2  ), //i
    .port_state_in_5_1_3   (shiftRows_port_state_out_5_1_3  ), //i
    .port_state_in_5_1_4   (shiftRows_port_state_out_5_1_4  ), //i
    .port_state_in_5_1_5   (shiftRows_port_state_out_5_1_5  ), //i
    .port_state_in_5_1_6   (shiftRows_port_state_out_5_1_6  ), //i
    .port_state_in_5_1_7   (shiftRows_port_state_out_5_1_7  ), //i
    .port_state_in_5_2_0   (shiftRows_port_state_out_5_2_0  ), //i
    .port_state_in_5_2_1   (shiftRows_port_state_out_5_2_1  ), //i
    .port_state_in_5_2_2   (shiftRows_port_state_out_5_2_2  ), //i
    .port_state_in_5_2_3   (shiftRows_port_state_out_5_2_3  ), //i
    .port_state_in_5_2_4   (shiftRows_port_state_out_5_2_4  ), //i
    .port_state_in_5_2_5   (shiftRows_port_state_out_5_2_5  ), //i
    .port_state_in_5_2_6   (shiftRows_port_state_out_5_2_6  ), //i
    .port_state_in_5_2_7   (shiftRows_port_state_out_5_2_7  ), //i
    .port_state_in_5_3_0   (shiftRows_port_state_out_5_3_0  ), //i
    .port_state_in_5_3_1   (shiftRows_port_state_out_5_3_1  ), //i
    .port_state_in_5_3_2   (shiftRows_port_state_out_5_3_2  ), //i
    .port_state_in_5_3_3   (shiftRows_port_state_out_5_3_3  ), //i
    .port_state_in_5_3_4   (shiftRows_port_state_out_5_3_4  ), //i
    .port_state_in_5_3_5   (shiftRows_port_state_out_5_3_5  ), //i
    .port_state_in_5_3_6   (shiftRows_port_state_out_5_3_6  ), //i
    .port_state_in_5_3_7   (shiftRows_port_state_out_5_3_7  ), //i
    .port_state_in_6_0_0   (shiftRows_port_state_out_6_0_0  ), //i
    .port_state_in_6_0_1   (shiftRows_port_state_out_6_0_1  ), //i
    .port_state_in_6_0_2   (shiftRows_port_state_out_6_0_2  ), //i
    .port_state_in_6_0_3   (shiftRows_port_state_out_6_0_3  ), //i
    .port_state_in_6_0_4   (shiftRows_port_state_out_6_0_4  ), //i
    .port_state_in_6_0_5   (shiftRows_port_state_out_6_0_5  ), //i
    .port_state_in_6_0_6   (shiftRows_port_state_out_6_0_6  ), //i
    .port_state_in_6_0_7   (shiftRows_port_state_out_6_0_7  ), //i
    .port_state_in_6_1_0   (shiftRows_port_state_out_6_1_0  ), //i
    .port_state_in_6_1_1   (shiftRows_port_state_out_6_1_1  ), //i
    .port_state_in_6_1_2   (shiftRows_port_state_out_6_1_2  ), //i
    .port_state_in_6_1_3   (shiftRows_port_state_out_6_1_3  ), //i
    .port_state_in_6_1_4   (shiftRows_port_state_out_6_1_4  ), //i
    .port_state_in_6_1_5   (shiftRows_port_state_out_6_1_5  ), //i
    .port_state_in_6_1_6   (shiftRows_port_state_out_6_1_6  ), //i
    .port_state_in_6_1_7   (shiftRows_port_state_out_6_1_7  ), //i
    .port_state_in_6_2_0   (shiftRows_port_state_out_6_2_0  ), //i
    .port_state_in_6_2_1   (shiftRows_port_state_out_6_2_1  ), //i
    .port_state_in_6_2_2   (shiftRows_port_state_out_6_2_2  ), //i
    .port_state_in_6_2_3   (shiftRows_port_state_out_6_2_3  ), //i
    .port_state_in_6_2_4   (shiftRows_port_state_out_6_2_4  ), //i
    .port_state_in_6_2_5   (shiftRows_port_state_out_6_2_5  ), //i
    .port_state_in_6_2_6   (shiftRows_port_state_out_6_2_6  ), //i
    .port_state_in_6_2_7   (shiftRows_port_state_out_6_2_7  ), //i
    .port_state_in_6_3_0   (shiftRows_port_state_out_6_3_0  ), //i
    .port_state_in_6_3_1   (shiftRows_port_state_out_6_3_1  ), //i
    .port_state_in_6_3_2   (shiftRows_port_state_out_6_3_2  ), //i
    .port_state_in_6_3_3   (shiftRows_port_state_out_6_3_3  ), //i
    .port_state_in_6_3_4   (shiftRows_port_state_out_6_3_4  ), //i
    .port_state_in_6_3_5   (shiftRows_port_state_out_6_3_5  ), //i
    .port_state_in_6_3_6   (shiftRows_port_state_out_6_3_6  ), //i
    .port_state_in_6_3_7   (shiftRows_port_state_out_6_3_7  ), //i
    .port_state_in_7_0_0   (shiftRows_port_state_out_7_0_0  ), //i
    .port_state_in_7_0_1   (shiftRows_port_state_out_7_0_1  ), //i
    .port_state_in_7_0_2   (shiftRows_port_state_out_7_0_2  ), //i
    .port_state_in_7_0_3   (shiftRows_port_state_out_7_0_3  ), //i
    .port_state_in_7_0_4   (shiftRows_port_state_out_7_0_4  ), //i
    .port_state_in_7_0_5   (shiftRows_port_state_out_7_0_5  ), //i
    .port_state_in_7_0_6   (shiftRows_port_state_out_7_0_6  ), //i
    .port_state_in_7_0_7   (shiftRows_port_state_out_7_0_7  ), //i
    .port_state_in_7_1_0   (shiftRows_port_state_out_7_1_0  ), //i
    .port_state_in_7_1_1   (shiftRows_port_state_out_7_1_1  ), //i
    .port_state_in_7_1_2   (shiftRows_port_state_out_7_1_2  ), //i
    .port_state_in_7_1_3   (shiftRows_port_state_out_7_1_3  ), //i
    .port_state_in_7_1_4   (shiftRows_port_state_out_7_1_4  ), //i
    .port_state_in_7_1_5   (shiftRows_port_state_out_7_1_5  ), //i
    .port_state_in_7_1_6   (shiftRows_port_state_out_7_1_6  ), //i
    .port_state_in_7_1_7   (shiftRows_port_state_out_7_1_7  ), //i
    .port_state_in_7_2_0   (shiftRows_port_state_out_7_2_0  ), //i
    .port_state_in_7_2_1   (shiftRows_port_state_out_7_2_1  ), //i
    .port_state_in_7_2_2   (shiftRows_port_state_out_7_2_2  ), //i
    .port_state_in_7_2_3   (shiftRows_port_state_out_7_2_3  ), //i
    .port_state_in_7_2_4   (shiftRows_port_state_out_7_2_4  ), //i
    .port_state_in_7_2_5   (shiftRows_port_state_out_7_2_5  ), //i
    .port_state_in_7_2_6   (shiftRows_port_state_out_7_2_6  ), //i
    .port_state_in_7_2_7   (shiftRows_port_state_out_7_2_7  ), //i
    .port_state_in_7_3_0   (shiftRows_port_state_out_7_3_0  ), //i
    .port_state_in_7_3_1   (shiftRows_port_state_out_7_3_1  ), //i
    .port_state_in_7_3_2   (shiftRows_port_state_out_7_3_2  ), //i
    .port_state_in_7_3_3   (shiftRows_port_state_out_7_3_3  ), //i
    .port_state_in_7_3_4   (shiftRows_port_state_out_7_3_4  ), //i
    .port_state_in_7_3_5   (shiftRows_port_state_out_7_3_5  ), //i
    .port_state_in_7_3_6   (shiftRows_port_state_out_7_3_6  ), //i
    .port_state_in_7_3_7   (shiftRows_port_state_out_7_3_7  ), //i
    .port_state_in_8_0_0   (shiftRows_port_state_out_8_0_0  ), //i
    .port_state_in_8_0_1   (shiftRows_port_state_out_8_0_1  ), //i
    .port_state_in_8_0_2   (shiftRows_port_state_out_8_0_2  ), //i
    .port_state_in_8_0_3   (shiftRows_port_state_out_8_0_3  ), //i
    .port_state_in_8_0_4   (shiftRows_port_state_out_8_0_4  ), //i
    .port_state_in_8_0_5   (shiftRows_port_state_out_8_0_5  ), //i
    .port_state_in_8_0_6   (shiftRows_port_state_out_8_0_6  ), //i
    .port_state_in_8_0_7   (shiftRows_port_state_out_8_0_7  ), //i
    .port_state_in_8_1_0   (shiftRows_port_state_out_8_1_0  ), //i
    .port_state_in_8_1_1   (shiftRows_port_state_out_8_1_1  ), //i
    .port_state_in_8_1_2   (shiftRows_port_state_out_8_1_2  ), //i
    .port_state_in_8_1_3   (shiftRows_port_state_out_8_1_3  ), //i
    .port_state_in_8_1_4   (shiftRows_port_state_out_8_1_4  ), //i
    .port_state_in_8_1_5   (shiftRows_port_state_out_8_1_5  ), //i
    .port_state_in_8_1_6   (shiftRows_port_state_out_8_1_6  ), //i
    .port_state_in_8_1_7   (shiftRows_port_state_out_8_1_7  ), //i
    .port_state_in_8_2_0   (shiftRows_port_state_out_8_2_0  ), //i
    .port_state_in_8_2_1   (shiftRows_port_state_out_8_2_1  ), //i
    .port_state_in_8_2_2   (shiftRows_port_state_out_8_2_2  ), //i
    .port_state_in_8_2_3   (shiftRows_port_state_out_8_2_3  ), //i
    .port_state_in_8_2_4   (shiftRows_port_state_out_8_2_4  ), //i
    .port_state_in_8_2_5   (shiftRows_port_state_out_8_2_5  ), //i
    .port_state_in_8_2_6   (shiftRows_port_state_out_8_2_6  ), //i
    .port_state_in_8_2_7   (shiftRows_port_state_out_8_2_7  ), //i
    .port_state_in_8_3_0   (shiftRows_port_state_out_8_3_0  ), //i
    .port_state_in_8_3_1   (shiftRows_port_state_out_8_3_1  ), //i
    .port_state_in_8_3_2   (shiftRows_port_state_out_8_3_2  ), //i
    .port_state_in_8_3_3   (shiftRows_port_state_out_8_3_3  ), //i
    .port_state_in_8_3_4   (shiftRows_port_state_out_8_3_4  ), //i
    .port_state_in_8_3_5   (shiftRows_port_state_out_8_3_5  ), //i
    .port_state_in_8_3_6   (shiftRows_port_state_out_8_3_6  ), //i
    .port_state_in_8_3_7   (shiftRows_port_state_out_8_3_7  ), //i
    .port_state_in_9_0_0   (shiftRows_port_state_out_9_0_0  ), //i
    .port_state_in_9_0_1   (shiftRows_port_state_out_9_0_1  ), //i
    .port_state_in_9_0_2   (shiftRows_port_state_out_9_0_2  ), //i
    .port_state_in_9_0_3   (shiftRows_port_state_out_9_0_3  ), //i
    .port_state_in_9_0_4   (shiftRows_port_state_out_9_0_4  ), //i
    .port_state_in_9_0_5   (shiftRows_port_state_out_9_0_5  ), //i
    .port_state_in_9_0_6   (shiftRows_port_state_out_9_0_6  ), //i
    .port_state_in_9_0_7   (shiftRows_port_state_out_9_0_7  ), //i
    .port_state_in_9_1_0   (shiftRows_port_state_out_9_1_0  ), //i
    .port_state_in_9_1_1   (shiftRows_port_state_out_9_1_1  ), //i
    .port_state_in_9_1_2   (shiftRows_port_state_out_9_1_2  ), //i
    .port_state_in_9_1_3   (shiftRows_port_state_out_9_1_3  ), //i
    .port_state_in_9_1_4   (shiftRows_port_state_out_9_1_4  ), //i
    .port_state_in_9_1_5   (shiftRows_port_state_out_9_1_5  ), //i
    .port_state_in_9_1_6   (shiftRows_port_state_out_9_1_6  ), //i
    .port_state_in_9_1_7   (shiftRows_port_state_out_9_1_7  ), //i
    .port_state_in_9_2_0   (shiftRows_port_state_out_9_2_0  ), //i
    .port_state_in_9_2_1   (shiftRows_port_state_out_9_2_1  ), //i
    .port_state_in_9_2_2   (shiftRows_port_state_out_9_2_2  ), //i
    .port_state_in_9_2_3   (shiftRows_port_state_out_9_2_3  ), //i
    .port_state_in_9_2_4   (shiftRows_port_state_out_9_2_4  ), //i
    .port_state_in_9_2_5   (shiftRows_port_state_out_9_2_5  ), //i
    .port_state_in_9_2_6   (shiftRows_port_state_out_9_2_6  ), //i
    .port_state_in_9_2_7   (shiftRows_port_state_out_9_2_7  ), //i
    .port_state_in_9_3_0   (shiftRows_port_state_out_9_3_0  ), //i
    .port_state_in_9_3_1   (shiftRows_port_state_out_9_3_1  ), //i
    .port_state_in_9_3_2   (shiftRows_port_state_out_9_3_2  ), //i
    .port_state_in_9_3_3   (shiftRows_port_state_out_9_3_3  ), //i
    .port_state_in_9_3_4   (shiftRows_port_state_out_9_3_4  ), //i
    .port_state_in_9_3_5   (shiftRows_port_state_out_9_3_5  ), //i
    .port_state_in_9_3_6   (shiftRows_port_state_out_9_3_6  ), //i
    .port_state_in_9_3_7   (shiftRows_port_state_out_9_3_7  ), //i
    .port_state_in_10_0_0  (shiftRows_port_state_out_10_0_0 ), //i
    .port_state_in_10_0_1  (shiftRows_port_state_out_10_0_1 ), //i
    .port_state_in_10_0_2  (shiftRows_port_state_out_10_0_2 ), //i
    .port_state_in_10_0_3  (shiftRows_port_state_out_10_0_3 ), //i
    .port_state_in_10_0_4  (shiftRows_port_state_out_10_0_4 ), //i
    .port_state_in_10_0_5  (shiftRows_port_state_out_10_0_5 ), //i
    .port_state_in_10_0_6  (shiftRows_port_state_out_10_0_6 ), //i
    .port_state_in_10_0_7  (shiftRows_port_state_out_10_0_7 ), //i
    .port_state_in_10_1_0  (shiftRows_port_state_out_10_1_0 ), //i
    .port_state_in_10_1_1  (shiftRows_port_state_out_10_1_1 ), //i
    .port_state_in_10_1_2  (shiftRows_port_state_out_10_1_2 ), //i
    .port_state_in_10_1_3  (shiftRows_port_state_out_10_1_3 ), //i
    .port_state_in_10_1_4  (shiftRows_port_state_out_10_1_4 ), //i
    .port_state_in_10_1_5  (shiftRows_port_state_out_10_1_5 ), //i
    .port_state_in_10_1_6  (shiftRows_port_state_out_10_1_6 ), //i
    .port_state_in_10_1_7  (shiftRows_port_state_out_10_1_7 ), //i
    .port_state_in_10_2_0  (shiftRows_port_state_out_10_2_0 ), //i
    .port_state_in_10_2_1  (shiftRows_port_state_out_10_2_1 ), //i
    .port_state_in_10_2_2  (shiftRows_port_state_out_10_2_2 ), //i
    .port_state_in_10_2_3  (shiftRows_port_state_out_10_2_3 ), //i
    .port_state_in_10_2_4  (shiftRows_port_state_out_10_2_4 ), //i
    .port_state_in_10_2_5  (shiftRows_port_state_out_10_2_5 ), //i
    .port_state_in_10_2_6  (shiftRows_port_state_out_10_2_6 ), //i
    .port_state_in_10_2_7  (shiftRows_port_state_out_10_2_7 ), //i
    .port_state_in_10_3_0  (shiftRows_port_state_out_10_3_0 ), //i
    .port_state_in_10_3_1  (shiftRows_port_state_out_10_3_1 ), //i
    .port_state_in_10_3_2  (shiftRows_port_state_out_10_3_2 ), //i
    .port_state_in_10_3_3  (shiftRows_port_state_out_10_3_3 ), //i
    .port_state_in_10_3_4  (shiftRows_port_state_out_10_3_4 ), //i
    .port_state_in_10_3_5  (shiftRows_port_state_out_10_3_5 ), //i
    .port_state_in_10_3_6  (shiftRows_port_state_out_10_3_6 ), //i
    .port_state_in_10_3_7  (shiftRows_port_state_out_10_3_7 ), //i
    .port_state_in_11_0_0  (shiftRows_port_state_out_11_0_0 ), //i
    .port_state_in_11_0_1  (shiftRows_port_state_out_11_0_1 ), //i
    .port_state_in_11_0_2  (shiftRows_port_state_out_11_0_2 ), //i
    .port_state_in_11_0_3  (shiftRows_port_state_out_11_0_3 ), //i
    .port_state_in_11_0_4  (shiftRows_port_state_out_11_0_4 ), //i
    .port_state_in_11_0_5  (shiftRows_port_state_out_11_0_5 ), //i
    .port_state_in_11_0_6  (shiftRows_port_state_out_11_0_6 ), //i
    .port_state_in_11_0_7  (shiftRows_port_state_out_11_0_7 ), //i
    .port_state_in_11_1_0  (shiftRows_port_state_out_11_1_0 ), //i
    .port_state_in_11_1_1  (shiftRows_port_state_out_11_1_1 ), //i
    .port_state_in_11_1_2  (shiftRows_port_state_out_11_1_2 ), //i
    .port_state_in_11_1_3  (shiftRows_port_state_out_11_1_3 ), //i
    .port_state_in_11_1_4  (shiftRows_port_state_out_11_1_4 ), //i
    .port_state_in_11_1_5  (shiftRows_port_state_out_11_1_5 ), //i
    .port_state_in_11_1_6  (shiftRows_port_state_out_11_1_6 ), //i
    .port_state_in_11_1_7  (shiftRows_port_state_out_11_1_7 ), //i
    .port_state_in_11_2_0  (shiftRows_port_state_out_11_2_0 ), //i
    .port_state_in_11_2_1  (shiftRows_port_state_out_11_2_1 ), //i
    .port_state_in_11_2_2  (shiftRows_port_state_out_11_2_2 ), //i
    .port_state_in_11_2_3  (shiftRows_port_state_out_11_2_3 ), //i
    .port_state_in_11_2_4  (shiftRows_port_state_out_11_2_4 ), //i
    .port_state_in_11_2_5  (shiftRows_port_state_out_11_2_5 ), //i
    .port_state_in_11_2_6  (shiftRows_port_state_out_11_2_6 ), //i
    .port_state_in_11_2_7  (shiftRows_port_state_out_11_2_7 ), //i
    .port_state_in_11_3_0  (shiftRows_port_state_out_11_3_0 ), //i
    .port_state_in_11_3_1  (shiftRows_port_state_out_11_3_1 ), //i
    .port_state_in_11_3_2  (shiftRows_port_state_out_11_3_2 ), //i
    .port_state_in_11_3_3  (shiftRows_port_state_out_11_3_3 ), //i
    .port_state_in_11_3_4  (shiftRows_port_state_out_11_3_4 ), //i
    .port_state_in_11_3_5  (shiftRows_port_state_out_11_3_5 ), //i
    .port_state_in_11_3_6  (shiftRows_port_state_out_11_3_6 ), //i
    .port_state_in_11_3_7  (shiftRows_port_state_out_11_3_7 ), //i
    .port_state_in_12_0_0  (shiftRows_port_state_out_12_0_0 ), //i
    .port_state_in_12_0_1  (shiftRows_port_state_out_12_0_1 ), //i
    .port_state_in_12_0_2  (shiftRows_port_state_out_12_0_2 ), //i
    .port_state_in_12_0_3  (shiftRows_port_state_out_12_0_3 ), //i
    .port_state_in_12_0_4  (shiftRows_port_state_out_12_0_4 ), //i
    .port_state_in_12_0_5  (shiftRows_port_state_out_12_0_5 ), //i
    .port_state_in_12_0_6  (shiftRows_port_state_out_12_0_6 ), //i
    .port_state_in_12_0_7  (shiftRows_port_state_out_12_0_7 ), //i
    .port_state_in_12_1_0  (shiftRows_port_state_out_12_1_0 ), //i
    .port_state_in_12_1_1  (shiftRows_port_state_out_12_1_1 ), //i
    .port_state_in_12_1_2  (shiftRows_port_state_out_12_1_2 ), //i
    .port_state_in_12_1_3  (shiftRows_port_state_out_12_1_3 ), //i
    .port_state_in_12_1_4  (shiftRows_port_state_out_12_1_4 ), //i
    .port_state_in_12_1_5  (shiftRows_port_state_out_12_1_5 ), //i
    .port_state_in_12_1_6  (shiftRows_port_state_out_12_1_6 ), //i
    .port_state_in_12_1_7  (shiftRows_port_state_out_12_1_7 ), //i
    .port_state_in_12_2_0  (shiftRows_port_state_out_12_2_0 ), //i
    .port_state_in_12_2_1  (shiftRows_port_state_out_12_2_1 ), //i
    .port_state_in_12_2_2  (shiftRows_port_state_out_12_2_2 ), //i
    .port_state_in_12_2_3  (shiftRows_port_state_out_12_2_3 ), //i
    .port_state_in_12_2_4  (shiftRows_port_state_out_12_2_4 ), //i
    .port_state_in_12_2_5  (shiftRows_port_state_out_12_2_5 ), //i
    .port_state_in_12_2_6  (shiftRows_port_state_out_12_2_6 ), //i
    .port_state_in_12_2_7  (shiftRows_port_state_out_12_2_7 ), //i
    .port_state_in_12_3_0  (shiftRows_port_state_out_12_3_0 ), //i
    .port_state_in_12_3_1  (shiftRows_port_state_out_12_3_1 ), //i
    .port_state_in_12_3_2  (shiftRows_port_state_out_12_3_2 ), //i
    .port_state_in_12_3_3  (shiftRows_port_state_out_12_3_3 ), //i
    .port_state_in_12_3_4  (shiftRows_port_state_out_12_3_4 ), //i
    .port_state_in_12_3_5  (shiftRows_port_state_out_12_3_5 ), //i
    .port_state_in_12_3_6  (shiftRows_port_state_out_12_3_6 ), //i
    .port_state_in_12_3_7  (shiftRows_port_state_out_12_3_7 ), //i
    .port_state_in_13_0_0  (shiftRows_port_state_out_13_0_0 ), //i
    .port_state_in_13_0_1  (shiftRows_port_state_out_13_0_1 ), //i
    .port_state_in_13_0_2  (shiftRows_port_state_out_13_0_2 ), //i
    .port_state_in_13_0_3  (shiftRows_port_state_out_13_0_3 ), //i
    .port_state_in_13_0_4  (shiftRows_port_state_out_13_0_4 ), //i
    .port_state_in_13_0_5  (shiftRows_port_state_out_13_0_5 ), //i
    .port_state_in_13_0_6  (shiftRows_port_state_out_13_0_6 ), //i
    .port_state_in_13_0_7  (shiftRows_port_state_out_13_0_7 ), //i
    .port_state_in_13_1_0  (shiftRows_port_state_out_13_1_0 ), //i
    .port_state_in_13_1_1  (shiftRows_port_state_out_13_1_1 ), //i
    .port_state_in_13_1_2  (shiftRows_port_state_out_13_1_2 ), //i
    .port_state_in_13_1_3  (shiftRows_port_state_out_13_1_3 ), //i
    .port_state_in_13_1_4  (shiftRows_port_state_out_13_1_4 ), //i
    .port_state_in_13_1_5  (shiftRows_port_state_out_13_1_5 ), //i
    .port_state_in_13_1_6  (shiftRows_port_state_out_13_1_6 ), //i
    .port_state_in_13_1_7  (shiftRows_port_state_out_13_1_7 ), //i
    .port_state_in_13_2_0  (shiftRows_port_state_out_13_2_0 ), //i
    .port_state_in_13_2_1  (shiftRows_port_state_out_13_2_1 ), //i
    .port_state_in_13_2_2  (shiftRows_port_state_out_13_2_2 ), //i
    .port_state_in_13_2_3  (shiftRows_port_state_out_13_2_3 ), //i
    .port_state_in_13_2_4  (shiftRows_port_state_out_13_2_4 ), //i
    .port_state_in_13_2_5  (shiftRows_port_state_out_13_2_5 ), //i
    .port_state_in_13_2_6  (shiftRows_port_state_out_13_2_6 ), //i
    .port_state_in_13_2_7  (shiftRows_port_state_out_13_2_7 ), //i
    .port_state_in_13_3_0  (shiftRows_port_state_out_13_3_0 ), //i
    .port_state_in_13_3_1  (shiftRows_port_state_out_13_3_1 ), //i
    .port_state_in_13_3_2  (shiftRows_port_state_out_13_3_2 ), //i
    .port_state_in_13_3_3  (shiftRows_port_state_out_13_3_3 ), //i
    .port_state_in_13_3_4  (shiftRows_port_state_out_13_3_4 ), //i
    .port_state_in_13_3_5  (shiftRows_port_state_out_13_3_5 ), //i
    .port_state_in_13_3_6  (shiftRows_port_state_out_13_3_6 ), //i
    .port_state_in_13_3_7  (shiftRows_port_state_out_13_3_7 ), //i
    .port_state_in_14_0_0  (shiftRows_port_state_out_14_0_0 ), //i
    .port_state_in_14_0_1  (shiftRows_port_state_out_14_0_1 ), //i
    .port_state_in_14_0_2  (shiftRows_port_state_out_14_0_2 ), //i
    .port_state_in_14_0_3  (shiftRows_port_state_out_14_0_3 ), //i
    .port_state_in_14_0_4  (shiftRows_port_state_out_14_0_4 ), //i
    .port_state_in_14_0_5  (shiftRows_port_state_out_14_0_5 ), //i
    .port_state_in_14_0_6  (shiftRows_port_state_out_14_0_6 ), //i
    .port_state_in_14_0_7  (shiftRows_port_state_out_14_0_7 ), //i
    .port_state_in_14_1_0  (shiftRows_port_state_out_14_1_0 ), //i
    .port_state_in_14_1_1  (shiftRows_port_state_out_14_1_1 ), //i
    .port_state_in_14_1_2  (shiftRows_port_state_out_14_1_2 ), //i
    .port_state_in_14_1_3  (shiftRows_port_state_out_14_1_3 ), //i
    .port_state_in_14_1_4  (shiftRows_port_state_out_14_1_4 ), //i
    .port_state_in_14_1_5  (shiftRows_port_state_out_14_1_5 ), //i
    .port_state_in_14_1_6  (shiftRows_port_state_out_14_1_6 ), //i
    .port_state_in_14_1_7  (shiftRows_port_state_out_14_1_7 ), //i
    .port_state_in_14_2_0  (shiftRows_port_state_out_14_2_0 ), //i
    .port_state_in_14_2_1  (shiftRows_port_state_out_14_2_1 ), //i
    .port_state_in_14_2_2  (shiftRows_port_state_out_14_2_2 ), //i
    .port_state_in_14_2_3  (shiftRows_port_state_out_14_2_3 ), //i
    .port_state_in_14_2_4  (shiftRows_port_state_out_14_2_4 ), //i
    .port_state_in_14_2_5  (shiftRows_port_state_out_14_2_5 ), //i
    .port_state_in_14_2_6  (shiftRows_port_state_out_14_2_6 ), //i
    .port_state_in_14_2_7  (shiftRows_port_state_out_14_2_7 ), //i
    .port_state_in_14_3_0  (shiftRows_port_state_out_14_3_0 ), //i
    .port_state_in_14_3_1  (shiftRows_port_state_out_14_3_1 ), //i
    .port_state_in_14_3_2  (shiftRows_port_state_out_14_3_2 ), //i
    .port_state_in_14_3_3  (shiftRows_port_state_out_14_3_3 ), //i
    .port_state_in_14_3_4  (shiftRows_port_state_out_14_3_4 ), //i
    .port_state_in_14_3_5  (shiftRows_port_state_out_14_3_5 ), //i
    .port_state_in_14_3_6  (shiftRows_port_state_out_14_3_6 ), //i
    .port_state_in_14_3_7  (shiftRows_port_state_out_14_3_7 ), //i
    .port_state_in_15_0_0  (shiftRows_port_state_out_15_0_0 ), //i
    .port_state_in_15_0_1  (shiftRows_port_state_out_15_0_1 ), //i
    .port_state_in_15_0_2  (shiftRows_port_state_out_15_0_2 ), //i
    .port_state_in_15_0_3  (shiftRows_port_state_out_15_0_3 ), //i
    .port_state_in_15_0_4  (shiftRows_port_state_out_15_0_4 ), //i
    .port_state_in_15_0_5  (shiftRows_port_state_out_15_0_5 ), //i
    .port_state_in_15_0_6  (shiftRows_port_state_out_15_0_6 ), //i
    .port_state_in_15_0_7  (shiftRows_port_state_out_15_0_7 ), //i
    .port_state_in_15_1_0  (shiftRows_port_state_out_15_1_0 ), //i
    .port_state_in_15_1_1  (shiftRows_port_state_out_15_1_1 ), //i
    .port_state_in_15_1_2  (shiftRows_port_state_out_15_1_2 ), //i
    .port_state_in_15_1_3  (shiftRows_port_state_out_15_1_3 ), //i
    .port_state_in_15_1_4  (shiftRows_port_state_out_15_1_4 ), //i
    .port_state_in_15_1_5  (shiftRows_port_state_out_15_1_5 ), //i
    .port_state_in_15_1_6  (shiftRows_port_state_out_15_1_6 ), //i
    .port_state_in_15_1_7  (shiftRows_port_state_out_15_1_7 ), //i
    .port_state_in_15_2_0  (shiftRows_port_state_out_15_2_0 ), //i
    .port_state_in_15_2_1  (shiftRows_port_state_out_15_2_1 ), //i
    .port_state_in_15_2_2  (shiftRows_port_state_out_15_2_2 ), //i
    .port_state_in_15_2_3  (shiftRows_port_state_out_15_2_3 ), //i
    .port_state_in_15_2_4  (shiftRows_port_state_out_15_2_4 ), //i
    .port_state_in_15_2_5  (shiftRows_port_state_out_15_2_5 ), //i
    .port_state_in_15_2_6  (shiftRows_port_state_out_15_2_6 ), //i
    .port_state_in_15_2_7  (shiftRows_port_state_out_15_2_7 ), //i
    .port_state_in_15_3_0  (shiftRows_port_state_out_15_3_0 ), //i
    .port_state_in_15_3_1  (shiftRows_port_state_out_15_3_1 ), //i
    .port_state_in_15_3_2  (shiftRows_port_state_out_15_3_2 ), //i
    .port_state_in_15_3_3  (shiftRows_port_state_out_15_3_3 ), //i
    .port_state_in_15_3_4  (shiftRows_port_state_out_15_3_4 ), //i
    .port_state_in_15_3_5  (shiftRows_port_state_out_15_3_5 ), //i
    .port_state_in_15_3_6  (shiftRows_port_state_out_15_3_6 ), //i
    .port_state_in_15_3_7  (shiftRows_port_state_out_15_3_7 ), //i
    .port_state_out_0_0_0  (mixColumns_port_state_out_0_0_0 ), //o
    .port_state_out_0_0_1  (mixColumns_port_state_out_0_0_1 ), //o
    .port_state_out_0_0_2  (mixColumns_port_state_out_0_0_2 ), //o
    .port_state_out_0_0_3  (mixColumns_port_state_out_0_0_3 ), //o
    .port_state_out_0_0_4  (mixColumns_port_state_out_0_0_4 ), //o
    .port_state_out_0_0_5  (mixColumns_port_state_out_0_0_5 ), //o
    .port_state_out_0_0_6  (mixColumns_port_state_out_0_0_6 ), //o
    .port_state_out_0_0_7  (mixColumns_port_state_out_0_0_7 ), //o
    .port_state_out_0_1_0  (mixColumns_port_state_out_0_1_0 ), //o
    .port_state_out_0_1_1  (mixColumns_port_state_out_0_1_1 ), //o
    .port_state_out_0_1_2  (mixColumns_port_state_out_0_1_2 ), //o
    .port_state_out_0_1_3  (mixColumns_port_state_out_0_1_3 ), //o
    .port_state_out_0_1_4  (mixColumns_port_state_out_0_1_4 ), //o
    .port_state_out_0_1_5  (mixColumns_port_state_out_0_1_5 ), //o
    .port_state_out_0_1_6  (mixColumns_port_state_out_0_1_6 ), //o
    .port_state_out_0_1_7  (mixColumns_port_state_out_0_1_7 ), //o
    .port_state_out_0_2_0  (mixColumns_port_state_out_0_2_0 ), //o
    .port_state_out_0_2_1  (mixColumns_port_state_out_0_2_1 ), //o
    .port_state_out_0_2_2  (mixColumns_port_state_out_0_2_2 ), //o
    .port_state_out_0_2_3  (mixColumns_port_state_out_0_2_3 ), //o
    .port_state_out_0_2_4  (mixColumns_port_state_out_0_2_4 ), //o
    .port_state_out_0_2_5  (mixColumns_port_state_out_0_2_5 ), //o
    .port_state_out_0_2_6  (mixColumns_port_state_out_0_2_6 ), //o
    .port_state_out_0_2_7  (mixColumns_port_state_out_0_2_7 ), //o
    .port_state_out_0_3_0  (mixColumns_port_state_out_0_3_0 ), //o
    .port_state_out_0_3_1  (mixColumns_port_state_out_0_3_1 ), //o
    .port_state_out_0_3_2  (mixColumns_port_state_out_0_3_2 ), //o
    .port_state_out_0_3_3  (mixColumns_port_state_out_0_3_3 ), //o
    .port_state_out_0_3_4  (mixColumns_port_state_out_0_3_4 ), //o
    .port_state_out_0_3_5  (mixColumns_port_state_out_0_3_5 ), //o
    .port_state_out_0_3_6  (mixColumns_port_state_out_0_3_6 ), //o
    .port_state_out_0_3_7  (mixColumns_port_state_out_0_3_7 ), //o
    .port_state_out_1_0_0  (mixColumns_port_state_out_1_0_0 ), //o
    .port_state_out_1_0_1  (mixColumns_port_state_out_1_0_1 ), //o
    .port_state_out_1_0_2  (mixColumns_port_state_out_1_0_2 ), //o
    .port_state_out_1_0_3  (mixColumns_port_state_out_1_0_3 ), //o
    .port_state_out_1_0_4  (mixColumns_port_state_out_1_0_4 ), //o
    .port_state_out_1_0_5  (mixColumns_port_state_out_1_0_5 ), //o
    .port_state_out_1_0_6  (mixColumns_port_state_out_1_0_6 ), //o
    .port_state_out_1_0_7  (mixColumns_port_state_out_1_0_7 ), //o
    .port_state_out_1_1_0  (mixColumns_port_state_out_1_1_0 ), //o
    .port_state_out_1_1_1  (mixColumns_port_state_out_1_1_1 ), //o
    .port_state_out_1_1_2  (mixColumns_port_state_out_1_1_2 ), //o
    .port_state_out_1_1_3  (mixColumns_port_state_out_1_1_3 ), //o
    .port_state_out_1_1_4  (mixColumns_port_state_out_1_1_4 ), //o
    .port_state_out_1_1_5  (mixColumns_port_state_out_1_1_5 ), //o
    .port_state_out_1_1_6  (mixColumns_port_state_out_1_1_6 ), //o
    .port_state_out_1_1_7  (mixColumns_port_state_out_1_1_7 ), //o
    .port_state_out_1_2_0  (mixColumns_port_state_out_1_2_0 ), //o
    .port_state_out_1_2_1  (mixColumns_port_state_out_1_2_1 ), //o
    .port_state_out_1_2_2  (mixColumns_port_state_out_1_2_2 ), //o
    .port_state_out_1_2_3  (mixColumns_port_state_out_1_2_3 ), //o
    .port_state_out_1_2_4  (mixColumns_port_state_out_1_2_4 ), //o
    .port_state_out_1_2_5  (mixColumns_port_state_out_1_2_5 ), //o
    .port_state_out_1_2_6  (mixColumns_port_state_out_1_2_6 ), //o
    .port_state_out_1_2_7  (mixColumns_port_state_out_1_2_7 ), //o
    .port_state_out_1_3_0  (mixColumns_port_state_out_1_3_0 ), //o
    .port_state_out_1_3_1  (mixColumns_port_state_out_1_3_1 ), //o
    .port_state_out_1_3_2  (mixColumns_port_state_out_1_3_2 ), //o
    .port_state_out_1_3_3  (mixColumns_port_state_out_1_3_3 ), //o
    .port_state_out_1_3_4  (mixColumns_port_state_out_1_3_4 ), //o
    .port_state_out_1_3_5  (mixColumns_port_state_out_1_3_5 ), //o
    .port_state_out_1_3_6  (mixColumns_port_state_out_1_3_6 ), //o
    .port_state_out_1_3_7  (mixColumns_port_state_out_1_3_7 ), //o
    .port_state_out_2_0_0  (mixColumns_port_state_out_2_0_0 ), //o
    .port_state_out_2_0_1  (mixColumns_port_state_out_2_0_1 ), //o
    .port_state_out_2_0_2  (mixColumns_port_state_out_2_0_2 ), //o
    .port_state_out_2_0_3  (mixColumns_port_state_out_2_0_3 ), //o
    .port_state_out_2_0_4  (mixColumns_port_state_out_2_0_4 ), //o
    .port_state_out_2_0_5  (mixColumns_port_state_out_2_0_5 ), //o
    .port_state_out_2_0_6  (mixColumns_port_state_out_2_0_6 ), //o
    .port_state_out_2_0_7  (mixColumns_port_state_out_2_0_7 ), //o
    .port_state_out_2_1_0  (mixColumns_port_state_out_2_1_0 ), //o
    .port_state_out_2_1_1  (mixColumns_port_state_out_2_1_1 ), //o
    .port_state_out_2_1_2  (mixColumns_port_state_out_2_1_2 ), //o
    .port_state_out_2_1_3  (mixColumns_port_state_out_2_1_3 ), //o
    .port_state_out_2_1_4  (mixColumns_port_state_out_2_1_4 ), //o
    .port_state_out_2_1_5  (mixColumns_port_state_out_2_1_5 ), //o
    .port_state_out_2_1_6  (mixColumns_port_state_out_2_1_6 ), //o
    .port_state_out_2_1_7  (mixColumns_port_state_out_2_1_7 ), //o
    .port_state_out_2_2_0  (mixColumns_port_state_out_2_2_0 ), //o
    .port_state_out_2_2_1  (mixColumns_port_state_out_2_2_1 ), //o
    .port_state_out_2_2_2  (mixColumns_port_state_out_2_2_2 ), //o
    .port_state_out_2_2_3  (mixColumns_port_state_out_2_2_3 ), //o
    .port_state_out_2_2_4  (mixColumns_port_state_out_2_2_4 ), //o
    .port_state_out_2_2_5  (mixColumns_port_state_out_2_2_5 ), //o
    .port_state_out_2_2_6  (mixColumns_port_state_out_2_2_6 ), //o
    .port_state_out_2_2_7  (mixColumns_port_state_out_2_2_7 ), //o
    .port_state_out_2_3_0  (mixColumns_port_state_out_2_3_0 ), //o
    .port_state_out_2_3_1  (mixColumns_port_state_out_2_3_1 ), //o
    .port_state_out_2_3_2  (mixColumns_port_state_out_2_3_2 ), //o
    .port_state_out_2_3_3  (mixColumns_port_state_out_2_3_3 ), //o
    .port_state_out_2_3_4  (mixColumns_port_state_out_2_3_4 ), //o
    .port_state_out_2_3_5  (mixColumns_port_state_out_2_3_5 ), //o
    .port_state_out_2_3_6  (mixColumns_port_state_out_2_3_6 ), //o
    .port_state_out_2_3_7  (mixColumns_port_state_out_2_3_7 ), //o
    .port_state_out_3_0_0  (mixColumns_port_state_out_3_0_0 ), //o
    .port_state_out_3_0_1  (mixColumns_port_state_out_3_0_1 ), //o
    .port_state_out_3_0_2  (mixColumns_port_state_out_3_0_2 ), //o
    .port_state_out_3_0_3  (mixColumns_port_state_out_3_0_3 ), //o
    .port_state_out_3_0_4  (mixColumns_port_state_out_3_0_4 ), //o
    .port_state_out_3_0_5  (mixColumns_port_state_out_3_0_5 ), //o
    .port_state_out_3_0_6  (mixColumns_port_state_out_3_0_6 ), //o
    .port_state_out_3_0_7  (mixColumns_port_state_out_3_0_7 ), //o
    .port_state_out_3_1_0  (mixColumns_port_state_out_3_1_0 ), //o
    .port_state_out_3_1_1  (mixColumns_port_state_out_3_1_1 ), //o
    .port_state_out_3_1_2  (mixColumns_port_state_out_3_1_2 ), //o
    .port_state_out_3_1_3  (mixColumns_port_state_out_3_1_3 ), //o
    .port_state_out_3_1_4  (mixColumns_port_state_out_3_1_4 ), //o
    .port_state_out_3_1_5  (mixColumns_port_state_out_3_1_5 ), //o
    .port_state_out_3_1_6  (mixColumns_port_state_out_3_1_6 ), //o
    .port_state_out_3_1_7  (mixColumns_port_state_out_3_1_7 ), //o
    .port_state_out_3_2_0  (mixColumns_port_state_out_3_2_0 ), //o
    .port_state_out_3_2_1  (mixColumns_port_state_out_3_2_1 ), //o
    .port_state_out_3_2_2  (mixColumns_port_state_out_3_2_2 ), //o
    .port_state_out_3_2_3  (mixColumns_port_state_out_3_2_3 ), //o
    .port_state_out_3_2_4  (mixColumns_port_state_out_3_2_4 ), //o
    .port_state_out_3_2_5  (mixColumns_port_state_out_3_2_5 ), //o
    .port_state_out_3_2_6  (mixColumns_port_state_out_3_2_6 ), //o
    .port_state_out_3_2_7  (mixColumns_port_state_out_3_2_7 ), //o
    .port_state_out_3_3_0  (mixColumns_port_state_out_3_3_0 ), //o
    .port_state_out_3_3_1  (mixColumns_port_state_out_3_3_1 ), //o
    .port_state_out_3_3_2  (mixColumns_port_state_out_3_3_2 ), //o
    .port_state_out_3_3_3  (mixColumns_port_state_out_3_3_3 ), //o
    .port_state_out_3_3_4  (mixColumns_port_state_out_3_3_4 ), //o
    .port_state_out_3_3_5  (mixColumns_port_state_out_3_3_5 ), //o
    .port_state_out_3_3_6  (mixColumns_port_state_out_3_3_6 ), //o
    .port_state_out_3_3_7  (mixColumns_port_state_out_3_3_7 ), //o
    .port_state_out_4_0_0  (mixColumns_port_state_out_4_0_0 ), //o
    .port_state_out_4_0_1  (mixColumns_port_state_out_4_0_1 ), //o
    .port_state_out_4_0_2  (mixColumns_port_state_out_4_0_2 ), //o
    .port_state_out_4_0_3  (mixColumns_port_state_out_4_0_3 ), //o
    .port_state_out_4_0_4  (mixColumns_port_state_out_4_0_4 ), //o
    .port_state_out_4_0_5  (mixColumns_port_state_out_4_0_5 ), //o
    .port_state_out_4_0_6  (mixColumns_port_state_out_4_0_6 ), //o
    .port_state_out_4_0_7  (mixColumns_port_state_out_4_0_7 ), //o
    .port_state_out_4_1_0  (mixColumns_port_state_out_4_1_0 ), //o
    .port_state_out_4_1_1  (mixColumns_port_state_out_4_1_1 ), //o
    .port_state_out_4_1_2  (mixColumns_port_state_out_4_1_2 ), //o
    .port_state_out_4_1_3  (mixColumns_port_state_out_4_1_3 ), //o
    .port_state_out_4_1_4  (mixColumns_port_state_out_4_1_4 ), //o
    .port_state_out_4_1_5  (mixColumns_port_state_out_4_1_5 ), //o
    .port_state_out_4_1_6  (mixColumns_port_state_out_4_1_6 ), //o
    .port_state_out_4_1_7  (mixColumns_port_state_out_4_1_7 ), //o
    .port_state_out_4_2_0  (mixColumns_port_state_out_4_2_0 ), //o
    .port_state_out_4_2_1  (mixColumns_port_state_out_4_2_1 ), //o
    .port_state_out_4_2_2  (mixColumns_port_state_out_4_2_2 ), //o
    .port_state_out_4_2_3  (mixColumns_port_state_out_4_2_3 ), //o
    .port_state_out_4_2_4  (mixColumns_port_state_out_4_2_4 ), //o
    .port_state_out_4_2_5  (mixColumns_port_state_out_4_2_5 ), //o
    .port_state_out_4_2_6  (mixColumns_port_state_out_4_2_6 ), //o
    .port_state_out_4_2_7  (mixColumns_port_state_out_4_2_7 ), //o
    .port_state_out_4_3_0  (mixColumns_port_state_out_4_3_0 ), //o
    .port_state_out_4_3_1  (mixColumns_port_state_out_4_3_1 ), //o
    .port_state_out_4_3_2  (mixColumns_port_state_out_4_3_2 ), //o
    .port_state_out_4_3_3  (mixColumns_port_state_out_4_3_3 ), //o
    .port_state_out_4_3_4  (mixColumns_port_state_out_4_3_4 ), //o
    .port_state_out_4_3_5  (mixColumns_port_state_out_4_3_5 ), //o
    .port_state_out_4_3_6  (mixColumns_port_state_out_4_3_6 ), //o
    .port_state_out_4_3_7  (mixColumns_port_state_out_4_3_7 ), //o
    .port_state_out_5_0_0  (mixColumns_port_state_out_5_0_0 ), //o
    .port_state_out_5_0_1  (mixColumns_port_state_out_5_0_1 ), //o
    .port_state_out_5_0_2  (mixColumns_port_state_out_5_0_2 ), //o
    .port_state_out_5_0_3  (mixColumns_port_state_out_5_0_3 ), //o
    .port_state_out_5_0_4  (mixColumns_port_state_out_5_0_4 ), //o
    .port_state_out_5_0_5  (mixColumns_port_state_out_5_0_5 ), //o
    .port_state_out_5_0_6  (mixColumns_port_state_out_5_0_6 ), //o
    .port_state_out_5_0_7  (mixColumns_port_state_out_5_0_7 ), //o
    .port_state_out_5_1_0  (mixColumns_port_state_out_5_1_0 ), //o
    .port_state_out_5_1_1  (mixColumns_port_state_out_5_1_1 ), //o
    .port_state_out_5_1_2  (mixColumns_port_state_out_5_1_2 ), //o
    .port_state_out_5_1_3  (mixColumns_port_state_out_5_1_3 ), //o
    .port_state_out_5_1_4  (mixColumns_port_state_out_5_1_4 ), //o
    .port_state_out_5_1_5  (mixColumns_port_state_out_5_1_5 ), //o
    .port_state_out_5_1_6  (mixColumns_port_state_out_5_1_6 ), //o
    .port_state_out_5_1_7  (mixColumns_port_state_out_5_1_7 ), //o
    .port_state_out_5_2_0  (mixColumns_port_state_out_5_2_0 ), //o
    .port_state_out_5_2_1  (mixColumns_port_state_out_5_2_1 ), //o
    .port_state_out_5_2_2  (mixColumns_port_state_out_5_2_2 ), //o
    .port_state_out_5_2_3  (mixColumns_port_state_out_5_2_3 ), //o
    .port_state_out_5_2_4  (mixColumns_port_state_out_5_2_4 ), //o
    .port_state_out_5_2_5  (mixColumns_port_state_out_5_2_5 ), //o
    .port_state_out_5_2_6  (mixColumns_port_state_out_5_2_6 ), //o
    .port_state_out_5_2_7  (mixColumns_port_state_out_5_2_7 ), //o
    .port_state_out_5_3_0  (mixColumns_port_state_out_5_3_0 ), //o
    .port_state_out_5_3_1  (mixColumns_port_state_out_5_3_1 ), //o
    .port_state_out_5_3_2  (mixColumns_port_state_out_5_3_2 ), //o
    .port_state_out_5_3_3  (mixColumns_port_state_out_5_3_3 ), //o
    .port_state_out_5_3_4  (mixColumns_port_state_out_5_3_4 ), //o
    .port_state_out_5_3_5  (mixColumns_port_state_out_5_3_5 ), //o
    .port_state_out_5_3_6  (mixColumns_port_state_out_5_3_6 ), //o
    .port_state_out_5_3_7  (mixColumns_port_state_out_5_3_7 ), //o
    .port_state_out_6_0_0  (mixColumns_port_state_out_6_0_0 ), //o
    .port_state_out_6_0_1  (mixColumns_port_state_out_6_0_1 ), //o
    .port_state_out_6_0_2  (mixColumns_port_state_out_6_0_2 ), //o
    .port_state_out_6_0_3  (mixColumns_port_state_out_6_0_3 ), //o
    .port_state_out_6_0_4  (mixColumns_port_state_out_6_0_4 ), //o
    .port_state_out_6_0_5  (mixColumns_port_state_out_6_0_5 ), //o
    .port_state_out_6_0_6  (mixColumns_port_state_out_6_0_6 ), //o
    .port_state_out_6_0_7  (mixColumns_port_state_out_6_0_7 ), //o
    .port_state_out_6_1_0  (mixColumns_port_state_out_6_1_0 ), //o
    .port_state_out_6_1_1  (mixColumns_port_state_out_6_1_1 ), //o
    .port_state_out_6_1_2  (mixColumns_port_state_out_6_1_2 ), //o
    .port_state_out_6_1_3  (mixColumns_port_state_out_6_1_3 ), //o
    .port_state_out_6_1_4  (mixColumns_port_state_out_6_1_4 ), //o
    .port_state_out_6_1_5  (mixColumns_port_state_out_6_1_5 ), //o
    .port_state_out_6_1_6  (mixColumns_port_state_out_6_1_6 ), //o
    .port_state_out_6_1_7  (mixColumns_port_state_out_6_1_7 ), //o
    .port_state_out_6_2_0  (mixColumns_port_state_out_6_2_0 ), //o
    .port_state_out_6_2_1  (mixColumns_port_state_out_6_2_1 ), //o
    .port_state_out_6_2_2  (mixColumns_port_state_out_6_2_2 ), //o
    .port_state_out_6_2_3  (mixColumns_port_state_out_6_2_3 ), //o
    .port_state_out_6_2_4  (mixColumns_port_state_out_6_2_4 ), //o
    .port_state_out_6_2_5  (mixColumns_port_state_out_6_2_5 ), //o
    .port_state_out_6_2_6  (mixColumns_port_state_out_6_2_6 ), //o
    .port_state_out_6_2_7  (mixColumns_port_state_out_6_2_7 ), //o
    .port_state_out_6_3_0  (mixColumns_port_state_out_6_3_0 ), //o
    .port_state_out_6_3_1  (mixColumns_port_state_out_6_3_1 ), //o
    .port_state_out_6_3_2  (mixColumns_port_state_out_6_3_2 ), //o
    .port_state_out_6_3_3  (mixColumns_port_state_out_6_3_3 ), //o
    .port_state_out_6_3_4  (mixColumns_port_state_out_6_3_4 ), //o
    .port_state_out_6_3_5  (mixColumns_port_state_out_6_3_5 ), //o
    .port_state_out_6_3_6  (mixColumns_port_state_out_6_3_6 ), //o
    .port_state_out_6_3_7  (mixColumns_port_state_out_6_3_7 ), //o
    .port_state_out_7_0_0  (mixColumns_port_state_out_7_0_0 ), //o
    .port_state_out_7_0_1  (mixColumns_port_state_out_7_0_1 ), //o
    .port_state_out_7_0_2  (mixColumns_port_state_out_7_0_2 ), //o
    .port_state_out_7_0_3  (mixColumns_port_state_out_7_0_3 ), //o
    .port_state_out_7_0_4  (mixColumns_port_state_out_7_0_4 ), //o
    .port_state_out_7_0_5  (mixColumns_port_state_out_7_0_5 ), //o
    .port_state_out_7_0_6  (mixColumns_port_state_out_7_0_6 ), //o
    .port_state_out_7_0_7  (mixColumns_port_state_out_7_0_7 ), //o
    .port_state_out_7_1_0  (mixColumns_port_state_out_7_1_0 ), //o
    .port_state_out_7_1_1  (mixColumns_port_state_out_7_1_1 ), //o
    .port_state_out_7_1_2  (mixColumns_port_state_out_7_1_2 ), //o
    .port_state_out_7_1_3  (mixColumns_port_state_out_7_1_3 ), //o
    .port_state_out_7_1_4  (mixColumns_port_state_out_7_1_4 ), //o
    .port_state_out_7_1_5  (mixColumns_port_state_out_7_1_5 ), //o
    .port_state_out_7_1_6  (mixColumns_port_state_out_7_1_6 ), //o
    .port_state_out_7_1_7  (mixColumns_port_state_out_7_1_7 ), //o
    .port_state_out_7_2_0  (mixColumns_port_state_out_7_2_0 ), //o
    .port_state_out_7_2_1  (mixColumns_port_state_out_7_2_1 ), //o
    .port_state_out_7_2_2  (mixColumns_port_state_out_7_2_2 ), //o
    .port_state_out_7_2_3  (mixColumns_port_state_out_7_2_3 ), //o
    .port_state_out_7_2_4  (mixColumns_port_state_out_7_2_4 ), //o
    .port_state_out_7_2_5  (mixColumns_port_state_out_7_2_5 ), //o
    .port_state_out_7_2_6  (mixColumns_port_state_out_7_2_6 ), //o
    .port_state_out_7_2_7  (mixColumns_port_state_out_7_2_7 ), //o
    .port_state_out_7_3_0  (mixColumns_port_state_out_7_3_0 ), //o
    .port_state_out_7_3_1  (mixColumns_port_state_out_7_3_1 ), //o
    .port_state_out_7_3_2  (mixColumns_port_state_out_7_3_2 ), //o
    .port_state_out_7_3_3  (mixColumns_port_state_out_7_3_3 ), //o
    .port_state_out_7_3_4  (mixColumns_port_state_out_7_3_4 ), //o
    .port_state_out_7_3_5  (mixColumns_port_state_out_7_3_5 ), //o
    .port_state_out_7_3_6  (mixColumns_port_state_out_7_3_6 ), //o
    .port_state_out_7_3_7  (mixColumns_port_state_out_7_3_7 ), //o
    .port_state_out_8_0_0  (mixColumns_port_state_out_8_0_0 ), //o
    .port_state_out_8_0_1  (mixColumns_port_state_out_8_0_1 ), //o
    .port_state_out_8_0_2  (mixColumns_port_state_out_8_0_2 ), //o
    .port_state_out_8_0_3  (mixColumns_port_state_out_8_0_3 ), //o
    .port_state_out_8_0_4  (mixColumns_port_state_out_8_0_4 ), //o
    .port_state_out_8_0_5  (mixColumns_port_state_out_8_0_5 ), //o
    .port_state_out_8_0_6  (mixColumns_port_state_out_8_0_6 ), //o
    .port_state_out_8_0_7  (mixColumns_port_state_out_8_0_7 ), //o
    .port_state_out_8_1_0  (mixColumns_port_state_out_8_1_0 ), //o
    .port_state_out_8_1_1  (mixColumns_port_state_out_8_1_1 ), //o
    .port_state_out_8_1_2  (mixColumns_port_state_out_8_1_2 ), //o
    .port_state_out_8_1_3  (mixColumns_port_state_out_8_1_3 ), //o
    .port_state_out_8_1_4  (mixColumns_port_state_out_8_1_4 ), //o
    .port_state_out_8_1_5  (mixColumns_port_state_out_8_1_5 ), //o
    .port_state_out_8_1_6  (mixColumns_port_state_out_8_1_6 ), //o
    .port_state_out_8_1_7  (mixColumns_port_state_out_8_1_7 ), //o
    .port_state_out_8_2_0  (mixColumns_port_state_out_8_2_0 ), //o
    .port_state_out_8_2_1  (mixColumns_port_state_out_8_2_1 ), //o
    .port_state_out_8_2_2  (mixColumns_port_state_out_8_2_2 ), //o
    .port_state_out_8_2_3  (mixColumns_port_state_out_8_2_3 ), //o
    .port_state_out_8_2_4  (mixColumns_port_state_out_8_2_4 ), //o
    .port_state_out_8_2_5  (mixColumns_port_state_out_8_2_5 ), //o
    .port_state_out_8_2_6  (mixColumns_port_state_out_8_2_6 ), //o
    .port_state_out_8_2_7  (mixColumns_port_state_out_8_2_7 ), //o
    .port_state_out_8_3_0  (mixColumns_port_state_out_8_3_0 ), //o
    .port_state_out_8_3_1  (mixColumns_port_state_out_8_3_1 ), //o
    .port_state_out_8_3_2  (mixColumns_port_state_out_8_3_2 ), //o
    .port_state_out_8_3_3  (mixColumns_port_state_out_8_3_3 ), //o
    .port_state_out_8_3_4  (mixColumns_port_state_out_8_3_4 ), //o
    .port_state_out_8_3_5  (mixColumns_port_state_out_8_3_5 ), //o
    .port_state_out_8_3_6  (mixColumns_port_state_out_8_3_6 ), //o
    .port_state_out_8_3_7  (mixColumns_port_state_out_8_3_7 ), //o
    .port_state_out_9_0_0  (mixColumns_port_state_out_9_0_0 ), //o
    .port_state_out_9_0_1  (mixColumns_port_state_out_9_0_1 ), //o
    .port_state_out_9_0_2  (mixColumns_port_state_out_9_0_2 ), //o
    .port_state_out_9_0_3  (mixColumns_port_state_out_9_0_3 ), //o
    .port_state_out_9_0_4  (mixColumns_port_state_out_9_0_4 ), //o
    .port_state_out_9_0_5  (mixColumns_port_state_out_9_0_5 ), //o
    .port_state_out_9_0_6  (mixColumns_port_state_out_9_0_6 ), //o
    .port_state_out_9_0_7  (mixColumns_port_state_out_9_0_7 ), //o
    .port_state_out_9_1_0  (mixColumns_port_state_out_9_1_0 ), //o
    .port_state_out_9_1_1  (mixColumns_port_state_out_9_1_1 ), //o
    .port_state_out_9_1_2  (mixColumns_port_state_out_9_1_2 ), //o
    .port_state_out_9_1_3  (mixColumns_port_state_out_9_1_3 ), //o
    .port_state_out_9_1_4  (mixColumns_port_state_out_9_1_4 ), //o
    .port_state_out_9_1_5  (mixColumns_port_state_out_9_1_5 ), //o
    .port_state_out_9_1_6  (mixColumns_port_state_out_9_1_6 ), //o
    .port_state_out_9_1_7  (mixColumns_port_state_out_9_1_7 ), //o
    .port_state_out_9_2_0  (mixColumns_port_state_out_9_2_0 ), //o
    .port_state_out_9_2_1  (mixColumns_port_state_out_9_2_1 ), //o
    .port_state_out_9_2_2  (mixColumns_port_state_out_9_2_2 ), //o
    .port_state_out_9_2_3  (mixColumns_port_state_out_9_2_3 ), //o
    .port_state_out_9_2_4  (mixColumns_port_state_out_9_2_4 ), //o
    .port_state_out_9_2_5  (mixColumns_port_state_out_9_2_5 ), //o
    .port_state_out_9_2_6  (mixColumns_port_state_out_9_2_6 ), //o
    .port_state_out_9_2_7  (mixColumns_port_state_out_9_2_7 ), //o
    .port_state_out_9_3_0  (mixColumns_port_state_out_9_3_0 ), //o
    .port_state_out_9_3_1  (mixColumns_port_state_out_9_3_1 ), //o
    .port_state_out_9_3_2  (mixColumns_port_state_out_9_3_2 ), //o
    .port_state_out_9_3_3  (mixColumns_port_state_out_9_3_3 ), //o
    .port_state_out_9_3_4  (mixColumns_port_state_out_9_3_4 ), //o
    .port_state_out_9_3_5  (mixColumns_port_state_out_9_3_5 ), //o
    .port_state_out_9_3_6  (mixColumns_port_state_out_9_3_6 ), //o
    .port_state_out_9_3_7  (mixColumns_port_state_out_9_3_7 ), //o
    .port_state_out_10_0_0 (mixColumns_port_state_out_10_0_0), //o
    .port_state_out_10_0_1 (mixColumns_port_state_out_10_0_1), //o
    .port_state_out_10_0_2 (mixColumns_port_state_out_10_0_2), //o
    .port_state_out_10_0_3 (mixColumns_port_state_out_10_0_3), //o
    .port_state_out_10_0_4 (mixColumns_port_state_out_10_0_4), //o
    .port_state_out_10_0_5 (mixColumns_port_state_out_10_0_5), //o
    .port_state_out_10_0_6 (mixColumns_port_state_out_10_0_6), //o
    .port_state_out_10_0_7 (mixColumns_port_state_out_10_0_7), //o
    .port_state_out_10_1_0 (mixColumns_port_state_out_10_1_0), //o
    .port_state_out_10_1_1 (mixColumns_port_state_out_10_1_1), //o
    .port_state_out_10_1_2 (mixColumns_port_state_out_10_1_2), //o
    .port_state_out_10_1_3 (mixColumns_port_state_out_10_1_3), //o
    .port_state_out_10_1_4 (mixColumns_port_state_out_10_1_4), //o
    .port_state_out_10_1_5 (mixColumns_port_state_out_10_1_5), //o
    .port_state_out_10_1_6 (mixColumns_port_state_out_10_1_6), //o
    .port_state_out_10_1_7 (mixColumns_port_state_out_10_1_7), //o
    .port_state_out_10_2_0 (mixColumns_port_state_out_10_2_0), //o
    .port_state_out_10_2_1 (mixColumns_port_state_out_10_2_1), //o
    .port_state_out_10_2_2 (mixColumns_port_state_out_10_2_2), //o
    .port_state_out_10_2_3 (mixColumns_port_state_out_10_2_3), //o
    .port_state_out_10_2_4 (mixColumns_port_state_out_10_2_4), //o
    .port_state_out_10_2_5 (mixColumns_port_state_out_10_2_5), //o
    .port_state_out_10_2_6 (mixColumns_port_state_out_10_2_6), //o
    .port_state_out_10_2_7 (mixColumns_port_state_out_10_2_7), //o
    .port_state_out_10_3_0 (mixColumns_port_state_out_10_3_0), //o
    .port_state_out_10_3_1 (mixColumns_port_state_out_10_3_1), //o
    .port_state_out_10_3_2 (mixColumns_port_state_out_10_3_2), //o
    .port_state_out_10_3_3 (mixColumns_port_state_out_10_3_3), //o
    .port_state_out_10_3_4 (mixColumns_port_state_out_10_3_4), //o
    .port_state_out_10_3_5 (mixColumns_port_state_out_10_3_5), //o
    .port_state_out_10_3_6 (mixColumns_port_state_out_10_3_6), //o
    .port_state_out_10_3_7 (mixColumns_port_state_out_10_3_7), //o
    .port_state_out_11_0_0 (mixColumns_port_state_out_11_0_0), //o
    .port_state_out_11_0_1 (mixColumns_port_state_out_11_0_1), //o
    .port_state_out_11_0_2 (mixColumns_port_state_out_11_0_2), //o
    .port_state_out_11_0_3 (mixColumns_port_state_out_11_0_3), //o
    .port_state_out_11_0_4 (mixColumns_port_state_out_11_0_4), //o
    .port_state_out_11_0_5 (mixColumns_port_state_out_11_0_5), //o
    .port_state_out_11_0_6 (mixColumns_port_state_out_11_0_6), //o
    .port_state_out_11_0_7 (mixColumns_port_state_out_11_0_7), //o
    .port_state_out_11_1_0 (mixColumns_port_state_out_11_1_0), //o
    .port_state_out_11_1_1 (mixColumns_port_state_out_11_1_1), //o
    .port_state_out_11_1_2 (mixColumns_port_state_out_11_1_2), //o
    .port_state_out_11_1_3 (mixColumns_port_state_out_11_1_3), //o
    .port_state_out_11_1_4 (mixColumns_port_state_out_11_1_4), //o
    .port_state_out_11_1_5 (mixColumns_port_state_out_11_1_5), //o
    .port_state_out_11_1_6 (mixColumns_port_state_out_11_1_6), //o
    .port_state_out_11_1_7 (mixColumns_port_state_out_11_1_7), //o
    .port_state_out_11_2_0 (mixColumns_port_state_out_11_2_0), //o
    .port_state_out_11_2_1 (mixColumns_port_state_out_11_2_1), //o
    .port_state_out_11_2_2 (mixColumns_port_state_out_11_2_2), //o
    .port_state_out_11_2_3 (mixColumns_port_state_out_11_2_3), //o
    .port_state_out_11_2_4 (mixColumns_port_state_out_11_2_4), //o
    .port_state_out_11_2_5 (mixColumns_port_state_out_11_2_5), //o
    .port_state_out_11_2_6 (mixColumns_port_state_out_11_2_6), //o
    .port_state_out_11_2_7 (mixColumns_port_state_out_11_2_7), //o
    .port_state_out_11_3_0 (mixColumns_port_state_out_11_3_0), //o
    .port_state_out_11_3_1 (mixColumns_port_state_out_11_3_1), //o
    .port_state_out_11_3_2 (mixColumns_port_state_out_11_3_2), //o
    .port_state_out_11_3_3 (mixColumns_port_state_out_11_3_3), //o
    .port_state_out_11_3_4 (mixColumns_port_state_out_11_3_4), //o
    .port_state_out_11_3_5 (mixColumns_port_state_out_11_3_5), //o
    .port_state_out_11_3_6 (mixColumns_port_state_out_11_3_6), //o
    .port_state_out_11_3_7 (mixColumns_port_state_out_11_3_7), //o
    .port_state_out_12_0_0 (mixColumns_port_state_out_12_0_0), //o
    .port_state_out_12_0_1 (mixColumns_port_state_out_12_0_1), //o
    .port_state_out_12_0_2 (mixColumns_port_state_out_12_0_2), //o
    .port_state_out_12_0_3 (mixColumns_port_state_out_12_0_3), //o
    .port_state_out_12_0_4 (mixColumns_port_state_out_12_0_4), //o
    .port_state_out_12_0_5 (mixColumns_port_state_out_12_0_5), //o
    .port_state_out_12_0_6 (mixColumns_port_state_out_12_0_6), //o
    .port_state_out_12_0_7 (mixColumns_port_state_out_12_0_7), //o
    .port_state_out_12_1_0 (mixColumns_port_state_out_12_1_0), //o
    .port_state_out_12_1_1 (mixColumns_port_state_out_12_1_1), //o
    .port_state_out_12_1_2 (mixColumns_port_state_out_12_1_2), //o
    .port_state_out_12_1_3 (mixColumns_port_state_out_12_1_3), //o
    .port_state_out_12_1_4 (mixColumns_port_state_out_12_1_4), //o
    .port_state_out_12_1_5 (mixColumns_port_state_out_12_1_5), //o
    .port_state_out_12_1_6 (mixColumns_port_state_out_12_1_6), //o
    .port_state_out_12_1_7 (mixColumns_port_state_out_12_1_7), //o
    .port_state_out_12_2_0 (mixColumns_port_state_out_12_2_0), //o
    .port_state_out_12_2_1 (mixColumns_port_state_out_12_2_1), //o
    .port_state_out_12_2_2 (mixColumns_port_state_out_12_2_2), //o
    .port_state_out_12_2_3 (mixColumns_port_state_out_12_2_3), //o
    .port_state_out_12_2_4 (mixColumns_port_state_out_12_2_4), //o
    .port_state_out_12_2_5 (mixColumns_port_state_out_12_2_5), //o
    .port_state_out_12_2_6 (mixColumns_port_state_out_12_2_6), //o
    .port_state_out_12_2_7 (mixColumns_port_state_out_12_2_7), //o
    .port_state_out_12_3_0 (mixColumns_port_state_out_12_3_0), //o
    .port_state_out_12_3_1 (mixColumns_port_state_out_12_3_1), //o
    .port_state_out_12_3_2 (mixColumns_port_state_out_12_3_2), //o
    .port_state_out_12_3_3 (mixColumns_port_state_out_12_3_3), //o
    .port_state_out_12_3_4 (mixColumns_port_state_out_12_3_4), //o
    .port_state_out_12_3_5 (mixColumns_port_state_out_12_3_5), //o
    .port_state_out_12_3_6 (mixColumns_port_state_out_12_3_6), //o
    .port_state_out_12_3_7 (mixColumns_port_state_out_12_3_7), //o
    .port_state_out_13_0_0 (mixColumns_port_state_out_13_0_0), //o
    .port_state_out_13_0_1 (mixColumns_port_state_out_13_0_1), //o
    .port_state_out_13_0_2 (mixColumns_port_state_out_13_0_2), //o
    .port_state_out_13_0_3 (mixColumns_port_state_out_13_0_3), //o
    .port_state_out_13_0_4 (mixColumns_port_state_out_13_0_4), //o
    .port_state_out_13_0_5 (mixColumns_port_state_out_13_0_5), //o
    .port_state_out_13_0_6 (mixColumns_port_state_out_13_0_6), //o
    .port_state_out_13_0_7 (mixColumns_port_state_out_13_0_7), //o
    .port_state_out_13_1_0 (mixColumns_port_state_out_13_1_0), //o
    .port_state_out_13_1_1 (mixColumns_port_state_out_13_1_1), //o
    .port_state_out_13_1_2 (mixColumns_port_state_out_13_1_2), //o
    .port_state_out_13_1_3 (mixColumns_port_state_out_13_1_3), //o
    .port_state_out_13_1_4 (mixColumns_port_state_out_13_1_4), //o
    .port_state_out_13_1_5 (mixColumns_port_state_out_13_1_5), //o
    .port_state_out_13_1_6 (mixColumns_port_state_out_13_1_6), //o
    .port_state_out_13_1_7 (mixColumns_port_state_out_13_1_7), //o
    .port_state_out_13_2_0 (mixColumns_port_state_out_13_2_0), //o
    .port_state_out_13_2_1 (mixColumns_port_state_out_13_2_1), //o
    .port_state_out_13_2_2 (mixColumns_port_state_out_13_2_2), //o
    .port_state_out_13_2_3 (mixColumns_port_state_out_13_2_3), //o
    .port_state_out_13_2_4 (mixColumns_port_state_out_13_2_4), //o
    .port_state_out_13_2_5 (mixColumns_port_state_out_13_2_5), //o
    .port_state_out_13_2_6 (mixColumns_port_state_out_13_2_6), //o
    .port_state_out_13_2_7 (mixColumns_port_state_out_13_2_7), //o
    .port_state_out_13_3_0 (mixColumns_port_state_out_13_3_0), //o
    .port_state_out_13_3_1 (mixColumns_port_state_out_13_3_1), //o
    .port_state_out_13_3_2 (mixColumns_port_state_out_13_3_2), //o
    .port_state_out_13_3_3 (mixColumns_port_state_out_13_3_3), //o
    .port_state_out_13_3_4 (mixColumns_port_state_out_13_3_4), //o
    .port_state_out_13_3_5 (mixColumns_port_state_out_13_3_5), //o
    .port_state_out_13_3_6 (mixColumns_port_state_out_13_3_6), //o
    .port_state_out_13_3_7 (mixColumns_port_state_out_13_3_7), //o
    .port_state_out_14_0_0 (mixColumns_port_state_out_14_0_0), //o
    .port_state_out_14_0_1 (mixColumns_port_state_out_14_0_1), //o
    .port_state_out_14_0_2 (mixColumns_port_state_out_14_0_2), //o
    .port_state_out_14_0_3 (mixColumns_port_state_out_14_0_3), //o
    .port_state_out_14_0_4 (mixColumns_port_state_out_14_0_4), //o
    .port_state_out_14_0_5 (mixColumns_port_state_out_14_0_5), //o
    .port_state_out_14_0_6 (mixColumns_port_state_out_14_0_6), //o
    .port_state_out_14_0_7 (mixColumns_port_state_out_14_0_7), //o
    .port_state_out_14_1_0 (mixColumns_port_state_out_14_1_0), //o
    .port_state_out_14_1_1 (mixColumns_port_state_out_14_1_1), //o
    .port_state_out_14_1_2 (mixColumns_port_state_out_14_1_2), //o
    .port_state_out_14_1_3 (mixColumns_port_state_out_14_1_3), //o
    .port_state_out_14_1_4 (mixColumns_port_state_out_14_1_4), //o
    .port_state_out_14_1_5 (mixColumns_port_state_out_14_1_5), //o
    .port_state_out_14_1_6 (mixColumns_port_state_out_14_1_6), //o
    .port_state_out_14_1_7 (mixColumns_port_state_out_14_1_7), //o
    .port_state_out_14_2_0 (mixColumns_port_state_out_14_2_0), //o
    .port_state_out_14_2_1 (mixColumns_port_state_out_14_2_1), //o
    .port_state_out_14_2_2 (mixColumns_port_state_out_14_2_2), //o
    .port_state_out_14_2_3 (mixColumns_port_state_out_14_2_3), //o
    .port_state_out_14_2_4 (mixColumns_port_state_out_14_2_4), //o
    .port_state_out_14_2_5 (mixColumns_port_state_out_14_2_5), //o
    .port_state_out_14_2_6 (mixColumns_port_state_out_14_2_6), //o
    .port_state_out_14_2_7 (mixColumns_port_state_out_14_2_7), //o
    .port_state_out_14_3_0 (mixColumns_port_state_out_14_3_0), //o
    .port_state_out_14_3_1 (mixColumns_port_state_out_14_3_1), //o
    .port_state_out_14_3_2 (mixColumns_port_state_out_14_3_2), //o
    .port_state_out_14_3_3 (mixColumns_port_state_out_14_3_3), //o
    .port_state_out_14_3_4 (mixColumns_port_state_out_14_3_4), //o
    .port_state_out_14_3_5 (mixColumns_port_state_out_14_3_5), //o
    .port_state_out_14_3_6 (mixColumns_port_state_out_14_3_6), //o
    .port_state_out_14_3_7 (mixColumns_port_state_out_14_3_7), //o
    .port_state_out_15_0_0 (mixColumns_port_state_out_15_0_0), //o
    .port_state_out_15_0_1 (mixColumns_port_state_out_15_0_1), //o
    .port_state_out_15_0_2 (mixColumns_port_state_out_15_0_2), //o
    .port_state_out_15_0_3 (mixColumns_port_state_out_15_0_3), //o
    .port_state_out_15_0_4 (mixColumns_port_state_out_15_0_4), //o
    .port_state_out_15_0_5 (mixColumns_port_state_out_15_0_5), //o
    .port_state_out_15_0_6 (mixColumns_port_state_out_15_0_6), //o
    .port_state_out_15_0_7 (mixColumns_port_state_out_15_0_7), //o
    .port_state_out_15_1_0 (mixColumns_port_state_out_15_1_0), //o
    .port_state_out_15_1_1 (mixColumns_port_state_out_15_1_1), //o
    .port_state_out_15_1_2 (mixColumns_port_state_out_15_1_2), //o
    .port_state_out_15_1_3 (mixColumns_port_state_out_15_1_3), //o
    .port_state_out_15_1_4 (mixColumns_port_state_out_15_1_4), //o
    .port_state_out_15_1_5 (mixColumns_port_state_out_15_1_5), //o
    .port_state_out_15_1_6 (mixColumns_port_state_out_15_1_6), //o
    .port_state_out_15_1_7 (mixColumns_port_state_out_15_1_7), //o
    .port_state_out_15_2_0 (mixColumns_port_state_out_15_2_0), //o
    .port_state_out_15_2_1 (mixColumns_port_state_out_15_2_1), //o
    .port_state_out_15_2_2 (mixColumns_port_state_out_15_2_2), //o
    .port_state_out_15_2_3 (mixColumns_port_state_out_15_2_3), //o
    .port_state_out_15_2_4 (mixColumns_port_state_out_15_2_4), //o
    .port_state_out_15_2_5 (mixColumns_port_state_out_15_2_5), //o
    .port_state_out_15_2_6 (mixColumns_port_state_out_15_2_6), //o
    .port_state_out_15_2_7 (mixColumns_port_state_out_15_2_7), //o
    .port_state_out_15_3_0 (mixColumns_port_state_out_15_3_0), //o
    .port_state_out_15_3_1 (mixColumns_port_state_out_15_3_1), //o
    .port_state_out_15_3_2 (mixColumns_port_state_out_15_3_2), //o
    .port_state_out_15_3_3 (mixColumns_port_state_out_15_3_3), //o
    .port_state_out_15_3_4 (mixColumns_port_state_out_15_3_4), //o
    .port_state_out_15_3_5 (mixColumns_port_state_out_15_3_5), //o
    .port_state_out_15_3_6 (mixColumns_port_state_out_15_3_6), //o
    .port_state_out_15_3_7 (mixColumns_port_state_out_15_3_7)  //o
  );
  assign subBytes_out_0_0_0 = sbox_AES_BoyarPeralta_16_port_o_0_0;
  assign subBytes_out_0_0_1 = sbox_AES_BoyarPeralta_16_port_o_0_1;
  assign subBytes_out_0_0_2 = sbox_AES_BoyarPeralta_16_port_o_0_2;
  assign subBytes_out_0_0_3 = sbox_AES_BoyarPeralta_16_port_o_0_3;
  assign subBytes_out_0_0_4 = sbox_AES_BoyarPeralta_16_port_o_0_4;
  assign subBytes_out_0_0_5 = sbox_AES_BoyarPeralta_16_port_o_0_5;
  assign subBytes_out_0_0_6 = sbox_AES_BoyarPeralta_16_port_o_0_6;
  assign subBytes_out_0_0_7 = sbox_AES_BoyarPeralta_16_port_o_0_7;
  assign subBytes_out_0_1_0 = sbox_AES_BoyarPeralta_16_port_o_1_0;
  assign subBytes_out_0_1_1 = sbox_AES_BoyarPeralta_16_port_o_1_1;
  assign subBytes_out_0_1_2 = sbox_AES_BoyarPeralta_16_port_o_1_2;
  assign subBytes_out_0_1_3 = sbox_AES_BoyarPeralta_16_port_o_1_3;
  assign subBytes_out_0_1_4 = sbox_AES_BoyarPeralta_16_port_o_1_4;
  assign subBytes_out_0_1_5 = sbox_AES_BoyarPeralta_16_port_o_1_5;
  assign subBytes_out_0_1_6 = sbox_AES_BoyarPeralta_16_port_o_1_6;
  assign subBytes_out_0_1_7 = sbox_AES_BoyarPeralta_16_port_o_1_7;
  assign subBytes_out_0_2_0 = sbox_AES_BoyarPeralta_16_port_o_2_0;
  assign subBytes_out_0_2_1 = sbox_AES_BoyarPeralta_16_port_o_2_1;
  assign subBytes_out_0_2_2 = sbox_AES_BoyarPeralta_16_port_o_2_2;
  assign subBytes_out_0_2_3 = sbox_AES_BoyarPeralta_16_port_o_2_3;
  assign subBytes_out_0_2_4 = sbox_AES_BoyarPeralta_16_port_o_2_4;
  assign subBytes_out_0_2_5 = sbox_AES_BoyarPeralta_16_port_o_2_5;
  assign subBytes_out_0_2_6 = sbox_AES_BoyarPeralta_16_port_o_2_6;
  assign subBytes_out_0_2_7 = sbox_AES_BoyarPeralta_16_port_o_2_7;
  assign subBytes_out_0_3_0 = sbox_AES_BoyarPeralta_16_port_o_3_0;
  assign subBytes_out_0_3_1 = sbox_AES_BoyarPeralta_16_port_o_3_1;
  assign subBytes_out_0_3_2 = sbox_AES_BoyarPeralta_16_port_o_3_2;
  assign subBytes_out_0_3_3 = sbox_AES_BoyarPeralta_16_port_o_3_3;
  assign subBytes_out_0_3_4 = sbox_AES_BoyarPeralta_16_port_o_3_4;
  assign subBytes_out_0_3_5 = sbox_AES_BoyarPeralta_16_port_o_3_5;
  assign subBytes_out_0_3_6 = sbox_AES_BoyarPeralta_16_port_o_3_6;
  assign subBytes_out_0_3_7 = sbox_AES_BoyarPeralta_16_port_o_3_7;
  assign subBytes_out_1_0_0 = sbox_AES_BoyarPeralta_17_port_o_0_0;
  assign subBytes_out_1_0_1 = sbox_AES_BoyarPeralta_17_port_o_0_1;
  assign subBytes_out_1_0_2 = sbox_AES_BoyarPeralta_17_port_o_0_2;
  assign subBytes_out_1_0_3 = sbox_AES_BoyarPeralta_17_port_o_0_3;
  assign subBytes_out_1_0_4 = sbox_AES_BoyarPeralta_17_port_o_0_4;
  assign subBytes_out_1_0_5 = sbox_AES_BoyarPeralta_17_port_o_0_5;
  assign subBytes_out_1_0_6 = sbox_AES_BoyarPeralta_17_port_o_0_6;
  assign subBytes_out_1_0_7 = sbox_AES_BoyarPeralta_17_port_o_0_7;
  assign subBytes_out_1_1_0 = sbox_AES_BoyarPeralta_17_port_o_1_0;
  assign subBytes_out_1_1_1 = sbox_AES_BoyarPeralta_17_port_o_1_1;
  assign subBytes_out_1_1_2 = sbox_AES_BoyarPeralta_17_port_o_1_2;
  assign subBytes_out_1_1_3 = sbox_AES_BoyarPeralta_17_port_o_1_3;
  assign subBytes_out_1_1_4 = sbox_AES_BoyarPeralta_17_port_o_1_4;
  assign subBytes_out_1_1_5 = sbox_AES_BoyarPeralta_17_port_o_1_5;
  assign subBytes_out_1_1_6 = sbox_AES_BoyarPeralta_17_port_o_1_6;
  assign subBytes_out_1_1_7 = sbox_AES_BoyarPeralta_17_port_o_1_7;
  assign subBytes_out_1_2_0 = sbox_AES_BoyarPeralta_17_port_o_2_0;
  assign subBytes_out_1_2_1 = sbox_AES_BoyarPeralta_17_port_o_2_1;
  assign subBytes_out_1_2_2 = sbox_AES_BoyarPeralta_17_port_o_2_2;
  assign subBytes_out_1_2_3 = sbox_AES_BoyarPeralta_17_port_o_2_3;
  assign subBytes_out_1_2_4 = sbox_AES_BoyarPeralta_17_port_o_2_4;
  assign subBytes_out_1_2_5 = sbox_AES_BoyarPeralta_17_port_o_2_5;
  assign subBytes_out_1_2_6 = sbox_AES_BoyarPeralta_17_port_o_2_6;
  assign subBytes_out_1_2_7 = sbox_AES_BoyarPeralta_17_port_o_2_7;
  assign subBytes_out_1_3_0 = sbox_AES_BoyarPeralta_17_port_o_3_0;
  assign subBytes_out_1_3_1 = sbox_AES_BoyarPeralta_17_port_o_3_1;
  assign subBytes_out_1_3_2 = sbox_AES_BoyarPeralta_17_port_o_3_2;
  assign subBytes_out_1_3_3 = sbox_AES_BoyarPeralta_17_port_o_3_3;
  assign subBytes_out_1_3_4 = sbox_AES_BoyarPeralta_17_port_o_3_4;
  assign subBytes_out_1_3_5 = sbox_AES_BoyarPeralta_17_port_o_3_5;
  assign subBytes_out_1_3_6 = sbox_AES_BoyarPeralta_17_port_o_3_6;
  assign subBytes_out_1_3_7 = sbox_AES_BoyarPeralta_17_port_o_3_7;
  assign subBytes_out_2_0_0 = sbox_AES_BoyarPeralta_18_port_o_0_0;
  assign subBytes_out_2_0_1 = sbox_AES_BoyarPeralta_18_port_o_0_1;
  assign subBytes_out_2_0_2 = sbox_AES_BoyarPeralta_18_port_o_0_2;
  assign subBytes_out_2_0_3 = sbox_AES_BoyarPeralta_18_port_o_0_3;
  assign subBytes_out_2_0_4 = sbox_AES_BoyarPeralta_18_port_o_0_4;
  assign subBytes_out_2_0_5 = sbox_AES_BoyarPeralta_18_port_o_0_5;
  assign subBytes_out_2_0_6 = sbox_AES_BoyarPeralta_18_port_o_0_6;
  assign subBytes_out_2_0_7 = sbox_AES_BoyarPeralta_18_port_o_0_7;
  assign subBytes_out_2_1_0 = sbox_AES_BoyarPeralta_18_port_o_1_0;
  assign subBytes_out_2_1_1 = sbox_AES_BoyarPeralta_18_port_o_1_1;
  assign subBytes_out_2_1_2 = sbox_AES_BoyarPeralta_18_port_o_1_2;
  assign subBytes_out_2_1_3 = sbox_AES_BoyarPeralta_18_port_o_1_3;
  assign subBytes_out_2_1_4 = sbox_AES_BoyarPeralta_18_port_o_1_4;
  assign subBytes_out_2_1_5 = sbox_AES_BoyarPeralta_18_port_o_1_5;
  assign subBytes_out_2_1_6 = sbox_AES_BoyarPeralta_18_port_o_1_6;
  assign subBytes_out_2_1_7 = sbox_AES_BoyarPeralta_18_port_o_1_7;
  assign subBytes_out_2_2_0 = sbox_AES_BoyarPeralta_18_port_o_2_0;
  assign subBytes_out_2_2_1 = sbox_AES_BoyarPeralta_18_port_o_2_1;
  assign subBytes_out_2_2_2 = sbox_AES_BoyarPeralta_18_port_o_2_2;
  assign subBytes_out_2_2_3 = sbox_AES_BoyarPeralta_18_port_o_2_3;
  assign subBytes_out_2_2_4 = sbox_AES_BoyarPeralta_18_port_o_2_4;
  assign subBytes_out_2_2_5 = sbox_AES_BoyarPeralta_18_port_o_2_5;
  assign subBytes_out_2_2_6 = sbox_AES_BoyarPeralta_18_port_o_2_6;
  assign subBytes_out_2_2_7 = sbox_AES_BoyarPeralta_18_port_o_2_7;
  assign subBytes_out_2_3_0 = sbox_AES_BoyarPeralta_18_port_o_3_0;
  assign subBytes_out_2_3_1 = sbox_AES_BoyarPeralta_18_port_o_3_1;
  assign subBytes_out_2_3_2 = sbox_AES_BoyarPeralta_18_port_o_3_2;
  assign subBytes_out_2_3_3 = sbox_AES_BoyarPeralta_18_port_o_3_3;
  assign subBytes_out_2_3_4 = sbox_AES_BoyarPeralta_18_port_o_3_4;
  assign subBytes_out_2_3_5 = sbox_AES_BoyarPeralta_18_port_o_3_5;
  assign subBytes_out_2_3_6 = sbox_AES_BoyarPeralta_18_port_o_3_6;
  assign subBytes_out_2_3_7 = sbox_AES_BoyarPeralta_18_port_o_3_7;
  assign subBytes_out_3_0_0 = sbox_AES_BoyarPeralta_19_port_o_0_0;
  assign subBytes_out_3_0_1 = sbox_AES_BoyarPeralta_19_port_o_0_1;
  assign subBytes_out_3_0_2 = sbox_AES_BoyarPeralta_19_port_o_0_2;
  assign subBytes_out_3_0_3 = sbox_AES_BoyarPeralta_19_port_o_0_3;
  assign subBytes_out_3_0_4 = sbox_AES_BoyarPeralta_19_port_o_0_4;
  assign subBytes_out_3_0_5 = sbox_AES_BoyarPeralta_19_port_o_0_5;
  assign subBytes_out_3_0_6 = sbox_AES_BoyarPeralta_19_port_o_0_6;
  assign subBytes_out_3_0_7 = sbox_AES_BoyarPeralta_19_port_o_0_7;
  assign subBytes_out_3_1_0 = sbox_AES_BoyarPeralta_19_port_o_1_0;
  assign subBytes_out_3_1_1 = sbox_AES_BoyarPeralta_19_port_o_1_1;
  assign subBytes_out_3_1_2 = sbox_AES_BoyarPeralta_19_port_o_1_2;
  assign subBytes_out_3_1_3 = sbox_AES_BoyarPeralta_19_port_o_1_3;
  assign subBytes_out_3_1_4 = sbox_AES_BoyarPeralta_19_port_o_1_4;
  assign subBytes_out_3_1_5 = sbox_AES_BoyarPeralta_19_port_o_1_5;
  assign subBytes_out_3_1_6 = sbox_AES_BoyarPeralta_19_port_o_1_6;
  assign subBytes_out_3_1_7 = sbox_AES_BoyarPeralta_19_port_o_1_7;
  assign subBytes_out_3_2_0 = sbox_AES_BoyarPeralta_19_port_o_2_0;
  assign subBytes_out_3_2_1 = sbox_AES_BoyarPeralta_19_port_o_2_1;
  assign subBytes_out_3_2_2 = sbox_AES_BoyarPeralta_19_port_o_2_2;
  assign subBytes_out_3_2_3 = sbox_AES_BoyarPeralta_19_port_o_2_3;
  assign subBytes_out_3_2_4 = sbox_AES_BoyarPeralta_19_port_o_2_4;
  assign subBytes_out_3_2_5 = sbox_AES_BoyarPeralta_19_port_o_2_5;
  assign subBytes_out_3_2_6 = sbox_AES_BoyarPeralta_19_port_o_2_6;
  assign subBytes_out_3_2_7 = sbox_AES_BoyarPeralta_19_port_o_2_7;
  assign subBytes_out_3_3_0 = sbox_AES_BoyarPeralta_19_port_o_3_0;
  assign subBytes_out_3_3_1 = sbox_AES_BoyarPeralta_19_port_o_3_1;
  assign subBytes_out_3_3_2 = sbox_AES_BoyarPeralta_19_port_o_3_2;
  assign subBytes_out_3_3_3 = sbox_AES_BoyarPeralta_19_port_o_3_3;
  assign subBytes_out_3_3_4 = sbox_AES_BoyarPeralta_19_port_o_3_4;
  assign subBytes_out_3_3_5 = sbox_AES_BoyarPeralta_19_port_o_3_5;
  assign subBytes_out_3_3_6 = sbox_AES_BoyarPeralta_19_port_o_3_6;
  assign subBytes_out_3_3_7 = sbox_AES_BoyarPeralta_19_port_o_3_7;
  assign subBytes_out_4_0_0 = sbox_AES_BoyarPeralta_20_port_o_0_0;
  assign subBytes_out_4_0_1 = sbox_AES_BoyarPeralta_20_port_o_0_1;
  assign subBytes_out_4_0_2 = sbox_AES_BoyarPeralta_20_port_o_0_2;
  assign subBytes_out_4_0_3 = sbox_AES_BoyarPeralta_20_port_o_0_3;
  assign subBytes_out_4_0_4 = sbox_AES_BoyarPeralta_20_port_o_0_4;
  assign subBytes_out_4_0_5 = sbox_AES_BoyarPeralta_20_port_o_0_5;
  assign subBytes_out_4_0_6 = sbox_AES_BoyarPeralta_20_port_o_0_6;
  assign subBytes_out_4_0_7 = sbox_AES_BoyarPeralta_20_port_o_0_7;
  assign subBytes_out_4_1_0 = sbox_AES_BoyarPeralta_20_port_o_1_0;
  assign subBytes_out_4_1_1 = sbox_AES_BoyarPeralta_20_port_o_1_1;
  assign subBytes_out_4_1_2 = sbox_AES_BoyarPeralta_20_port_o_1_2;
  assign subBytes_out_4_1_3 = sbox_AES_BoyarPeralta_20_port_o_1_3;
  assign subBytes_out_4_1_4 = sbox_AES_BoyarPeralta_20_port_o_1_4;
  assign subBytes_out_4_1_5 = sbox_AES_BoyarPeralta_20_port_o_1_5;
  assign subBytes_out_4_1_6 = sbox_AES_BoyarPeralta_20_port_o_1_6;
  assign subBytes_out_4_1_7 = sbox_AES_BoyarPeralta_20_port_o_1_7;
  assign subBytes_out_4_2_0 = sbox_AES_BoyarPeralta_20_port_o_2_0;
  assign subBytes_out_4_2_1 = sbox_AES_BoyarPeralta_20_port_o_2_1;
  assign subBytes_out_4_2_2 = sbox_AES_BoyarPeralta_20_port_o_2_2;
  assign subBytes_out_4_2_3 = sbox_AES_BoyarPeralta_20_port_o_2_3;
  assign subBytes_out_4_2_4 = sbox_AES_BoyarPeralta_20_port_o_2_4;
  assign subBytes_out_4_2_5 = sbox_AES_BoyarPeralta_20_port_o_2_5;
  assign subBytes_out_4_2_6 = sbox_AES_BoyarPeralta_20_port_o_2_6;
  assign subBytes_out_4_2_7 = sbox_AES_BoyarPeralta_20_port_o_2_7;
  assign subBytes_out_4_3_0 = sbox_AES_BoyarPeralta_20_port_o_3_0;
  assign subBytes_out_4_3_1 = sbox_AES_BoyarPeralta_20_port_o_3_1;
  assign subBytes_out_4_3_2 = sbox_AES_BoyarPeralta_20_port_o_3_2;
  assign subBytes_out_4_3_3 = sbox_AES_BoyarPeralta_20_port_o_3_3;
  assign subBytes_out_4_3_4 = sbox_AES_BoyarPeralta_20_port_o_3_4;
  assign subBytes_out_4_3_5 = sbox_AES_BoyarPeralta_20_port_o_3_5;
  assign subBytes_out_4_3_6 = sbox_AES_BoyarPeralta_20_port_o_3_6;
  assign subBytes_out_4_3_7 = sbox_AES_BoyarPeralta_20_port_o_3_7;
  assign subBytes_out_5_0_0 = sbox_AES_BoyarPeralta_21_port_o_0_0;
  assign subBytes_out_5_0_1 = sbox_AES_BoyarPeralta_21_port_o_0_1;
  assign subBytes_out_5_0_2 = sbox_AES_BoyarPeralta_21_port_o_0_2;
  assign subBytes_out_5_0_3 = sbox_AES_BoyarPeralta_21_port_o_0_3;
  assign subBytes_out_5_0_4 = sbox_AES_BoyarPeralta_21_port_o_0_4;
  assign subBytes_out_5_0_5 = sbox_AES_BoyarPeralta_21_port_o_0_5;
  assign subBytes_out_5_0_6 = sbox_AES_BoyarPeralta_21_port_o_0_6;
  assign subBytes_out_5_0_7 = sbox_AES_BoyarPeralta_21_port_o_0_7;
  assign subBytes_out_5_1_0 = sbox_AES_BoyarPeralta_21_port_o_1_0;
  assign subBytes_out_5_1_1 = sbox_AES_BoyarPeralta_21_port_o_1_1;
  assign subBytes_out_5_1_2 = sbox_AES_BoyarPeralta_21_port_o_1_2;
  assign subBytes_out_5_1_3 = sbox_AES_BoyarPeralta_21_port_o_1_3;
  assign subBytes_out_5_1_4 = sbox_AES_BoyarPeralta_21_port_o_1_4;
  assign subBytes_out_5_1_5 = sbox_AES_BoyarPeralta_21_port_o_1_5;
  assign subBytes_out_5_1_6 = sbox_AES_BoyarPeralta_21_port_o_1_6;
  assign subBytes_out_5_1_7 = sbox_AES_BoyarPeralta_21_port_o_1_7;
  assign subBytes_out_5_2_0 = sbox_AES_BoyarPeralta_21_port_o_2_0;
  assign subBytes_out_5_2_1 = sbox_AES_BoyarPeralta_21_port_o_2_1;
  assign subBytes_out_5_2_2 = sbox_AES_BoyarPeralta_21_port_o_2_2;
  assign subBytes_out_5_2_3 = sbox_AES_BoyarPeralta_21_port_o_2_3;
  assign subBytes_out_5_2_4 = sbox_AES_BoyarPeralta_21_port_o_2_4;
  assign subBytes_out_5_2_5 = sbox_AES_BoyarPeralta_21_port_o_2_5;
  assign subBytes_out_5_2_6 = sbox_AES_BoyarPeralta_21_port_o_2_6;
  assign subBytes_out_5_2_7 = sbox_AES_BoyarPeralta_21_port_o_2_7;
  assign subBytes_out_5_3_0 = sbox_AES_BoyarPeralta_21_port_o_3_0;
  assign subBytes_out_5_3_1 = sbox_AES_BoyarPeralta_21_port_o_3_1;
  assign subBytes_out_5_3_2 = sbox_AES_BoyarPeralta_21_port_o_3_2;
  assign subBytes_out_5_3_3 = sbox_AES_BoyarPeralta_21_port_o_3_3;
  assign subBytes_out_5_3_4 = sbox_AES_BoyarPeralta_21_port_o_3_4;
  assign subBytes_out_5_3_5 = sbox_AES_BoyarPeralta_21_port_o_3_5;
  assign subBytes_out_5_3_6 = sbox_AES_BoyarPeralta_21_port_o_3_6;
  assign subBytes_out_5_3_7 = sbox_AES_BoyarPeralta_21_port_o_3_7;
  assign subBytes_out_6_0_0 = sbox_AES_BoyarPeralta_22_port_o_0_0;
  assign subBytes_out_6_0_1 = sbox_AES_BoyarPeralta_22_port_o_0_1;
  assign subBytes_out_6_0_2 = sbox_AES_BoyarPeralta_22_port_o_0_2;
  assign subBytes_out_6_0_3 = sbox_AES_BoyarPeralta_22_port_o_0_3;
  assign subBytes_out_6_0_4 = sbox_AES_BoyarPeralta_22_port_o_0_4;
  assign subBytes_out_6_0_5 = sbox_AES_BoyarPeralta_22_port_o_0_5;
  assign subBytes_out_6_0_6 = sbox_AES_BoyarPeralta_22_port_o_0_6;
  assign subBytes_out_6_0_7 = sbox_AES_BoyarPeralta_22_port_o_0_7;
  assign subBytes_out_6_1_0 = sbox_AES_BoyarPeralta_22_port_o_1_0;
  assign subBytes_out_6_1_1 = sbox_AES_BoyarPeralta_22_port_o_1_1;
  assign subBytes_out_6_1_2 = sbox_AES_BoyarPeralta_22_port_o_1_2;
  assign subBytes_out_6_1_3 = sbox_AES_BoyarPeralta_22_port_o_1_3;
  assign subBytes_out_6_1_4 = sbox_AES_BoyarPeralta_22_port_o_1_4;
  assign subBytes_out_6_1_5 = sbox_AES_BoyarPeralta_22_port_o_1_5;
  assign subBytes_out_6_1_6 = sbox_AES_BoyarPeralta_22_port_o_1_6;
  assign subBytes_out_6_1_7 = sbox_AES_BoyarPeralta_22_port_o_1_7;
  assign subBytes_out_6_2_0 = sbox_AES_BoyarPeralta_22_port_o_2_0;
  assign subBytes_out_6_2_1 = sbox_AES_BoyarPeralta_22_port_o_2_1;
  assign subBytes_out_6_2_2 = sbox_AES_BoyarPeralta_22_port_o_2_2;
  assign subBytes_out_6_2_3 = sbox_AES_BoyarPeralta_22_port_o_2_3;
  assign subBytes_out_6_2_4 = sbox_AES_BoyarPeralta_22_port_o_2_4;
  assign subBytes_out_6_2_5 = sbox_AES_BoyarPeralta_22_port_o_2_5;
  assign subBytes_out_6_2_6 = sbox_AES_BoyarPeralta_22_port_o_2_6;
  assign subBytes_out_6_2_7 = sbox_AES_BoyarPeralta_22_port_o_2_7;
  assign subBytes_out_6_3_0 = sbox_AES_BoyarPeralta_22_port_o_3_0;
  assign subBytes_out_6_3_1 = sbox_AES_BoyarPeralta_22_port_o_3_1;
  assign subBytes_out_6_3_2 = sbox_AES_BoyarPeralta_22_port_o_3_2;
  assign subBytes_out_6_3_3 = sbox_AES_BoyarPeralta_22_port_o_3_3;
  assign subBytes_out_6_3_4 = sbox_AES_BoyarPeralta_22_port_o_3_4;
  assign subBytes_out_6_3_5 = sbox_AES_BoyarPeralta_22_port_o_3_5;
  assign subBytes_out_6_3_6 = sbox_AES_BoyarPeralta_22_port_o_3_6;
  assign subBytes_out_6_3_7 = sbox_AES_BoyarPeralta_22_port_o_3_7;
  assign subBytes_out_7_0_0 = sbox_AES_BoyarPeralta_23_port_o_0_0;
  assign subBytes_out_7_0_1 = sbox_AES_BoyarPeralta_23_port_o_0_1;
  assign subBytes_out_7_0_2 = sbox_AES_BoyarPeralta_23_port_o_0_2;
  assign subBytes_out_7_0_3 = sbox_AES_BoyarPeralta_23_port_o_0_3;
  assign subBytes_out_7_0_4 = sbox_AES_BoyarPeralta_23_port_o_0_4;
  assign subBytes_out_7_0_5 = sbox_AES_BoyarPeralta_23_port_o_0_5;
  assign subBytes_out_7_0_6 = sbox_AES_BoyarPeralta_23_port_o_0_6;
  assign subBytes_out_7_0_7 = sbox_AES_BoyarPeralta_23_port_o_0_7;
  assign subBytes_out_7_1_0 = sbox_AES_BoyarPeralta_23_port_o_1_0;
  assign subBytes_out_7_1_1 = sbox_AES_BoyarPeralta_23_port_o_1_1;
  assign subBytes_out_7_1_2 = sbox_AES_BoyarPeralta_23_port_o_1_2;
  assign subBytes_out_7_1_3 = sbox_AES_BoyarPeralta_23_port_o_1_3;
  assign subBytes_out_7_1_4 = sbox_AES_BoyarPeralta_23_port_o_1_4;
  assign subBytes_out_7_1_5 = sbox_AES_BoyarPeralta_23_port_o_1_5;
  assign subBytes_out_7_1_6 = sbox_AES_BoyarPeralta_23_port_o_1_6;
  assign subBytes_out_7_1_7 = sbox_AES_BoyarPeralta_23_port_o_1_7;
  assign subBytes_out_7_2_0 = sbox_AES_BoyarPeralta_23_port_o_2_0;
  assign subBytes_out_7_2_1 = sbox_AES_BoyarPeralta_23_port_o_2_1;
  assign subBytes_out_7_2_2 = sbox_AES_BoyarPeralta_23_port_o_2_2;
  assign subBytes_out_7_2_3 = sbox_AES_BoyarPeralta_23_port_o_2_3;
  assign subBytes_out_7_2_4 = sbox_AES_BoyarPeralta_23_port_o_2_4;
  assign subBytes_out_7_2_5 = sbox_AES_BoyarPeralta_23_port_o_2_5;
  assign subBytes_out_7_2_6 = sbox_AES_BoyarPeralta_23_port_o_2_6;
  assign subBytes_out_7_2_7 = sbox_AES_BoyarPeralta_23_port_o_2_7;
  assign subBytes_out_7_3_0 = sbox_AES_BoyarPeralta_23_port_o_3_0;
  assign subBytes_out_7_3_1 = sbox_AES_BoyarPeralta_23_port_o_3_1;
  assign subBytes_out_7_3_2 = sbox_AES_BoyarPeralta_23_port_o_3_2;
  assign subBytes_out_7_3_3 = sbox_AES_BoyarPeralta_23_port_o_3_3;
  assign subBytes_out_7_3_4 = sbox_AES_BoyarPeralta_23_port_o_3_4;
  assign subBytes_out_7_3_5 = sbox_AES_BoyarPeralta_23_port_o_3_5;
  assign subBytes_out_7_3_6 = sbox_AES_BoyarPeralta_23_port_o_3_6;
  assign subBytes_out_7_3_7 = sbox_AES_BoyarPeralta_23_port_o_3_7;
  assign subBytes_out_8_0_0 = sbox_AES_BoyarPeralta_24_port_o_0_0;
  assign subBytes_out_8_0_1 = sbox_AES_BoyarPeralta_24_port_o_0_1;
  assign subBytes_out_8_0_2 = sbox_AES_BoyarPeralta_24_port_o_0_2;
  assign subBytes_out_8_0_3 = sbox_AES_BoyarPeralta_24_port_o_0_3;
  assign subBytes_out_8_0_4 = sbox_AES_BoyarPeralta_24_port_o_0_4;
  assign subBytes_out_8_0_5 = sbox_AES_BoyarPeralta_24_port_o_0_5;
  assign subBytes_out_8_0_6 = sbox_AES_BoyarPeralta_24_port_o_0_6;
  assign subBytes_out_8_0_7 = sbox_AES_BoyarPeralta_24_port_o_0_7;
  assign subBytes_out_8_1_0 = sbox_AES_BoyarPeralta_24_port_o_1_0;
  assign subBytes_out_8_1_1 = sbox_AES_BoyarPeralta_24_port_o_1_1;
  assign subBytes_out_8_1_2 = sbox_AES_BoyarPeralta_24_port_o_1_2;
  assign subBytes_out_8_1_3 = sbox_AES_BoyarPeralta_24_port_o_1_3;
  assign subBytes_out_8_1_4 = sbox_AES_BoyarPeralta_24_port_o_1_4;
  assign subBytes_out_8_1_5 = sbox_AES_BoyarPeralta_24_port_o_1_5;
  assign subBytes_out_8_1_6 = sbox_AES_BoyarPeralta_24_port_o_1_6;
  assign subBytes_out_8_1_7 = sbox_AES_BoyarPeralta_24_port_o_1_7;
  assign subBytes_out_8_2_0 = sbox_AES_BoyarPeralta_24_port_o_2_0;
  assign subBytes_out_8_2_1 = sbox_AES_BoyarPeralta_24_port_o_2_1;
  assign subBytes_out_8_2_2 = sbox_AES_BoyarPeralta_24_port_o_2_2;
  assign subBytes_out_8_2_3 = sbox_AES_BoyarPeralta_24_port_o_2_3;
  assign subBytes_out_8_2_4 = sbox_AES_BoyarPeralta_24_port_o_2_4;
  assign subBytes_out_8_2_5 = sbox_AES_BoyarPeralta_24_port_o_2_5;
  assign subBytes_out_8_2_6 = sbox_AES_BoyarPeralta_24_port_o_2_6;
  assign subBytes_out_8_2_7 = sbox_AES_BoyarPeralta_24_port_o_2_7;
  assign subBytes_out_8_3_0 = sbox_AES_BoyarPeralta_24_port_o_3_0;
  assign subBytes_out_8_3_1 = sbox_AES_BoyarPeralta_24_port_o_3_1;
  assign subBytes_out_8_3_2 = sbox_AES_BoyarPeralta_24_port_o_3_2;
  assign subBytes_out_8_3_3 = sbox_AES_BoyarPeralta_24_port_o_3_3;
  assign subBytes_out_8_3_4 = sbox_AES_BoyarPeralta_24_port_o_3_4;
  assign subBytes_out_8_3_5 = sbox_AES_BoyarPeralta_24_port_o_3_5;
  assign subBytes_out_8_3_6 = sbox_AES_BoyarPeralta_24_port_o_3_6;
  assign subBytes_out_8_3_7 = sbox_AES_BoyarPeralta_24_port_o_3_7;
  assign subBytes_out_9_0_0 = sbox_AES_BoyarPeralta_25_port_o_0_0;
  assign subBytes_out_9_0_1 = sbox_AES_BoyarPeralta_25_port_o_0_1;
  assign subBytes_out_9_0_2 = sbox_AES_BoyarPeralta_25_port_o_0_2;
  assign subBytes_out_9_0_3 = sbox_AES_BoyarPeralta_25_port_o_0_3;
  assign subBytes_out_9_0_4 = sbox_AES_BoyarPeralta_25_port_o_0_4;
  assign subBytes_out_9_0_5 = sbox_AES_BoyarPeralta_25_port_o_0_5;
  assign subBytes_out_9_0_6 = sbox_AES_BoyarPeralta_25_port_o_0_6;
  assign subBytes_out_9_0_7 = sbox_AES_BoyarPeralta_25_port_o_0_7;
  assign subBytes_out_9_1_0 = sbox_AES_BoyarPeralta_25_port_o_1_0;
  assign subBytes_out_9_1_1 = sbox_AES_BoyarPeralta_25_port_o_1_1;
  assign subBytes_out_9_1_2 = sbox_AES_BoyarPeralta_25_port_o_1_2;
  assign subBytes_out_9_1_3 = sbox_AES_BoyarPeralta_25_port_o_1_3;
  assign subBytes_out_9_1_4 = sbox_AES_BoyarPeralta_25_port_o_1_4;
  assign subBytes_out_9_1_5 = sbox_AES_BoyarPeralta_25_port_o_1_5;
  assign subBytes_out_9_1_6 = sbox_AES_BoyarPeralta_25_port_o_1_6;
  assign subBytes_out_9_1_7 = sbox_AES_BoyarPeralta_25_port_o_1_7;
  assign subBytes_out_9_2_0 = sbox_AES_BoyarPeralta_25_port_o_2_0;
  assign subBytes_out_9_2_1 = sbox_AES_BoyarPeralta_25_port_o_2_1;
  assign subBytes_out_9_2_2 = sbox_AES_BoyarPeralta_25_port_o_2_2;
  assign subBytes_out_9_2_3 = sbox_AES_BoyarPeralta_25_port_o_2_3;
  assign subBytes_out_9_2_4 = sbox_AES_BoyarPeralta_25_port_o_2_4;
  assign subBytes_out_9_2_5 = sbox_AES_BoyarPeralta_25_port_o_2_5;
  assign subBytes_out_9_2_6 = sbox_AES_BoyarPeralta_25_port_o_2_6;
  assign subBytes_out_9_2_7 = sbox_AES_BoyarPeralta_25_port_o_2_7;
  assign subBytes_out_9_3_0 = sbox_AES_BoyarPeralta_25_port_o_3_0;
  assign subBytes_out_9_3_1 = sbox_AES_BoyarPeralta_25_port_o_3_1;
  assign subBytes_out_9_3_2 = sbox_AES_BoyarPeralta_25_port_o_3_2;
  assign subBytes_out_9_3_3 = sbox_AES_BoyarPeralta_25_port_o_3_3;
  assign subBytes_out_9_3_4 = sbox_AES_BoyarPeralta_25_port_o_3_4;
  assign subBytes_out_9_3_5 = sbox_AES_BoyarPeralta_25_port_o_3_5;
  assign subBytes_out_9_3_6 = sbox_AES_BoyarPeralta_25_port_o_3_6;
  assign subBytes_out_9_3_7 = sbox_AES_BoyarPeralta_25_port_o_3_7;
  assign subBytes_out_10_0_0 = sbox_AES_BoyarPeralta_26_port_o_0_0;
  assign subBytes_out_10_0_1 = sbox_AES_BoyarPeralta_26_port_o_0_1;
  assign subBytes_out_10_0_2 = sbox_AES_BoyarPeralta_26_port_o_0_2;
  assign subBytes_out_10_0_3 = sbox_AES_BoyarPeralta_26_port_o_0_3;
  assign subBytes_out_10_0_4 = sbox_AES_BoyarPeralta_26_port_o_0_4;
  assign subBytes_out_10_0_5 = sbox_AES_BoyarPeralta_26_port_o_0_5;
  assign subBytes_out_10_0_6 = sbox_AES_BoyarPeralta_26_port_o_0_6;
  assign subBytes_out_10_0_7 = sbox_AES_BoyarPeralta_26_port_o_0_7;
  assign subBytes_out_10_1_0 = sbox_AES_BoyarPeralta_26_port_o_1_0;
  assign subBytes_out_10_1_1 = sbox_AES_BoyarPeralta_26_port_o_1_1;
  assign subBytes_out_10_1_2 = sbox_AES_BoyarPeralta_26_port_o_1_2;
  assign subBytes_out_10_1_3 = sbox_AES_BoyarPeralta_26_port_o_1_3;
  assign subBytes_out_10_1_4 = sbox_AES_BoyarPeralta_26_port_o_1_4;
  assign subBytes_out_10_1_5 = sbox_AES_BoyarPeralta_26_port_o_1_5;
  assign subBytes_out_10_1_6 = sbox_AES_BoyarPeralta_26_port_o_1_6;
  assign subBytes_out_10_1_7 = sbox_AES_BoyarPeralta_26_port_o_1_7;
  assign subBytes_out_10_2_0 = sbox_AES_BoyarPeralta_26_port_o_2_0;
  assign subBytes_out_10_2_1 = sbox_AES_BoyarPeralta_26_port_o_2_1;
  assign subBytes_out_10_2_2 = sbox_AES_BoyarPeralta_26_port_o_2_2;
  assign subBytes_out_10_2_3 = sbox_AES_BoyarPeralta_26_port_o_2_3;
  assign subBytes_out_10_2_4 = sbox_AES_BoyarPeralta_26_port_o_2_4;
  assign subBytes_out_10_2_5 = sbox_AES_BoyarPeralta_26_port_o_2_5;
  assign subBytes_out_10_2_6 = sbox_AES_BoyarPeralta_26_port_o_2_6;
  assign subBytes_out_10_2_7 = sbox_AES_BoyarPeralta_26_port_o_2_7;
  assign subBytes_out_10_3_0 = sbox_AES_BoyarPeralta_26_port_o_3_0;
  assign subBytes_out_10_3_1 = sbox_AES_BoyarPeralta_26_port_o_3_1;
  assign subBytes_out_10_3_2 = sbox_AES_BoyarPeralta_26_port_o_3_2;
  assign subBytes_out_10_3_3 = sbox_AES_BoyarPeralta_26_port_o_3_3;
  assign subBytes_out_10_3_4 = sbox_AES_BoyarPeralta_26_port_o_3_4;
  assign subBytes_out_10_3_5 = sbox_AES_BoyarPeralta_26_port_o_3_5;
  assign subBytes_out_10_3_6 = sbox_AES_BoyarPeralta_26_port_o_3_6;
  assign subBytes_out_10_3_7 = sbox_AES_BoyarPeralta_26_port_o_3_7;
  assign subBytes_out_11_0_0 = sbox_AES_BoyarPeralta_27_port_o_0_0;
  assign subBytes_out_11_0_1 = sbox_AES_BoyarPeralta_27_port_o_0_1;
  assign subBytes_out_11_0_2 = sbox_AES_BoyarPeralta_27_port_o_0_2;
  assign subBytes_out_11_0_3 = sbox_AES_BoyarPeralta_27_port_o_0_3;
  assign subBytes_out_11_0_4 = sbox_AES_BoyarPeralta_27_port_o_0_4;
  assign subBytes_out_11_0_5 = sbox_AES_BoyarPeralta_27_port_o_0_5;
  assign subBytes_out_11_0_6 = sbox_AES_BoyarPeralta_27_port_o_0_6;
  assign subBytes_out_11_0_7 = sbox_AES_BoyarPeralta_27_port_o_0_7;
  assign subBytes_out_11_1_0 = sbox_AES_BoyarPeralta_27_port_o_1_0;
  assign subBytes_out_11_1_1 = sbox_AES_BoyarPeralta_27_port_o_1_1;
  assign subBytes_out_11_1_2 = sbox_AES_BoyarPeralta_27_port_o_1_2;
  assign subBytes_out_11_1_3 = sbox_AES_BoyarPeralta_27_port_o_1_3;
  assign subBytes_out_11_1_4 = sbox_AES_BoyarPeralta_27_port_o_1_4;
  assign subBytes_out_11_1_5 = sbox_AES_BoyarPeralta_27_port_o_1_5;
  assign subBytes_out_11_1_6 = sbox_AES_BoyarPeralta_27_port_o_1_6;
  assign subBytes_out_11_1_7 = sbox_AES_BoyarPeralta_27_port_o_1_7;
  assign subBytes_out_11_2_0 = sbox_AES_BoyarPeralta_27_port_o_2_0;
  assign subBytes_out_11_2_1 = sbox_AES_BoyarPeralta_27_port_o_2_1;
  assign subBytes_out_11_2_2 = sbox_AES_BoyarPeralta_27_port_o_2_2;
  assign subBytes_out_11_2_3 = sbox_AES_BoyarPeralta_27_port_o_2_3;
  assign subBytes_out_11_2_4 = sbox_AES_BoyarPeralta_27_port_o_2_4;
  assign subBytes_out_11_2_5 = sbox_AES_BoyarPeralta_27_port_o_2_5;
  assign subBytes_out_11_2_6 = sbox_AES_BoyarPeralta_27_port_o_2_6;
  assign subBytes_out_11_2_7 = sbox_AES_BoyarPeralta_27_port_o_2_7;
  assign subBytes_out_11_3_0 = sbox_AES_BoyarPeralta_27_port_o_3_0;
  assign subBytes_out_11_3_1 = sbox_AES_BoyarPeralta_27_port_o_3_1;
  assign subBytes_out_11_3_2 = sbox_AES_BoyarPeralta_27_port_o_3_2;
  assign subBytes_out_11_3_3 = sbox_AES_BoyarPeralta_27_port_o_3_3;
  assign subBytes_out_11_3_4 = sbox_AES_BoyarPeralta_27_port_o_3_4;
  assign subBytes_out_11_3_5 = sbox_AES_BoyarPeralta_27_port_o_3_5;
  assign subBytes_out_11_3_6 = sbox_AES_BoyarPeralta_27_port_o_3_6;
  assign subBytes_out_11_3_7 = sbox_AES_BoyarPeralta_27_port_o_3_7;
  assign subBytes_out_12_0_0 = sbox_AES_BoyarPeralta_28_port_o_0_0;
  assign subBytes_out_12_0_1 = sbox_AES_BoyarPeralta_28_port_o_0_1;
  assign subBytes_out_12_0_2 = sbox_AES_BoyarPeralta_28_port_o_0_2;
  assign subBytes_out_12_0_3 = sbox_AES_BoyarPeralta_28_port_o_0_3;
  assign subBytes_out_12_0_4 = sbox_AES_BoyarPeralta_28_port_o_0_4;
  assign subBytes_out_12_0_5 = sbox_AES_BoyarPeralta_28_port_o_0_5;
  assign subBytes_out_12_0_6 = sbox_AES_BoyarPeralta_28_port_o_0_6;
  assign subBytes_out_12_0_7 = sbox_AES_BoyarPeralta_28_port_o_0_7;
  assign subBytes_out_12_1_0 = sbox_AES_BoyarPeralta_28_port_o_1_0;
  assign subBytes_out_12_1_1 = sbox_AES_BoyarPeralta_28_port_o_1_1;
  assign subBytes_out_12_1_2 = sbox_AES_BoyarPeralta_28_port_o_1_2;
  assign subBytes_out_12_1_3 = sbox_AES_BoyarPeralta_28_port_o_1_3;
  assign subBytes_out_12_1_4 = sbox_AES_BoyarPeralta_28_port_o_1_4;
  assign subBytes_out_12_1_5 = sbox_AES_BoyarPeralta_28_port_o_1_5;
  assign subBytes_out_12_1_6 = sbox_AES_BoyarPeralta_28_port_o_1_6;
  assign subBytes_out_12_1_7 = sbox_AES_BoyarPeralta_28_port_o_1_7;
  assign subBytes_out_12_2_0 = sbox_AES_BoyarPeralta_28_port_o_2_0;
  assign subBytes_out_12_2_1 = sbox_AES_BoyarPeralta_28_port_o_2_1;
  assign subBytes_out_12_2_2 = sbox_AES_BoyarPeralta_28_port_o_2_2;
  assign subBytes_out_12_2_3 = sbox_AES_BoyarPeralta_28_port_o_2_3;
  assign subBytes_out_12_2_4 = sbox_AES_BoyarPeralta_28_port_o_2_4;
  assign subBytes_out_12_2_5 = sbox_AES_BoyarPeralta_28_port_o_2_5;
  assign subBytes_out_12_2_6 = sbox_AES_BoyarPeralta_28_port_o_2_6;
  assign subBytes_out_12_2_7 = sbox_AES_BoyarPeralta_28_port_o_2_7;
  assign subBytes_out_12_3_0 = sbox_AES_BoyarPeralta_28_port_o_3_0;
  assign subBytes_out_12_3_1 = sbox_AES_BoyarPeralta_28_port_o_3_1;
  assign subBytes_out_12_3_2 = sbox_AES_BoyarPeralta_28_port_o_3_2;
  assign subBytes_out_12_3_3 = sbox_AES_BoyarPeralta_28_port_o_3_3;
  assign subBytes_out_12_3_4 = sbox_AES_BoyarPeralta_28_port_o_3_4;
  assign subBytes_out_12_3_5 = sbox_AES_BoyarPeralta_28_port_o_3_5;
  assign subBytes_out_12_3_6 = sbox_AES_BoyarPeralta_28_port_o_3_6;
  assign subBytes_out_12_3_7 = sbox_AES_BoyarPeralta_28_port_o_3_7;
  assign subBytes_out_13_0_0 = sbox_AES_BoyarPeralta_29_port_o_0_0;
  assign subBytes_out_13_0_1 = sbox_AES_BoyarPeralta_29_port_o_0_1;
  assign subBytes_out_13_0_2 = sbox_AES_BoyarPeralta_29_port_o_0_2;
  assign subBytes_out_13_0_3 = sbox_AES_BoyarPeralta_29_port_o_0_3;
  assign subBytes_out_13_0_4 = sbox_AES_BoyarPeralta_29_port_o_0_4;
  assign subBytes_out_13_0_5 = sbox_AES_BoyarPeralta_29_port_o_0_5;
  assign subBytes_out_13_0_6 = sbox_AES_BoyarPeralta_29_port_o_0_6;
  assign subBytes_out_13_0_7 = sbox_AES_BoyarPeralta_29_port_o_0_7;
  assign subBytes_out_13_1_0 = sbox_AES_BoyarPeralta_29_port_o_1_0;
  assign subBytes_out_13_1_1 = sbox_AES_BoyarPeralta_29_port_o_1_1;
  assign subBytes_out_13_1_2 = sbox_AES_BoyarPeralta_29_port_o_1_2;
  assign subBytes_out_13_1_3 = sbox_AES_BoyarPeralta_29_port_o_1_3;
  assign subBytes_out_13_1_4 = sbox_AES_BoyarPeralta_29_port_o_1_4;
  assign subBytes_out_13_1_5 = sbox_AES_BoyarPeralta_29_port_o_1_5;
  assign subBytes_out_13_1_6 = sbox_AES_BoyarPeralta_29_port_o_1_6;
  assign subBytes_out_13_1_7 = sbox_AES_BoyarPeralta_29_port_o_1_7;
  assign subBytes_out_13_2_0 = sbox_AES_BoyarPeralta_29_port_o_2_0;
  assign subBytes_out_13_2_1 = sbox_AES_BoyarPeralta_29_port_o_2_1;
  assign subBytes_out_13_2_2 = sbox_AES_BoyarPeralta_29_port_o_2_2;
  assign subBytes_out_13_2_3 = sbox_AES_BoyarPeralta_29_port_o_2_3;
  assign subBytes_out_13_2_4 = sbox_AES_BoyarPeralta_29_port_o_2_4;
  assign subBytes_out_13_2_5 = sbox_AES_BoyarPeralta_29_port_o_2_5;
  assign subBytes_out_13_2_6 = sbox_AES_BoyarPeralta_29_port_o_2_6;
  assign subBytes_out_13_2_7 = sbox_AES_BoyarPeralta_29_port_o_2_7;
  assign subBytes_out_13_3_0 = sbox_AES_BoyarPeralta_29_port_o_3_0;
  assign subBytes_out_13_3_1 = sbox_AES_BoyarPeralta_29_port_o_3_1;
  assign subBytes_out_13_3_2 = sbox_AES_BoyarPeralta_29_port_o_3_2;
  assign subBytes_out_13_3_3 = sbox_AES_BoyarPeralta_29_port_o_3_3;
  assign subBytes_out_13_3_4 = sbox_AES_BoyarPeralta_29_port_o_3_4;
  assign subBytes_out_13_3_5 = sbox_AES_BoyarPeralta_29_port_o_3_5;
  assign subBytes_out_13_3_6 = sbox_AES_BoyarPeralta_29_port_o_3_6;
  assign subBytes_out_13_3_7 = sbox_AES_BoyarPeralta_29_port_o_3_7;
  assign subBytes_out_14_0_0 = sbox_AES_BoyarPeralta_30_port_o_0_0;
  assign subBytes_out_14_0_1 = sbox_AES_BoyarPeralta_30_port_o_0_1;
  assign subBytes_out_14_0_2 = sbox_AES_BoyarPeralta_30_port_o_0_2;
  assign subBytes_out_14_0_3 = sbox_AES_BoyarPeralta_30_port_o_0_3;
  assign subBytes_out_14_0_4 = sbox_AES_BoyarPeralta_30_port_o_0_4;
  assign subBytes_out_14_0_5 = sbox_AES_BoyarPeralta_30_port_o_0_5;
  assign subBytes_out_14_0_6 = sbox_AES_BoyarPeralta_30_port_o_0_6;
  assign subBytes_out_14_0_7 = sbox_AES_BoyarPeralta_30_port_o_0_7;
  assign subBytes_out_14_1_0 = sbox_AES_BoyarPeralta_30_port_o_1_0;
  assign subBytes_out_14_1_1 = sbox_AES_BoyarPeralta_30_port_o_1_1;
  assign subBytes_out_14_1_2 = sbox_AES_BoyarPeralta_30_port_o_1_2;
  assign subBytes_out_14_1_3 = sbox_AES_BoyarPeralta_30_port_o_1_3;
  assign subBytes_out_14_1_4 = sbox_AES_BoyarPeralta_30_port_o_1_4;
  assign subBytes_out_14_1_5 = sbox_AES_BoyarPeralta_30_port_o_1_5;
  assign subBytes_out_14_1_6 = sbox_AES_BoyarPeralta_30_port_o_1_6;
  assign subBytes_out_14_1_7 = sbox_AES_BoyarPeralta_30_port_o_1_7;
  assign subBytes_out_14_2_0 = sbox_AES_BoyarPeralta_30_port_o_2_0;
  assign subBytes_out_14_2_1 = sbox_AES_BoyarPeralta_30_port_o_2_1;
  assign subBytes_out_14_2_2 = sbox_AES_BoyarPeralta_30_port_o_2_2;
  assign subBytes_out_14_2_3 = sbox_AES_BoyarPeralta_30_port_o_2_3;
  assign subBytes_out_14_2_4 = sbox_AES_BoyarPeralta_30_port_o_2_4;
  assign subBytes_out_14_2_5 = sbox_AES_BoyarPeralta_30_port_o_2_5;
  assign subBytes_out_14_2_6 = sbox_AES_BoyarPeralta_30_port_o_2_6;
  assign subBytes_out_14_2_7 = sbox_AES_BoyarPeralta_30_port_o_2_7;
  assign subBytes_out_14_3_0 = sbox_AES_BoyarPeralta_30_port_o_3_0;
  assign subBytes_out_14_3_1 = sbox_AES_BoyarPeralta_30_port_o_3_1;
  assign subBytes_out_14_3_2 = sbox_AES_BoyarPeralta_30_port_o_3_2;
  assign subBytes_out_14_3_3 = sbox_AES_BoyarPeralta_30_port_o_3_3;
  assign subBytes_out_14_3_4 = sbox_AES_BoyarPeralta_30_port_o_3_4;
  assign subBytes_out_14_3_5 = sbox_AES_BoyarPeralta_30_port_o_3_5;
  assign subBytes_out_14_3_6 = sbox_AES_BoyarPeralta_30_port_o_3_6;
  assign subBytes_out_14_3_7 = sbox_AES_BoyarPeralta_30_port_o_3_7;
  assign subBytes_out_15_0_0 = sbox_AES_BoyarPeralta_31_port_o_0_0;
  assign subBytes_out_15_0_1 = sbox_AES_BoyarPeralta_31_port_o_0_1;
  assign subBytes_out_15_0_2 = sbox_AES_BoyarPeralta_31_port_o_0_2;
  assign subBytes_out_15_0_3 = sbox_AES_BoyarPeralta_31_port_o_0_3;
  assign subBytes_out_15_0_4 = sbox_AES_BoyarPeralta_31_port_o_0_4;
  assign subBytes_out_15_0_5 = sbox_AES_BoyarPeralta_31_port_o_0_5;
  assign subBytes_out_15_0_6 = sbox_AES_BoyarPeralta_31_port_o_0_6;
  assign subBytes_out_15_0_7 = sbox_AES_BoyarPeralta_31_port_o_0_7;
  assign subBytes_out_15_1_0 = sbox_AES_BoyarPeralta_31_port_o_1_0;
  assign subBytes_out_15_1_1 = sbox_AES_BoyarPeralta_31_port_o_1_1;
  assign subBytes_out_15_1_2 = sbox_AES_BoyarPeralta_31_port_o_1_2;
  assign subBytes_out_15_1_3 = sbox_AES_BoyarPeralta_31_port_o_1_3;
  assign subBytes_out_15_1_4 = sbox_AES_BoyarPeralta_31_port_o_1_4;
  assign subBytes_out_15_1_5 = sbox_AES_BoyarPeralta_31_port_o_1_5;
  assign subBytes_out_15_1_6 = sbox_AES_BoyarPeralta_31_port_o_1_6;
  assign subBytes_out_15_1_7 = sbox_AES_BoyarPeralta_31_port_o_1_7;
  assign subBytes_out_15_2_0 = sbox_AES_BoyarPeralta_31_port_o_2_0;
  assign subBytes_out_15_2_1 = sbox_AES_BoyarPeralta_31_port_o_2_1;
  assign subBytes_out_15_2_2 = sbox_AES_BoyarPeralta_31_port_o_2_2;
  assign subBytes_out_15_2_3 = sbox_AES_BoyarPeralta_31_port_o_2_3;
  assign subBytes_out_15_2_4 = sbox_AES_BoyarPeralta_31_port_o_2_4;
  assign subBytes_out_15_2_5 = sbox_AES_BoyarPeralta_31_port_o_2_5;
  assign subBytes_out_15_2_6 = sbox_AES_BoyarPeralta_31_port_o_2_6;
  assign subBytes_out_15_2_7 = sbox_AES_BoyarPeralta_31_port_o_2_7;
  assign subBytes_out_15_3_0 = sbox_AES_BoyarPeralta_31_port_o_3_0;
  assign subBytes_out_15_3_1 = sbox_AES_BoyarPeralta_31_port_o_3_1;
  assign subBytes_out_15_3_2 = sbox_AES_BoyarPeralta_31_port_o_3_2;
  assign subBytes_out_15_3_3 = sbox_AES_BoyarPeralta_31_port_o_3_3;
  assign subBytes_out_15_3_4 = sbox_AES_BoyarPeralta_31_port_o_3_4;
  assign subBytes_out_15_3_5 = sbox_AES_BoyarPeralta_31_port_o_3_5;
  assign subBytes_out_15_3_6 = sbox_AES_BoyarPeralta_31_port_o_3_6;
  assign subBytes_out_15_3_7 = sbox_AES_BoyarPeralta_31_port_o_3_7;
  assign port_state_out_0_0_0 = roundReg_0_0_0;
  assign port_state_out_0_0_1 = roundReg_0_0_1;
  assign port_state_out_0_0_2 = roundReg_0_0_2;
  assign port_state_out_0_0_3 = roundReg_0_0_3;
  assign port_state_out_0_0_4 = roundReg_0_0_4;
  assign port_state_out_0_0_5 = roundReg_0_0_5;
  assign port_state_out_0_0_6 = roundReg_0_0_6;
  assign port_state_out_0_0_7 = roundReg_0_0_7;
  assign port_state_out_0_1_0 = roundReg_0_1_0;
  assign port_state_out_0_1_1 = roundReg_0_1_1;
  assign port_state_out_0_1_2 = roundReg_0_1_2;
  assign port_state_out_0_1_3 = roundReg_0_1_3;
  assign port_state_out_0_1_4 = roundReg_0_1_4;
  assign port_state_out_0_1_5 = roundReg_0_1_5;
  assign port_state_out_0_1_6 = roundReg_0_1_6;
  assign port_state_out_0_1_7 = roundReg_0_1_7;
  assign port_state_out_0_2_0 = roundReg_0_2_0;
  assign port_state_out_0_2_1 = roundReg_0_2_1;
  assign port_state_out_0_2_2 = roundReg_0_2_2;
  assign port_state_out_0_2_3 = roundReg_0_2_3;
  assign port_state_out_0_2_4 = roundReg_0_2_4;
  assign port_state_out_0_2_5 = roundReg_0_2_5;
  assign port_state_out_0_2_6 = roundReg_0_2_6;
  assign port_state_out_0_2_7 = roundReg_0_2_7;
  assign port_state_out_0_3_0 = roundReg_0_3_0;
  assign port_state_out_0_3_1 = roundReg_0_3_1;
  assign port_state_out_0_3_2 = roundReg_0_3_2;
  assign port_state_out_0_3_3 = roundReg_0_3_3;
  assign port_state_out_0_3_4 = roundReg_0_3_4;
  assign port_state_out_0_3_5 = roundReg_0_3_5;
  assign port_state_out_0_3_6 = roundReg_0_3_6;
  assign port_state_out_0_3_7 = roundReg_0_3_7;
  assign port_state_out_1_0_0 = roundReg_1_0_0;
  assign port_state_out_1_0_1 = roundReg_1_0_1;
  assign port_state_out_1_0_2 = roundReg_1_0_2;
  assign port_state_out_1_0_3 = roundReg_1_0_3;
  assign port_state_out_1_0_4 = roundReg_1_0_4;
  assign port_state_out_1_0_5 = roundReg_1_0_5;
  assign port_state_out_1_0_6 = roundReg_1_0_6;
  assign port_state_out_1_0_7 = roundReg_1_0_7;
  assign port_state_out_1_1_0 = roundReg_1_1_0;
  assign port_state_out_1_1_1 = roundReg_1_1_1;
  assign port_state_out_1_1_2 = roundReg_1_1_2;
  assign port_state_out_1_1_3 = roundReg_1_1_3;
  assign port_state_out_1_1_4 = roundReg_1_1_4;
  assign port_state_out_1_1_5 = roundReg_1_1_5;
  assign port_state_out_1_1_6 = roundReg_1_1_6;
  assign port_state_out_1_1_7 = roundReg_1_1_7;
  assign port_state_out_1_2_0 = roundReg_1_2_0;
  assign port_state_out_1_2_1 = roundReg_1_2_1;
  assign port_state_out_1_2_2 = roundReg_1_2_2;
  assign port_state_out_1_2_3 = roundReg_1_2_3;
  assign port_state_out_1_2_4 = roundReg_1_2_4;
  assign port_state_out_1_2_5 = roundReg_1_2_5;
  assign port_state_out_1_2_6 = roundReg_1_2_6;
  assign port_state_out_1_2_7 = roundReg_1_2_7;
  assign port_state_out_1_3_0 = roundReg_1_3_0;
  assign port_state_out_1_3_1 = roundReg_1_3_1;
  assign port_state_out_1_3_2 = roundReg_1_3_2;
  assign port_state_out_1_3_3 = roundReg_1_3_3;
  assign port_state_out_1_3_4 = roundReg_1_3_4;
  assign port_state_out_1_3_5 = roundReg_1_3_5;
  assign port_state_out_1_3_6 = roundReg_1_3_6;
  assign port_state_out_1_3_7 = roundReg_1_3_7;
  assign port_state_out_2_0_0 = roundReg_2_0_0;
  assign port_state_out_2_0_1 = roundReg_2_0_1;
  assign port_state_out_2_0_2 = roundReg_2_0_2;
  assign port_state_out_2_0_3 = roundReg_2_0_3;
  assign port_state_out_2_0_4 = roundReg_2_0_4;
  assign port_state_out_2_0_5 = roundReg_2_0_5;
  assign port_state_out_2_0_6 = roundReg_2_0_6;
  assign port_state_out_2_0_7 = roundReg_2_0_7;
  assign port_state_out_2_1_0 = roundReg_2_1_0;
  assign port_state_out_2_1_1 = roundReg_2_1_1;
  assign port_state_out_2_1_2 = roundReg_2_1_2;
  assign port_state_out_2_1_3 = roundReg_2_1_3;
  assign port_state_out_2_1_4 = roundReg_2_1_4;
  assign port_state_out_2_1_5 = roundReg_2_1_5;
  assign port_state_out_2_1_6 = roundReg_2_1_6;
  assign port_state_out_2_1_7 = roundReg_2_1_7;
  assign port_state_out_2_2_0 = roundReg_2_2_0;
  assign port_state_out_2_2_1 = roundReg_2_2_1;
  assign port_state_out_2_2_2 = roundReg_2_2_2;
  assign port_state_out_2_2_3 = roundReg_2_2_3;
  assign port_state_out_2_2_4 = roundReg_2_2_4;
  assign port_state_out_2_2_5 = roundReg_2_2_5;
  assign port_state_out_2_2_6 = roundReg_2_2_6;
  assign port_state_out_2_2_7 = roundReg_2_2_7;
  assign port_state_out_2_3_0 = roundReg_2_3_0;
  assign port_state_out_2_3_1 = roundReg_2_3_1;
  assign port_state_out_2_3_2 = roundReg_2_3_2;
  assign port_state_out_2_3_3 = roundReg_2_3_3;
  assign port_state_out_2_3_4 = roundReg_2_3_4;
  assign port_state_out_2_3_5 = roundReg_2_3_5;
  assign port_state_out_2_3_6 = roundReg_2_3_6;
  assign port_state_out_2_3_7 = roundReg_2_3_7;
  assign port_state_out_3_0_0 = roundReg_3_0_0;
  assign port_state_out_3_0_1 = roundReg_3_0_1;
  assign port_state_out_3_0_2 = roundReg_3_0_2;
  assign port_state_out_3_0_3 = roundReg_3_0_3;
  assign port_state_out_3_0_4 = roundReg_3_0_4;
  assign port_state_out_3_0_5 = roundReg_3_0_5;
  assign port_state_out_3_0_6 = roundReg_3_0_6;
  assign port_state_out_3_0_7 = roundReg_3_0_7;
  assign port_state_out_3_1_0 = roundReg_3_1_0;
  assign port_state_out_3_1_1 = roundReg_3_1_1;
  assign port_state_out_3_1_2 = roundReg_3_1_2;
  assign port_state_out_3_1_3 = roundReg_3_1_3;
  assign port_state_out_3_1_4 = roundReg_3_1_4;
  assign port_state_out_3_1_5 = roundReg_3_1_5;
  assign port_state_out_3_1_6 = roundReg_3_1_6;
  assign port_state_out_3_1_7 = roundReg_3_1_7;
  assign port_state_out_3_2_0 = roundReg_3_2_0;
  assign port_state_out_3_2_1 = roundReg_3_2_1;
  assign port_state_out_3_2_2 = roundReg_3_2_2;
  assign port_state_out_3_2_3 = roundReg_3_2_3;
  assign port_state_out_3_2_4 = roundReg_3_2_4;
  assign port_state_out_3_2_5 = roundReg_3_2_5;
  assign port_state_out_3_2_6 = roundReg_3_2_6;
  assign port_state_out_3_2_7 = roundReg_3_2_7;
  assign port_state_out_3_3_0 = roundReg_3_3_0;
  assign port_state_out_3_3_1 = roundReg_3_3_1;
  assign port_state_out_3_3_2 = roundReg_3_3_2;
  assign port_state_out_3_3_3 = roundReg_3_3_3;
  assign port_state_out_3_3_4 = roundReg_3_3_4;
  assign port_state_out_3_3_5 = roundReg_3_3_5;
  assign port_state_out_3_3_6 = roundReg_3_3_6;
  assign port_state_out_3_3_7 = roundReg_3_3_7;
  assign port_state_out_4_0_0 = roundReg_4_0_0;
  assign port_state_out_4_0_1 = roundReg_4_0_1;
  assign port_state_out_4_0_2 = roundReg_4_0_2;
  assign port_state_out_4_0_3 = roundReg_4_0_3;
  assign port_state_out_4_0_4 = roundReg_4_0_4;
  assign port_state_out_4_0_5 = roundReg_4_0_5;
  assign port_state_out_4_0_6 = roundReg_4_0_6;
  assign port_state_out_4_0_7 = roundReg_4_0_7;
  assign port_state_out_4_1_0 = roundReg_4_1_0;
  assign port_state_out_4_1_1 = roundReg_4_1_1;
  assign port_state_out_4_1_2 = roundReg_4_1_2;
  assign port_state_out_4_1_3 = roundReg_4_1_3;
  assign port_state_out_4_1_4 = roundReg_4_1_4;
  assign port_state_out_4_1_5 = roundReg_4_1_5;
  assign port_state_out_4_1_6 = roundReg_4_1_6;
  assign port_state_out_4_1_7 = roundReg_4_1_7;
  assign port_state_out_4_2_0 = roundReg_4_2_0;
  assign port_state_out_4_2_1 = roundReg_4_2_1;
  assign port_state_out_4_2_2 = roundReg_4_2_2;
  assign port_state_out_4_2_3 = roundReg_4_2_3;
  assign port_state_out_4_2_4 = roundReg_4_2_4;
  assign port_state_out_4_2_5 = roundReg_4_2_5;
  assign port_state_out_4_2_6 = roundReg_4_2_6;
  assign port_state_out_4_2_7 = roundReg_4_2_7;
  assign port_state_out_4_3_0 = roundReg_4_3_0;
  assign port_state_out_4_3_1 = roundReg_4_3_1;
  assign port_state_out_4_3_2 = roundReg_4_3_2;
  assign port_state_out_4_3_3 = roundReg_4_3_3;
  assign port_state_out_4_3_4 = roundReg_4_3_4;
  assign port_state_out_4_3_5 = roundReg_4_3_5;
  assign port_state_out_4_3_6 = roundReg_4_3_6;
  assign port_state_out_4_3_7 = roundReg_4_3_7;
  assign port_state_out_5_0_0 = roundReg_5_0_0;
  assign port_state_out_5_0_1 = roundReg_5_0_1;
  assign port_state_out_5_0_2 = roundReg_5_0_2;
  assign port_state_out_5_0_3 = roundReg_5_0_3;
  assign port_state_out_5_0_4 = roundReg_5_0_4;
  assign port_state_out_5_0_5 = roundReg_5_0_5;
  assign port_state_out_5_0_6 = roundReg_5_0_6;
  assign port_state_out_5_0_7 = roundReg_5_0_7;
  assign port_state_out_5_1_0 = roundReg_5_1_0;
  assign port_state_out_5_1_1 = roundReg_5_1_1;
  assign port_state_out_5_1_2 = roundReg_5_1_2;
  assign port_state_out_5_1_3 = roundReg_5_1_3;
  assign port_state_out_5_1_4 = roundReg_5_1_4;
  assign port_state_out_5_1_5 = roundReg_5_1_5;
  assign port_state_out_5_1_6 = roundReg_5_1_6;
  assign port_state_out_5_1_7 = roundReg_5_1_7;
  assign port_state_out_5_2_0 = roundReg_5_2_0;
  assign port_state_out_5_2_1 = roundReg_5_2_1;
  assign port_state_out_5_2_2 = roundReg_5_2_2;
  assign port_state_out_5_2_3 = roundReg_5_2_3;
  assign port_state_out_5_2_4 = roundReg_5_2_4;
  assign port_state_out_5_2_5 = roundReg_5_2_5;
  assign port_state_out_5_2_6 = roundReg_5_2_6;
  assign port_state_out_5_2_7 = roundReg_5_2_7;
  assign port_state_out_5_3_0 = roundReg_5_3_0;
  assign port_state_out_5_3_1 = roundReg_5_3_1;
  assign port_state_out_5_3_2 = roundReg_5_3_2;
  assign port_state_out_5_3_3 = roundReg_5_3_3;
  assign port_state_out_5_3_4 = roundReg_5_3_4;
  assign port_state_out_5_3_5 = roundReg_5_3_5;
  assign port_state_out_5_3_6 = roundReg_5_3_6;
  assign port_state_out_5_3_7 = roundReg_5_3_7;
  assign port_state_out_6_0_0 = roundReg_6_0_0;
  assign port_state_out_6_0_1 = roundReg_6_0_1;
  assign port_state_out_6_0_2 = roundReg_6_0_2;
  assign port_state_out_6_0_3 = roundReg_6_0_3;
  assign port_state_out_6_0_4 = roundReg_6_0_4;
  assign port_state_out_6_0_5 = roundReg_6_0_5;
  assign port_state_out_6_0_6 = roundReg_6_0_6;
  assign port_state_out_6_0_7 = roundReg_6_0_7;
  assign port_state_out_6_1_0 = roundReg_6_1_0;
  assign port_state_out_6_1_1 = roundReg_6_1_1;
  assign port_state_out_6_1_2 = roundReg_6_1_2;
  assign port_state_out_6_1_3 = roundReg_6_1_3;
  assign port_state_out_6_1_4 = roundReg_6_1_4;
  assign port_state_out_6_1_5 = roundReg_6_1_5;
  assign port_state_out_6_1_6 = roundReg_6_1_6;
  assign port_state_out_6_1_7 = roundReg_6_1_7;
  assign port_state_out_6_2_0 = roundReg_6_2_0;
  assign port_state_out_6_2_1 = roundReg_6_2_1;
  assign port_state_out_6_2_2 = roundReg_6_2_2;
  assign port_state_out_6_2_3 = roundReg_6_2_3;
  assign port_state_out_6_2_4 = roundReg_6_2_4;
  assign port_state_out_6_2_5 = roundReg_6_2_5;
  assign port_state_out_6_2_6 = roundReg_6_2_6;
  assign port_state_out_6_2_7 = roundReg_6_2_7;
  assign port_state_out_6_3_0 = roundReg_6_3_0;
  assign port_state_out_6_3_1 = roundReg_6_3_1;
  assign port_state_out_6_3_2 = roundReg_6_3_2;
  assign port_state_out_6_3_3 = roundReg_6_3_3;
  assign port_state_out_6_3_4 = roundReg_6_3_4;
  assign port_state_out_6_3_5 = roundReg_6_3_5;
  assign port_state_out_6_3_6 = roundReg_6_3_6;
  assign port_state_out_6_3_7 = roundReg_6_3_7;
  assign port_state_out_7_0_0 = roundReg_7_0_0;
  assign port_state_out_7_0_1 = roundReg_7_0_1;
  assign port_state_out_7_0_2 = roundReg_7_0_2;
  assign port_state_out_7_0_3 = roundReg_7_0_3;
  assign port_state_out_7_0_4 = roundReg_7_0_4;
  assign port_state_out_7_0_5 = roundReg_7_0_5;
  assign port_state_out_7_0_6 = roundReg_7_0_6;
  assign port_state_out_7_0_7 = roundReg_7_0_7;
  assign port_state_out_7_1_0 = roundReg_7_1_0;
  assign port_state_out_7_1_1 = roundReg_7_1_1;
  assign port_state_out_7_1_2 = roundReg_7_1_2;
  assign port_state_out_7_1_3 = roundReg_7_1_3;
  assign port_state_out_7_1_4 = roundReg_7_1_4;
  assign port_state_out_7_1_5 = roundReg_7_1_5;
  assign port_state_out_7_1_6 = roundReg_7_1_6;
  assign port_state_out_7_1_7 = roundReg_7_1_7;
  assign port_state_out_7_2_0 = roundReg_7_2_0;
  assign port_state_out_7_2_1 = roundReg_7_2_1;
  assign port_state_out_7_2_2 = roundReg_7_2_2;
  assign port_state_out_7_2_3 = roundReg_7_2_3;
  assign port_state_out_7_2_4 = roundReg_7_2_4;
  assign port_state_out_7_2_5 = roundReg_7_2_5;
  assign port_state_out_7_2_6 = roundReg_7_2_6;
  assign port_state_out_7_2_7 = roundReg_7_2_7;
  assign port_state_out_7_3_0 = roundReg_7_3_0;
  assign port_state_out_7_3_1 = roundReg_7_3_1;
  assign port_state_out_7_3_2 = roundReg_7_3_2;
  assign port_state_out_7_3_3 = roundReg_7_3_3;
  assign port_state_out_7_3_4 = roundReg_7_3_4;
  assign port_state_out_7_3_5 = roundReg_7_3_5;
  assign port_state_out_7_3_6 = roundReg_7_3_6;
  assign port_state_out_7_3_7 = roundReg_7_3_7;
  assign port_state_out_8_0_0 = roundReg_8_0_0;
  assign port_state_out_8_0_1 = roundReg_8_0_1;
  assign port_state_out_8_0_2 = roundReg_8_0_2;
  assign port_state_out_8_0_3 = roundReg_8_0_3;
  assign port_state_out_8_0_4 = roundReg_8_0_4;
  assign port_state_out_8_0_5 = roundReg_8_0_5;
  assign port_state_out_8_0_6 = roundReg_8_0_6;
  assign port_state_out_8_0_7 = roundReg_8_0_7;
  assign port_state_out_8_1_0 = roundReg_8_1_0;
  assign port_state_out_8_1_1 = roundReg_8_1_1;
  assign port_state_out_8_1_2 = roundReg_8_1_2;
  assign port_state_out_8_1_3 = roundReg_8_1_3;
  assign port_state_out_8_1_4 = roundReg_8_1_4;
  assign port_state_out_8_1_5 = roundReg_8_1_5;
  assign port_state_out_8_1_6 = roundReg_8_1_6;
  assign port_state_out_8_1_7 = roundReg_8_1_7;
  assign port_state_out_8_2_0 = roundReg_8_2_0;
  assign port_state_out_8_2_1 = roundReg_8_2_1;
  assign port_state_out_8_2_2 = roundReg_8_2_2;
  assign port_state_out_8_2_3 = roundReg_8_2_3;
  assign port_state_out_8_2_4 = roundReg_8_2_4;
  assign port_state_out_8_2_5 = roundReg_8_2_5;
  assign port_state_out_8_2_6 = roundReg_8_2_6;
  assign port_state_out_8_2_7 = roundReg_8_2_7;
  assign port_state_out_8_3_0 = roundReg_8_3_0;
  assign port_state_out_8_3_1 = roundReg_8_3_1;
  assign port_state_out_8_3_2 = roundReg_8_3_2;
  assign port_state_out_8_3_3 = roundReg_8_3_3;
  assign port_state_out_8_3_4 = roundReg_8_3_4;
  assign port_state_out_8_3_5 = roundReg_8_3_5;
  assign port_state_out_8_3_6 = roundReg_8_3_6;
  assign port_state_out_8_3_7 = roundReg_8_3_7;
  assign port_state_out_9_0_0 = roundReg_9_0_0;
  assign port_state_out_9_0_1 = roundReg_9_0_1;
  assign port_state_out_9_0_2 = roundReg_9_0_2;
  assign port_state_out_9_0_3 = roundReg_9_0_3;
  assign port_state_out_9_0_4 = roundReg_9_0_4;
  assign port_state_out_9_0_5 = roundReg_9_0_5;
  assign port_state_out_9_0_6 = roundReg_9_0_6;
  assign port_state_out_9_0_7 = roundReg_9_0_7;
  assign port_state_out_9_1_0 = roundReg_9_1_0;
  assign port_state_out_9_1_1 = roundReg_9_1_1;
  assign port_state_out_9_1_2 = roundReg_9_1_2;
  assign port_state_out_9_1_3 = roundReg_9_1_3;
  assign port_state_out_9_1_4 = roundReg_9_1_4;
  assign port_state_out_9_1_5 = roundReg_9_1_5;
  assign port_state_out_9_1_6 = roundReg_9_1_6;
  assign port_state_out_9_1_7 = roundReg_9_1_7;
  assign port_state_out_9_2_0 = roundReg_9_2_0;
  assign port_state_out_9_2_1 = roundReg_9_2_1;
  assign port_state_out_9_2_2 = roundReg_9_2_2;
  assign port_state_out_9_2_3 = roundReg_9_2_3;
  assign port_state_out_9_2_4 = roundReg_9_2_4;
  assign port_state_out_9_2_5 = roundReg_9_2_5;
  assign port_state_out_9_2_6 = roundReg_9_2_6;
  assign port_state_out_9_2_7 = roundReg_9_2_7;
  assign port_state_out_9_3_0 = roundReg_9_3_0;
  assign port_state_out_9_3_1 = roundReg_9_3_1;
  assign port_state_out_9_3_2 = roundReg_9_3_2;
  assign port_state_out_9_3_3 = roundReg_9_3_3;
  assign port_state_out_9_3_4 = roundReg_9_3_4;
  assign port_state_out_9_3_5 = roundReg_9_3_5;
  assign port_state_out_9_3_6 = roundReg_9_3_6;
  assign port_state_out_9_3_7 = roundReg_9_3_7;
  assign port_state_out_10_0_0 = roundReg_10_0_0;
  assign port_state_out_10_0_1 = roundReg_10_0_1;
  assign port_state_out_10_0_2 = roundReg_10_0_2;
  assign port_state_out_10_0_3 = roundReg_10_0_3;
  assign port_state_out_10_0_4 = roundReg_10_0_4;
  assign port_state_out_10_0_5 = roundReg_10_0_5;
  assign port_state_out_10_0_6 = roundReg_10_0_6;
  assign port_state_out_10_0_7 = roundReg_10_0_7;
  assign port_state_out_10_1_0 = roundReg_10_1_0;
  assign port_state_out_10_1_1 = roundReg_10_1_1;
  assign port_state_out_10_1_2 = roundReg_10_1_2;
  assign port_state_out_10_1_3 = roundReg_10_1_3;
  assign port_state_out_10_1_4 = roundReg_10_1_4;
  assign port_state_out_10_1_5 = roundReg_10_1_5;
  assign port_state_out_10_1_6 = roundReg_10_1_6;
  assign port_state_out_10_1_7 = roundReg_10_1_7;
  assign port_state_out_10_2_0 = roundReg_10_2_0;
  assign port_state_out_10_2_1 = roundReg_10_2_1;
  assign port_state_out_10_2_2 = roundReg_10_2_2;
  assign port_state_out_10_2_3 = roundReg_10_2_3;
  assign port_state_out_10_2_4 = roundReg_10_2_4;
  assign port_state_out_10_2_5 = roundReg_10_2_5;
  assign port_state_out_10_2_6 = roundReg_10_2_6;
  assign port_state_out_10_2_7 = roundReg_10_2_7;
  assign port_state_out_10_3_0 = roundReg_10_3_0;
  assign port_state_out_10_3_1 = roundReg_10_3_1;
  assign port_state_out_10_3_2 = roundReg_10_3_2;
  assign port_state_out_10_3_3 = roundReg_10_3_3;
  assign port_state_out_10_3_4 = roundReg_10_3_4;
  assign port_state_out_10_3_5 = roundReg_10_3_5;
  assign port_state_out_10_3_6 = roundReg_10_3_6;
  assign port_state_out_10_3_7 = roundReg_10_3_7;
  assign port_state_out_11_0_0 = roundReg_11_0_0;
  assign port_state_out_11_0_1 = roundReg_11_0_1;
  assign port_state_out_11_0_2 = roundReg_11_0_2;
  assign port_state_out_11_0_3 = roundReg_11_0_3;
  assign port_state_out_11_0_4 = roundReg_11_0_4;
  assign port_state_out_11_0_5 = roundReg_11_0_5;
  assign port_state_out_11_0_6 = roundReg_11_0_6;
  assign port_state_out_11_0_7 = roundReg_11_0_7;
  assign port_state_out_11_1_0 = roundReg_11_1_0;
  assign port_state_out_11_1_1 = roundReg_11_1_1;
  assign port_state_out_11_1_2 = roundReg_11_1_2;
  assign port_state_out_11_1_3 = roundReg_11_1_3;
  assign port_state_out_11_1_4 = roundReg_11_1_4;
  assign port_state_out_11_1_5 = roundReg_11_1_5;
  assign port_state_out_11_1_6 = roundReg_11_1_6;
  assign port_state_out_11_1_7 = roundReg_11_1_7;
  assign port_state_out_11_2_0 = roundReg_11_2_0;
  assign port_state_out_11_2_1 = roundReg_11_2_1;
  assign port_state_out_11_2_2 = roundReg_11_2_2;
  assign port_state_out_11_2_3 = roundReg_11_2_3;
  assign port_state_out_11_2_4 = roundReg_11_2_4;
  assign port_state_out_11_2_5 = roundReg_11_2_5;
  assign port_state_out_11_2_6 = roundReg_11_2_6;
  assign port_state_out_11_2_7 = roundReg_11_2_7;
  assign port_state_out_11_3_0 = roundReg_11_3_0;
  assign port_state_out_11_3_1 = roundReg_11_3_1;
  assign port_state_out_11_3_2 = roundReg_11_3_2;
  assign port_state_out_11_3_3 = roundReg_11_3_3;
  assign port_state_out_11_3_4 = roundReg_11_3_4;
  assign port_state_out_11_3_5 = roundReg_11_3_5;
  assign port_state_out_11_3_6 = roundReg_11_3_6;
  assign port_state_out_11_3_7 = roundReg_11_3_7;
  assign port_state_out_12_0_0 = roundReg_12_0_0;
  assign port_state_out_12_0_1 = roundReg_12_0_1;
  assign port_state_out_12_0_2 = roundReg_12_0_2;
  assign port_state_out_12_0_3 = roundReg_12_0_3;
  assign port_state_out_12_0_4 = roundReg_12_0_4;
  assign port_state_out_12_0_5 = roundReg_12_0_5;
  assign port_state_out_12_0_6 = roundReg_12_0_6;
  assign port_state_out_12_0_7 = roundReg_12_0_7;
  assign port_state_out_12_1_0 = roundReg_12_1_0;
  assign port_state_out_12_1_1 = roundReg_12_1_1;
  assign port_state_out_12_1_2 = roundReg_12_1_2;
  assign port_state_out_12_1_3 = roundReg_12_1_3;
  assign port_state_out_12_1_4 = roundReg_12_1_4;
  assign port_state_out_12_1_5 = roundReg_12_1_5;
  assign port_state_out_12_1_6 = roundReg_12_1_6;
  assign port_state_out_12_1_7 = roundReg_12_1_7;
  assign port_state_out_12_2_0 = roundReg_12_2_0;
  assign port_state_out_12_2_1 = roundReg_12_2_1;
  assign port_state_out_12_2_2 = roundReg_12_2_2;
  assign port_state_out_12_2_3 = roundReg_12_2_3;
  assign port_state_out_12_2_4 = roundReg_12_2_4;
  assign port_state_out_12_2_5 = roundReg_12_2_5;
  assign port_state_out_12_2_6 = roundReg_12_2_6;
  assign port_state_out_12_2_7 = roundReg_12_2_7;
  assign port_state_out_12_3_0 = roundReg_12_3_0;
  assign port_state_out_12_3_1 = roundReg_12_3_1;
  assign port_state_out_12_3_2 = roundReg_12_3_2;
  assign port_state_out_12_3_3 = roundReg_12_3_3;
  assign port_state_out_12_3_4 = roundReg_12_3_4;
  assign port_state_out_12_3_5 = roundReg_12_3_5;
  assign port_state_out_12_3_6 = roundReg_12_3_6;
  assign port_state_out_12_3_7 = roundReg_12_3_7;
  assign port_state_out_13_0_0 = roundReg_13_0_0;
  assign port_state_out_13_0_1 = roundReg_13_0_1;
  assign port_state_out_13_0_2 = roundReg_13_0_2;
  assign port_state_out_13_0_3 = roundReg_13_0_3;
  assign port_state_out_13_0_4 = roundReg_13_0_4;
  assign port_state_out_13_0_5 = roundReg_13_0_5;
  assign port_state_out_13_0_6 = roundReg_13_0_6;
  assign port_state_out_13_0_7 = roundReg_13_0_7;
  assign port_state_out_13_1_0 = roundReg_13_1_0;
  assign port_state_out_13_1_1 = roundReg_13_1_1;
  assign port_state_out_13_1_2 = roundReg_13_1_2;
  assign port_state_out_13_1_3 = roundReg_13_1_3;
  assign port_state_out_13_1_4 = roundReg_13_1_4;
  assign port_state_out_13_1_5 = roundReg_13_1_5;
  assign port_state_out_13_1_6 = roundReg_13_1_6;
  assign port_state_out_13_1_7 = roundReg_13_1_7;
  assign port_state_out_13_2_0 = roundReg_13_2_0;
  assign port_state_out_13_2_1 = roundReg_13_2_1;
  assign port_state_out_13_2_2 = roundReg_13_2_2;
  assign port_state_out_13_2_3 = roundReg_13_2_3;
  assign port_state_out_13_2_4 = roundReg_13_2_4;
  assign port_state_out_13_2_5 = roundReg_13_2_5;
  assign port_state_out_13_2_6 = roundReg_13_2_6;
  assign port_state_out_13_2_7 = roundReg_13_2_7;
  assign port_state_out_13_3_0 = roundReg_13_3_0;
  assign port_state_out_13_3_1 = roundReg_13_3_1;
  assign port_state_out_13_3_2 = roundReg_13_3_2;
  assign port_state_out_13_3_3 = roundReg_13_3_3;
  assign port_state_out_13_3_4 = roundReg_13_3_4;
  assign port_state_out_13_3_5 = roundReg_13_3_5;
  assign port_state_out_13_3_6 = roundReg_13_3_6;
  assign port_state_out_13_3_7 = roundReg_13_3_7;
  assign port_state_out_14_0_0 = roundReg_14_0_0;
  assign port_state_out_14_0_1 = roundReg_14_0_1;
  assign port_state_out_14_0_2 = roundReg_14_0_2;
  assign port_state_out_14_0_3 = roundReg_14_0_3;
  assign port_state_out_14_0_4 = roundReg_14_0_4;
  assign port_state_out_14_0_5 = roundReg_14_0_5;
  assign port_state_out_14_0_6 = roundReg_14_0_6;
  assign port_state_out_14_0_7 = roundReg_14_0_7;
  assign port_state_out_14_1_0 = roundReg_14_1_0;
  assign port_state_out_14_1_1 = roundReg_14_1_1;
  assign port_state_out_14_1_2 = roundReg_14_1_2;
  assign port_state_out_14_1_3 = roundReg_14_1_3;
  assign port_state_out_14_1_4 = roundReg_14_1_4;
  assign port_state_out_14_1_5 = roundReg_14_1_5;
  assign port_state_out_14_1_6 = roundReg_14_1_6;
  assign port_state_out_14_1_7 = roundReg_14_1_7;
  assign port_state_out_14_2_0 = roundReg_14_2_0;
  assign port_state_out_14_2_1 = roundReg_14_2_1;
  assign port_state_out_14_2_2 = roundReg_14_2_2;
  assign port_state_out_14_2_3 = roundReg_14_2_3;
  assign port_state_out_14_2_4 = roundReg_14_2_4;
  assign port_state_out_14_2_5 = roundReg_14_2_5;
  assign port_state_out_14_2_6 = roundReg_14_2_6;
  assign port_state_out_14_2_7 = roundReg_14_2_7;
  assign port_state_out_14_3_0 = roundReg_14_3_0;
  assign port_state_out_14_3_1 = roundReg_14_3_1;
  assign port_state_out_14_3_2 = roundReg_14_3_2;
  assign port_state_out_14_3_3 = roundReg_14_3_3;
  assign port_state_out_14_3_4 = roundReg_14_3_4;
  assign port_state_out_14_3_5 = roundReg_14_3_5;
  assign port_state_out_14_3_6 = roundReg_14_3_6;
  assign port_state_out_14_3_7 = roundReg_14_3_7;
  assign port_state_out_15_0_0 = roundReg_15_0_0;
  assign port_state_out_15_0_1 = roundReg_15_0_1;
  assign port_state_out_15_0_2 = roundReg_15_0_2;
  assign port_state_out_15_0_3 = roundReg_15_0_3;
  assign port_state_out_15_0_4 = roundReg_15_0_4;
  assign port_state_out_15_0_5 = roundReg_15_0_5;
  assign port_state_out_15_0_6 = roundReg_15_0_6;
  assign port_state_out_15_0_7 = roundReg_15_0_7;
  assign port_state_out_15_1_0 = roundReg_15_1_0;
  assign port_state_out_15_1_1 = roundReg_15_1_1;
  assign port_state_out_15_1_2 = roundReg_15_1_2;
  assign port_state_out_15_1_3 = roundReg_15_1_3;
  assign port_state_out_15_1_4 = roundReg_15_1_4;
  assign port_state_out_15_1_5 = roundReg_15_1_5;
  assign port_state_out_15_1_6 = roundReg_15_1_6;
  assign port_state_out_15_1_7 = roundReg_15_1_7;
  assign port_state_out_15_2_0 = roundReg_15_2_0;
  assign port_state_out_15_2_1 = roundReg_15_2_1;
  assign port_state_out_15_2_2 = roundReg_15_2_2;
  assign port_state_out_15_2_3 = roundReg_15_2_3;
  assign port_state_out_15_2_4 = roundReg_15_2_4;
  assign port_state_out_15_2_5 = roundReg_15_2_5;
  assign port_state_out_15_2_6 = roundReg_15_2_6;
  assign port_state_out_15_2_7 = roundReg_15_2_7;
  assign port_state_out_15_3_0 = roundReg_15_3_0;
  assign port_state_out_15_3_1 = roundReg_15_3_1;
  assign port_state_out_15_3_2 = roundReg_15_3_2;
  assign port_state_out_15_3_3 = roundReg_15_3_3;
  assign port_state_out_15_3_4 = roundReg_15_3_4;
  assign port_state_out_15_3_5 = roundReg_15_3_5;
  assign port_state_out_15_3_6 = roundReg_15_3_6;
  assign port_state_out_15_3_7 = roundReg_15_3_7;
  always @(posedge clk) begin
    roundReg_0_0_0 <= mixColumns_port_state_out_0_0_0;
    roundReg_0_0_1 <= mixColumns_port_state_out_0_0_1;
    roundReg_0_0_2 <= mixColumns_port_state_out_0_0_2;
    roundReg_0_0_3 <= mixColumns_port_state_out_0_0_3;
    roundReg_0_0_4 <= mixColumns_port_state_out_0_0_4;
    roundReg_0_0_5 <= mixColumns_port_state_out_0_0_5;
    roundReg_0_0_6 <= mixColumns_port_state_out_0_0_6;
    roundReg_0_0_7 <= mixColumns_port_state_out_0_0_7;
    roundReg_0_1_0 <= mixColumns_port_state_out_0_1_0;
    roundReg_0_1_1 <= mixColumns_port_state_out_0_1_1;
    roundReg_0_1_2 <= mixColumns_port_state_out_0_1_2;
    roundReg_0_1_3 <= mixColumns_port_state_out_0_1_3;
    roundReg_0_1_4 <= mixColumns_port_state_out_0_1_4;
    roundReg_0_1_5 <= mixColumns_port_state_out_0_1_5;
    roundReg_0_1_6 <= mixColumns_port_state_out_0_1_6;
    roundReg_0_1_7 <= mixColumns_port_state_out_0_1_7;
    roundReg_0_2_0 <= mixColumns_port_state_out_0_2_0;
    roundReg_0_2_1 <= mixColumns_port_state_out_0_2_1;
    roundReg_0_2_2 <= mixColumns_port_state_out_0_2_2;
    roundReg_0_2_3 <= mixColumns_port_state_out_0_2_3;
    roundReg_0_2_4 <= mixColumns_port_state_out_0_2_4;
    roundReg_0_2_5 <= mixColumns_port_state_out_0_2_5;
    roundReg_0_2_6 <= mixColumns_port_state_out_0_2_6;
    roundReg_0_2_7 <= mixColumns_port_state_out_0_2_7;
    roundReg_0_3_0 <= mixColumns_port_state_out_0_3_0;
    roundReg_0_3_1 <= mixColumns_port_state_out_0_3_1;
    roundReg_0_3_2 <= mixColumns_port_state_out_0_3_2;
    roundReg_0_3_3 <= mixColumns_port_state_out_0_3_3;
    roundReg_0_3_4 <= mixColumns_port_state_out_0_3_4;
    roundReg_0_3_5 <= mixColumns_port_state_out_0_3_5;
    roundReg_0_3_6 <= mixColumns_port_state_out_0_3_6;
    roundReg_0_3_7 <= mixColumns_port_state_out_0_3_7;
    roundReg_1_0_0 <= mixColumns_port_state_out_1_0_0;
    roundReg_1_0_1 <= mixColumns_port_state_out_1_0_1;
    roundReg_1_0_2 <= mixColumns_port_state_out_1_0_2;
    roundReg_1_0_3 <= mixColumns_port_state_out_1_0_3;
    roundReg_1_0_4 <= mixColumns_port_state_out_1_0_4;
    roundReg_1_0_5 <= mixColumns_port_state_out_1_0_5;
    roundReg_1_0_6 <= mixColumns_port_state_out_1_0_6;
    roundReg_1_0_7 <= mixColumns_port_state_out_1_0_7;
    roundReg_1_1_0 <= mixColumns_port_state_out_1_1_0;
    roundReg_1_1_1 <= mixColumns_port_state_out_1_1_1;
    roundReg_1_1_2 <= mixColumns_port_state_out_1_1_2;
    roundReg_1_1_3 <= mixColumns_port_state_out_1_1_3;
    roundReg_1_1_4 <= mixColumns_port_state_out_1_1_4;
    roundReg_1_1_5 <= mixColumns_port_state_out_1_1_5;
    roundReg_1_1_6 <= mixColumns_port_state_out_1_1_6;
    roundReg_1_1_7 <= mixColumns_port_state_out_1_1_7;
    roundReg_1_2_0 <= mixColumns_port_state_out_1_2_0;
    roundReg_1_2_1 <= mixColumns_port_state_out_1_2_1;
    roundReg_1_2_2 <= mixColumns_port_state_out_1_2_2;
    roundReg_1_2_3 <= mixColumns_port_state_out_1_2_3;
    roundReg_1_2_4 <= mixColumns_port_state_out_1_2_4;
    roundReg_1_2_5 <= mixColumns_port_state_out_1_2_5;
    roundReg_1_2_6 <= mixColumns_port_state_out_1_2_6;
    roundReg_1_2_7 <= mixColumns_port_state_out_1_2_7;
    roundReg_1_3_0 <= mixColumns_port_state_out_1_3_0;
    roundReg_1_3_1 <= mixColumns_port_state_out_1_3_1;
    roundReg_1_3_2 <= mixColumns_port_state_out_1_3_2;
    roundReg_1_3_3 <= mixColumns_port_state_out_1_3_3;
    roundReg_1_3_4 <= mixColumns_port_state_out_1_3_4;
    roundReg_1_3_5 <= mixColumns_port_state_out_1_3_5;
    roundReg_1_3_6 <= mixColumns_port_state_out_1_3_6;
    roundReg_1_3_7 <= mixColumns_port_state_out_1_3_7;
    roundReg_2_0_0 <= mixColumns_port_state_out_2_0_0;
    roundReg_2_0_1 <= mixColumns_port_state_out_2_0_1;
    roundReg_2_0_2 <= mixColumns_port_state_out_2_0_2;
    roundReg_2_0_3 <= mixColumns_port_state_out_2_0_3;
    roundReg_2_0_4 <= mixColumns_port_state_out_2_0_4;
    roundReg_2_0_5 <= mixColumns_port_state_out_2_0_5;
    roundReg_2_0_6 <= mixColumns_port_state_out_2_0_6;
    roundReg_2_0_7 <= mixColumns_port_state_out_2_0_7;
    roundReg_2_1_0 <= mixColumns_port_state_out_2_1_0;
    roundReg_2_1_1 <= mixColumns_port_state_out_2_1_1;
    roundReg_2_1_2 <= mixColumns_port_state_out_2_1_2;
    roundReg_2_1_3 <= mixColumns_port_state_out_2_1_3;
    roundReg_2_1_4 <= mixColumns_port_state_out_2_1_4;
    roundReg_2_1_5 <= mixColumns_port_state_out_2_1_5;
    roundReg_2_1_6 <= mixColumns_port_state_out_2_1_6;
    roundReg_2_1_7 <= mixColumns_port_state_out_2_1_7;
    roundReg_2_2_0 <= mixColumns_port_state_out_2_2_0;
    roundReg_2_2_1 <= mixColumns_port_state_out_2_2_1;
    roundReg_2_2_2 <= mixColumns_port_state_out_2_2_2;
    roundReg_2_2_3 <= mixColumns_port_state_out_2_2_3;
    roundReg_2_2_4 <= mixColumns_port_state_out_2_2_4;
    roundReg_2_2_5 <= mixColumns_port_state_out_2_2_5;
    roundReg_2_2_6 <= mixColumns_port_state_out_2_2_6;
    roundReg_2_2_7 <= mixColumns_port_state_out_2_2_7;
    roundReg_2_3_0 <= mixColumns_port_state_out_2_3_0;
    roundReg_2_3_1 <= mixColumns_port_state_out_2_3_1;
    roundReg_2_3_2 <= mixColumns_port_state_out_2_3_2;
    roundReg_2_3_3 <= mixColumns_port_state_out_2_3_3;
    roundReg_2_3_4 <= mixColumns_port_state_out_2_3_4;
    roundReg_2_3_5 <= mixColumns_port_state_out_2_3_5;
    roundReg_2_3_6 <= mixColumns_port_state_out_2_3_6;
    roundReg_2_3_7 <= mixColumns_port_state_out_2_3_7;
    roundReg_3_0_0 <= mixColumns_port_state_out_3_0_0;
    roundReg_3_0_1 <= mixColumns_port_state_out_3_0_1;
    roundReg_3_0_2 <= mixColumns_port_state_out_3_0_2;
    roundReg_3_0_3 <= mixColumns_port_state_out_3_0_3;
    roundReg_3_0_4 <= mixColumns_port_state_out_3_0_4;
    roundReg_3_0_5 <= mixColumns_port_state_out_3_0_5;
    roundReg_3_0_6 <= mixColumns_port_state_out_3_0_6;
    roundReg_3_0_7 <= mixColumns_port_state_out_3_0_7;
    roundReg_3_1_0 <= mixColumns_port_state_out_3_1_0;
    roundReg_3_1_1 <= mixColumns_port_state_out_3_1_1;
    roundReg_3_1_2 <= mixColumns_port_state_out_3_1_2;
    roundReg_3_1_3 <= mixColumns_port_state_out_3_1_3;
    roundReg_3_1_4 <= mixColumns_port_state_out_3_1_4;
    roundReg_3_1_5 <= mixColumns_port_state_out_3_1_5;
    roundReg_3_1_6 <= mixColumns_port_state_out_3_1_6;
    roundReg_3_1_7 <= mixColumns_port_state_out_3_1_7;
    roundReg_3_2_0 <= mixColumns_port_state_out_3_2_0;
    roundReg_3_2_1 <= mixColumns_port_state_out_3_2_1;
    roundReg_3_2_2 <= mixColumns_port_state_out_3_2_2;
    roundReg_3_2_3 <= mixColumns_port_state_out_3_2_3;
    roundReg_3_2_4 <= mixColumns_port_state_out_3_2_4;
    roundReg_3_2_5 <= mixColumns_port_state_out_3_2_5;
    roundReg_3_2_6 <= mixColumns_port_state_out_3_2_6;
    roundReg_3_2_7 <= mixColumns_port_state_out_3_2_7;
    roundReg_3_3_0 <= mixColumns_port_state_out_3_3_0;
    roundReg_3_3_1 <= mixColumns_port_state_out_3_3_1;
    roundReg_3_3_2 <= mixColumns_port_state_out_3_3_2;
    roundReg_3_3_3 <= mixColumns_port_state_out_3_3_3;
    roundReg_3_3_4 <= mixColumns_port_state_out_3_3_4;
    roundReg_3_3_5 <= mixColumns_port_state_out_3_3_5;
    roundReg_3_3_6 <= mixColumns_port_state_out_3_3_6;
    roundReg_3_3_7 <= mixColumns_port_state_out_3_3_7;
    roundReg_4_0_0 <= mixColumns_port_state_out_4_0_0;
    roundReg_4_0_1 <= mixColumns_port_state_out_4_0_1;
    roundReg_4_0_2 <= mixColumns_port_state_out_4_0_2;
    roundReg_4_0_3 <= mixColumns_port_state_out_4_0_3;
    roundReg_4_0_4 <= mixColumns_port_state_out_4_0_4;
    roundReg_4_0_5 <= mixColumns_port_state_out_4_0_5;
    roundReg_4_0_6 <= mixColumns_port_state_out_4_0_6;
    roundReg_4_0_7 <= mixColumns_port_state_out_4_0_7;
    roundReg_4_1_0 <= mixColumns_port_state_out_4_1_0;
    roundReg_4_1_1 <= mixColumns_port_state_out_4_1_1;
    roundReg_4_1_2 <= mixColumns_port_state_out_4_1_2;
    roundReg_4_1_3 <= mixColumns_port_state_out_4_1_3;
    roundReg_4_1_4 <= mixColumns_port_state_out_4_1_4;
    roundReg_4_1_5 <= mixColumns_port_state_out_4_1_5;
    roundReg_4_1_6 <= mixColumns_port_state_out_4_1_6;
    roundReg_4_1_7 <= mixColumns_port_state_out_4_1_7;
    roundReg_4_2_0 <= mixColumns_port_state_out_4_2_0;
    roundReg_4_2_1 <= mixColumns_port_state_out_4_2_1;
    roundReg_4_2_2 <= mixColumns_port_state_out_4_2_2;
    roundReg_4_2_3 <= mixColumns_port_state_out_4_2_3;
    roundReg_4_2_4 <= mixColumns_port_state_out_4_2_4;
    roundReg_4_2_5 <= mixColumns_port_state_out_4_2_5;
    roundReg_4_2_6 <= mixColumns_port_state_out_4_2_6;
    roundReg_4_2_7 <= mixColumns_port_state_out_4_2_7;
    roundReg_4_3_0 <= mixColumns_port_state_out_4_3_0;
    roundReg_4_3_1 <= mixColumns_port_state_out_4_3_1;
    roundReg_4_3_2 <= mixColumns_port_state_out_4_3_2;
    roundReg_4_3_3 <= mixColumns_port_state_out_4_3_3;
    roundReg_4_3_4 <= mixColumns_port_state_out_4_3_4;
    roundReg_4_3_5 <= mixColumns_port_state_out_4_3_5;
    roundReg_4_3_6 <= mixColumns_port_state_out_4_3_6;
    roundReg_4_3_7 <= mixColumns_port_state_out_4_3_7;
    roundReg_5_0_0 <= mixColumns_port_state_out_5_0_0;
    roundReg_5_0_1 <= mixColumns_port_state_out_5_0_1;
    roundReg_5_0_2 <= mixColumns_port_state_out_5_0_2;
    roundReg_5_0_3 <= mixColumns_port_state_out_5_0_3;
    roundReg_5_0_4 <= mixColumns_port_state_out_5_0_4;
    roundReg_5_0_5 <= mixColumns_port_state_out_5_0_5;
    roundReg_5_0_6 <= mixColumns_port_state_out_5_0_6;
    roundReg_5_0_7 <= mixColumns_port_state_out_5_0_7;
    roundReg_5_1_0 <= mixColumns_port_state_out_5_1_0;
    roundReg_5_1_1 <= mixColumns_port_state_out_5_1_1;
    roundReg_5_1_2 <= mixColumns_port_state_out_5_1_2;
    roundReg_5_1_3 <= mixColumns_port_state_out_5_1_3;
    roundReg_5_1_4 <= mixColumns_port_state_out_5_1_4;
    roundReg_5_1_5 <= mixColumns_port_state_out_5_1_5;
    roundReg_5_1_6 <= mixColumns_port_state_out_5_1_6;
    roundReg_5_1_7 <= mixColumns_port_state_out_5_1_7;
    roundReg_5_2_0 <= mixColumns_port_state_out_5_2_0;
    roundReg_5_2_1 <= mixColumns_port_state_out_5_2_1;
    roundReg_5_2_2 <= mixColumns_port_state_out_5_2_2;
    roundReg_5_2_3 <= mixColumns_port_state_out_5_2_3;
    roundReg_5_2_4 <= mixColumns_port_state_out_5_2_4;
    roundReg_5_2_5 <= mixColumns_port_state_out_5_2_5;
    roundReg_5_2_6 <= mixColumns_port_state_out_5_2_6;
    roundReg_5_2_7 <= mixColumns_port_state_out_5_2_7;
    roundReg_5_3_0 <= mixColumns_port_state_out_5_3_0;
    roundReg_5_3_1 <= mixColumns_port_state_out_5_3_1;
    roundReg_5_3_2 <= mixColumns_port_state_out_5_3_2;
    roundReg_5_3_3 <= mixColumns_port_state_out_5_3_3;
    roundReg_5_3_4 <= mixColumns_port_state_out_5_3_4;
    roundReg_5_3_5 <= mixColumns_port_state_out_5_3_5;
    roundReg_5_3_6 <= mixColumns_port_state_out_5_3_6;
    roundReg_5_3_7 <= mixColumns_port_state_out_5_3_7;
    roundReg_6_0_0 <= mixColumns_port_state_out_6_0_0;
    roundReg_6_0_1 <= mixColumns_port_state_out_6_0_1;
    roundReg_6_0_2 <= mixColumns_port_state_out_6_0_2;
    roundReg_6_0_3 <= mixColumns_port_state_out_6_0_3;
    roundReg_6_0_4 <= mixColumns_port_state_out_6_0_4;
    roundReg_6_0_5 <= mixColumns_port_state_out_6_0_5;
    roundReg_6_0_6 <= mixColumns_port_state_out_6_0_6;
    roundReg_6_0_7 <= mixColumns_port_state_out_6_0_7;
    roundReg_6_1_0 <= mixColumns_port_state_out_6_1_0;
    roundReg_6_1_1 <= mixColumns_port_state_out_6_1_1;
    roundReg_6_1_2 <= mixColumns_port_state_out_6_1_2;
    roundReg_6_1_3 <= mixColumns_port_state_out_6_1_3;
    roundReg_6_1_4 <= mixColumns_port_state_out_6_1_4;
    roundReg_6_1_5 <= mixColumns_port_state_out_6_1_5;
    roundReg_6_1_6 <= mixColumns_port_state_out_6_1_6;
    roundReg_6_1_7 <= mixColumns_port_state_out_6_1_7;
    roundReg_6_2_0 <= mixColumns_port_state_out_6_2_0;
    roundReg_6_2_1 <= mixColumns_port_state_out_6_2_1;
    roundReg_6_2_2 <= mixColumns_port_state_out_6_2_2;
    roundReg_6_2_3 <= mixColumns_port_state_out_6_2_3;
    roundReg_6_2_4 <= mixColumns_port_state_out_6_2_4;
    roundReg_6_2_5 <= mixColumns_port_state_out_6_2_5;
    roundReg_6_2_6 <= mixColumns_port_state_out_6_2_6;
    roundReg_6_2_7 <= mixColumns_port_state_out_6_2_7;
    roundReg_6_3_0 <= mixColumns_port_state_out_6_3_0;
    roundReg_6_3_1 <= mixColumns_port_state_out_6_3_1;
    roundReg_6_3_2 <= mixColumns_port_state_out_6_3_2;
    roundReg_6_3_3 <= mixColumns_port_state_out_6_3_3;
    roundReg_6_3_4 <= mixColumns_port_state_out_6_3_4;
    roundReg_6_3_5 <= mixColumns_port_state_out_6_3_5;
    roundReg_6_3_6 <= mixColumns_port_state_out_6_3_6;
    roundReg_6_3_7 <= mixColumns_port_state_out_6_3_7;
    roundReg_7_0_0 <= mixColumns_port_state_out_7_0_0;
    roundReg_7_0_1 <= mixColumns_port_state_out_7_0_1;
    roundReg_7_0_2 <= mixColumns_port_state_out_7_0_2;
    roundReg_7_0_3 <= mixColumns_port_state_out_7_0_3;
    roundReg_7_0_4 <= mixColumns_port_state_out_7_0_4;
    roundReg_7_0_5 <= mixColumns_port_state_out_7_0_5;
    roundReg_7_0_6 <= mixColumns_port_state_out_7_0_6;
    roundReg_7_0_7 <= mixColumns_port_state_out_7_0_7;
    roundReg_7_1_0 <= mixColumns_port_state_out_7_1_0;
    roundReg_7_1_1 <= mixColumns_port_state_out_7_1_1;
    roundReg_7_1_2 <= mixColumns_port_state_out_7_1_2;
    roundReg_7_1_3 <= mixColumns_port_state_out_7_1_3;
    roundReg_7_1_4 <= mixColumns_port_state_out_7_1_4;
    roundReg_7_1_5 <= mixColumns_port_state_out_7_1_5;
    roundReg_7_1_6 <= mixColumns_port_state_out_7_1_6;
    roundReg_7_1_7 <= mixColumns_port_state_out_7_1_7;
    roundReg_7_2_0 <= mixColumns_port_state_out_7_2_0;
    roundReg_7_2_1 <= mixColumns_port_state_out_7_2_1;
    roundReg_7_2_2 <= mixColumns_port_state_out_7_2_2;
    roundReg_7_2_3 <= mixColumns_port_state_out_7_2_3;
    roundReg_7_2_4 <= mixColumns_port_state_out_7_2_4;
    roundReg_7_2_5 <= mixColumns_port_state_out_7_2_5;
    roundReg_7_2_6 <= mixColumns_port_state_out_7_2_6;
    roundReg_7_2_7 <= mixColumns_port_state_out_7_2_7;
    roundReg_7_3_0 <= mixColumns_port_state_out_7_3_0;
    roundReg_7_3_1 <= mixColumns_port_state_out_7_3_1;
    roundReg_7_3_2 <= mixColumns_port_state_out_7_3_2;
    roundReg_7_3_3 <= mixColumns_port_state_out_7_3_3;
    roundReg_7_3_4 <= mixColumns_port_state_out_7_3_4;
    roundReg_7_3_5 <= mixColumns_port_state_out_7_3_5;
    roundReg_7_3_6 <= mixColumns_port_state_out_7_3_6;
    roundReg_7_3_7 <= mixColumns_port_state_out_7_3_7;
    roundReg_8_0_0 <= mixColumns_port_state_out_8_0_0;
    roundReg_8_0_1 <= mixColumns_port_state_out_8_0_1;
    roundReg_8_0_2 <= mixColumns_port_state_out_8_0_2;
    roundReg_8_0_3 <= mixColumns_port_state_out_8_0_3;
    roundReg_8_0_4 <= mixColumns_port_state_out_8_0_4;
    roundReg_8_0_5 <= mixColumns_port_state_out_8_0_5;
    roundReg_8_0_6 <= mixColumns_port_state_out_8_0_6;
    roundReg_8_0_7 <= mixColumns_port_state_out_8_0_7;
    roundReg_8_1_0 <= mixColumns_port_state_out_8_1_0;
    roundReg_8_1_1 <= mixColumns_port_state_out_8_1_1;
    roundReg_8_1_2 <= mixColumns_port_state_out_8_1_2;
    roundReg_8_1_3 <= mixColumns_port_state_out_8_1_3;
    roundReg_8_1_4 <= mixColumns_port_state_out_8_1_4;
    roundReg_8_1_5 <= mixColumns_port_state_out_8_1_5;
    roundReg_8_1_6 <= mixColumns_port_state_out_8_1_6;
    roundReg_8_1_7 <= mixColumns_port_state_out_8_1_7;
    roundReg_8_2_0 <= mixColumns_port_state_out_8_2_0;
    roundReg_8_2_1 <= mixColumns_port_state_out_8_2_1;
    roundReg_8_2_2 <= mixColumns_port_state_out_8_2_2;
    roundReg_8_2_3 <= mixColumns_port_state_out_8_2_3;
    roundReg_8_2_4 <= mixColumns_port_state_out_8_2_4;
    roundReg_8_2_5 <= mixColumns_port_state_out_8_2_5;
    roundReg_8_2_6 <= mixColumns_port_state_out_8_2_6;
    roundReg_8_2_7 <= mixColumns_port_state_out_8_2_7;
    roundReg_8_3_0 <= mixColumns_port_state_out_8_3_0;
    roundReg_8_3_1 <= mixColumns_port_state_out_8_3_1;
    roundReg_8_3_2 <= mixColumns_port_state_out_8_3_2;
    roundReg_8_3_3 <= mixColumns_port_state_out_8_3_3;
    roundReg_8_3_4 <= mixColumns_port_state_out_8_3_4;
    roundReg_8_3_5 <= mixColumns_port_state_out_8_3_5;
    roundReg_8_3_6 <= mixColumns_port_state_out_8_3_6;
    roundReg_8_3_7 <= mixColumns_port_state_out_8_3_7;
    roundReg_9_0_0 <= mixColumns_port_state_out_9_0_0;
    roundReg_9_0_1 <= mixColumns_port_state_out_9_0_1;
    roundReg_9_0_2 <= mixColumns_port_state_out_9_0_2;
    roundReg_9_0_3 <= mixColumns_port_state_out_9_0_3;
    roundReg_9_0_4 <= mixColumns_port_state_out_9_0_4;
    roundReg_9_0_5 <= mixColumns_port_state_out_9_0_5;
    roundReg_9_0_6 <= mixColumns_port_state_out_9_0_6;
    roundReg_9_0_7 <= mixColumns_port_state_out_9_0_7;
    roundReg_9_1_0 <= mixColumns_port_state_out_9_1_0;
    roundReg_9_1_1 <= mixColumns_port_state_out_9_1_1;
    roundReg_9_1_2 <= mixColumns_port_state_out_9_1_2;
    roundReg_9_1_3 <= mixColumns_port_state_out_9_1_3;
    roundReg_9_1_4 <= mixColumns_port_state_out_9_1_4;
    roundReg_9_1_5 <= mixColumns_port_state_out_9_1_5;
    roundReg_9_1_6 <= mixColumns_port_state_out_9_1_6;
    roundReg_9_1_7 <= mixColumns_port_state_out_9_1_7;
    roundReg_9_2_0 <= mixColumns_port_state_out_9_2_0;
    roundReg_9_2_1 <= mixColumns_port_state_out_9_2_1;
    roundReg_9_2_2 <= mixColumns_port_state_out_9_2_2;
    roundReg_9_2_3 <= mixColumns_port_state_out_9_2_3;
    roundReg_9_2_4 <= mixColumns_port_state_out_9_2_4;
    roundReg_9_2_5 <= mixColumns_port_state_out_9_2_5;
    roundReg_9_2_6 <= mixColumns_port_state_out_9_2_6;
    roundReg_9_2_7 <= mixColumns_port_state_out_9_2_7;
    roundReg_9_3_0 <= mixColumns_port_state_out_9_3_0;
    roundReg_9_3_1 <= mixColumns_port_state_out_9_3_1;
    roundReg_9_3_2 <= mixColumns_port_state_out_9_3_2;
    roundReg_9_3_3 <= mixColumns_port_state_out_9_3_3;
    roundReg_9_3_4 <= mixColumns_port_state_out_9_3_4;
    roundReg_9_3_5 <= mixColumns_port_state_out_9_3_5;
    roundReg_9_3_6 <= mixColumns_port_state_out_9_3_6;
    roundReg_9_3_7 <= mixColumns_port_state_out_9_3_7;
    roundReg_10_0_0 <= mixColumns_port_state_out_10_0_0;
    roundReg_10_0_1 <= mixColumns_port_state_out_10_0_1;
    roundReg_10_0_2 <= mixColumns_port_state_out_10_0_2;
    roundReg_10_0_3 <= mixColumns_port_state_out_10_0_3;
    roundReg_10_0_4 <= mixColumns_port_state_out_10_0_4;
    roundReg_10_0_5 <= mixColumns_port_state_out_10_0_5;
    roundReg_10_0_6 <= mixColumns_port_state_out_10_0_6;
    roundReg_10_0_7 <= mixColumns_port_state_out_10_0_7;
    roundReg_10_1_0 <= mixColumns_port_state_out_10_1_0;
    roundReg_10_1_1 <= mixColumns_port_state_out_10_1_1;
    roundReg_10_1_2 <= mixColumns_port_state_out_10_1_2;
    roundReg_10_1_3 <= mixColumns_port_state_out_10_1_3;
    roundReg_10_1_4 <= mixColumns_port_state_out_10_1_4;
    roundReg_10_1_5 <= mixColumns_port_state_out_10_1_5;
    roundReg_10_1_6 <= mixColumns_port_state_out_10_1_6;
    roundReg_10_1_7 <= mixColumns_port_state_out_10_1_7;
    roundReg_10_2_0 <= mixColumns_port_state_out_10_2_0;
    roundReg_10_2_1 <= mixColumns_port_state_out_10_2_1;
    roundReg_10_2_2 <= mixColumns_port_state_out_10_2_2;
    roundReg_10_2_3 <= mixColumns_port_state_out_10_2_3;
    roundReg_10_2_4 <= mixColumns_port_state_out_10_2_4;
    roundReg_10_2_5 <= mixColumns_port_state_out_10_2_5;
    roundReg_10_2_6 <= mixColumns_port_state_out_10_2_6;
    roundReg_10_2_7 <= mixColumns_port_state_out_10_2_7;
    roundReg_10_3_0 <= mixColumns_port_state_out_10_3_0;
    roundReg_10_3_1 <= mixColumns_port_state_out_10_3_1;
    roundReg_10_3_2 <= mixColumns_port_state_out_10_3_2;
    roundReg_10_3_3 <= mixColumns_port_state_out_10_3_3;
    roundReg_10_3_4 <= mixColumns_port_state_out_10_3_4;
    roundReg_10_3_5 <= mixColumns_port_state_out_10_3_5;
    roundReg_10_3_6 <= mixColumns_port_state_out_10_3_6;
    roundReg_10_3_7 <= mixColumns_port_state_out_10_3_7;
    roundReg_11_0_0 <= mixColumns_port_state_out_11_0_0;
    roundReg_11_0_1 <= mixColumns_port_state_out_11_0_1;
    roundReg_11_0_2 <= mixColumns_port_state_out_11_0_2;
    roundReg_11_0_3 <= mixColumns_port_state_out_11_0_3;
    roundReg_11_0_4 <= mixColumns_port_state_out_11_0_4;
    roundReg_11_0_5 <= mixColumns_port_state_out_11_0_5;
    roundReg_11_0_6 <= mixColumns_port_state_out_11_0_6;
    roundReg_11_0_7 <= mixColumns_port_state_out_11_0_7;
    roundReg_11_1_0 <= mixColumns_port_state_out_11_1_0;
    roundReg_11_1_1 <= mixColumns_port_state_out_11_1_1;
    roundReg_11_1_2 <= mixColumns_port_state_out_11_1_2;
    roundReg_11_1_3 <= mixColumns_port_state_out_11_1_3;
    roundReg_11_1_4 <= mixColumns_port_state_out_11_1_4;
    roundReg_11_1_5 <= mixColumns_port_state_out_11_1_5;
    roundReg_11_1_6 <= mixColumns_port_state_out_11_1_6;
    roundReg_11_1_7 <= mixColumns_port_state_out_11_1_7;
    roundReg_11_2_0 <= mixColumns_port_state_out_11_2_0;
    roundReg_11_2_1 <= mixColumns_port_state_out_11_2_1;
    roundReg_11_2_2 <= mixColumns_port_state_out_11_2_2;
    roundReg_11_2_3 <= mixColumns_port_state_out_11_2_3;
    roundReg_11_2_4 <= mixColumns_port_state_out_11_2_4;
    roundReg_11_2_5 <= mixColumns_port_state_out_11_2_5;
    roundReg_11_2_6 <= mixColumns_port_state_out_11_2_6;
    roundReg_11_2_7 <= mixColumns_port_state_out_11_2_7;
    roundReg_11_3_0 <= mixColumns_port_state_out_11_3_0;
    roundReg_11_3_1 <= mixColumns_port_state_out_11_3_1;
    roundReg_11_3_2 <= mixColumns_port_state_out_11_3_2;
    roundReg_11_3_3 <= mixColumns_port_state_out_11_3_3;
    roundReg_11_3_4 <= mixColumns_port_state_out_11_3_4;
    roundReg_11_3_5 <= mixColumns_port_state_out_11_3_5;
    roundReg_11_3_6 <= mixColumns_port_state_out_11_3_6;
    roundReg_11_3_7 <= mixColumns_port_state_out_11_3_7;
    roundReg_12_0_0 <= mixColumns_port_state_out_12_0_0;
    roundReg_12_0_1 <= mixColumns_port_state_out_12_0_1;
    roundReg_12_0_2 <= mixColumns_port_state_out_12_0_2;
    roundReg_12_0_3 <= mixColumns_port_state_out_12_0_3;
    roundReg_12_0_4 <= mixColumns_port_state_out_12_0_4;
    roundReg_12_0_5 <= mixColumns_port_state_out_12_0_5;
    roundReg_12_0_6 <= mixColumns_port_state_out_12_0_6;
    roundReg_12_0_7 <= mixColumns_port_state_out_12_0_7;
    roundReg_12_1_0 <= mixColumns_port_state_out_12_1_0;
    roundReg_12_1_1 <= mixColumns_port_state_out_12_1_1;
    roundReg_12_1_2 <= mixColumns_port_state_out_12_1_2;
    roundReg_12_1_3 <= mixColumns_port_state_out_12_1_3;
    roundReg_12_1_4 <= mixColumns_port_state_out_12_1_4;
    roundReg_12_1_5 <= mixColumns_port_state_out_12_1_5;
    roundReg_12_1_6 <= mixColumns_port_state_out_12_1_6;
    roundReg_12_1_7 <= mixColumns_port_state_out_12_1_7;
    roundReg_12_2_0 <= mixColumns_port_state_out_12_2_0;
    roundReg_12_2_1 <= mixColumns_port_state_out_12_2_1;
    roundReg_12_2_2 <= mixColumns_port_state_out_12_2_2;
    roundReg_12_2_3 <= mixColumns_port_state_out_12_2_3;
    roundReg_12_2_4 <= mixColumns_port_state_out_12_2_4;
    roundReg_12_2_5 <= mixColumns_port_state_out_12_2_5;
    roundReg_12_2_6 <= mixColumns_port_state_out_12_2_6;
    roundReg_12_2_7 <= mixColumns_port_state_out_12_2_7;
    roundReg_12_3_0 <= mixColumns_port_state_out_12_3_0;
    roundReg_12_3_1 <= mixColumns_port_state_out_12_3_1;
    roundReg_12_3_2 <= mixColumns_port_state_out_12_3_2;
    roundReg_12_3_3 <= mixColumns_port_state_out_12_3_3;
    roundReg_12_3_4 <= mixColumns_port_state_out_12_3_4;
    roundReg_12_3_5 <= mixColumns_port_state_out_12_3_5;
    roundReg_12_3_6 <= mixColumns_port_state_out_12_3_6;
    roundReg_12_3_7 <= mixColumns_port_state_out_12_3_7;
    roundReg_13_0_0 <= mixColumns_port_state_out_13_0_0;
    roundReg_13_0_1 <= mixColumns_port_state_out_13_0_1;
    roundReg_13_0_2 <= mixColumns_port_state_out_13_0_2;
    roundReg_13_0_3 <= mixColumns_port_state_out_13_0_3;
    roundReg_13_0_4 <= mixColumns_port_state_out_13_0_4;
    roundReg_13_0_5 <= mixColumns_port_state_out_13_0_5;
    roundReg_13_0_6 <= mixColumns_port_state_out_13_0_6;
    roundReg_13_0_7 <= mixColumns_port_state_out_13_0_7;
    roundReg_13_1_0 <= mixColumns_port_state_out_13_1_0;
    roundReg_13_1_1 <= mixColumns_port_state_out_13_1_1;
    roundReg_13_1_2 <= mixColumns_port_state_out_13_1_2;
    roundReg_13_1_3 <= mixColumns_port_state_out_13_1_3;
    roundReg_13_1_4 <= mixColumns_port_state_out_13_1_4;
    roundReg_13_1_5 <= mixColumns_port_state_out_13_1_5;
    roundReg_13_1_6 <= mixColumns_port_state_out_13_1_6;
    roundReg_13_1_7 <= mixColumns_port_state_out_13_1_7;
    roundReg_13_2_0 <= mixColumns_port_state_out_13_2_0;
    roundReg_13_2_1 <= mixColumns_port_state_out_13_2_1;
    roundReg_13_2_2 <= mixColumns_port_state_out_13_2_2;
    roundReg_13_2_3 <= mixColumns_port_state_out_13_2_3;
    roundReg_13_2_4 <= mixColumns_port_state_out_13_2_4;
    roundReg_13_2_5 <= mixColumns_port_state_out_13_2_5;
    roundReg_13_2_6 <= mixColumns_port_state_out_13_2_6;
    roundReg_13_2_7 <= mixColumns_port_state_out_13_2_7;
    roundReg_13_3_0 <= mixColumns_port_state_out_13_3_0;
    roundReg_13_3_1 <= mixColumns_port_state_out_13_3_1;
    roundReg_13_3_2 <= mixColumns_port_state_out_13_3_2;
    roundReg_13_3_3 <= mixColumns_port_state_out_13_3_3;
    roundReg_13_3_4 <= mixColumns_port_state_out_13_3_4;
    roundReg_13_3_5 <= mixColumns_port_state_out_13_3_5;
    roundReg_13_3_6 <= mixColumns_port_state_out_13_3_6;
    roundReg_13_3_7 <= mixColumns_port_state_out_13_3_7;
    roundReg_14_0_0 <= mixColumns_port_state_out_14_0_0;
    roundReg_14_0_1 <= mixColumns_port_state_out_14_0_1;
    roundReg_14_0_2 <= mixColumns_port_state_out_14_0_2;
    roundReg_14_0_3 <= mixColumns_port_state_out_14_0_3;
    roundReg_14_0_4 <= mixColumns_port_state_out_14_0_4;
    roundReg_14_0_5 <= mixColumns_port_state_out_14_0_5;
    roundReg_14_0_6 <= mixColumns_port_state_out_14_0_6;
    roundReg_14_0_7 <= mixColumns_port_state_out_14_0_7;
    roundReg_14_1_0 <= mixColumns_port_state_out_14_1_0;
    roundReg_14_1_1 <= mixColumns_port_state_out_14_1_1;
    roundReg_14_1_2 <= mixColumns_port_state_out_14_1_2;
    roundReg_14_1_3 <= mixColumns_port_state_out_14_1_3;
    roundReg_14_1_4 <= mixColumns_port_state_out_14_1_4;
    roundReg_14_1_5 <= mixColumns_port_state_out_14_1_5;
    roundReg_14_1_6 <= mixColumns_port_state_out_14_1_6;
    roundReg_14_1_7 <= mixColumns_port_state_out_14_1_7;
    roundReg_14_2_0 <= mixColumns_port_state_out_14_2_0;
    roundReg_14_2_1 <= mixColumns_port_state_out_14_2_1;
    roundReg_14_2_2 <= mixColumns_port_state_out_14_2_2;
    roundReg_14_2_3 <= mixColumns_port_state_out_14_2_3;
    roundReg_14_2_4 <= mixColumns_port_state_out_14_2_4;
    roundReg_14_2_5 <= mixColumns_port_state_out_14_2_5;
    roundReg_14_2_6 <= mixColumns_port_state_out_14_2_6;
    roundReg_14_2_7 <= mixColumns_port_state_out_14_2_7;
    roundReg_14_3_0 <= mixColumns_port_state_out_14_3_0;
    roundReg_14_3_1 <= mixColumns_port_state_out_14_3_1;
    roundReg_14_3_2 <= mixColumns_port_state_out_14_3_2;
    roundReg_14_3_3 <= mixColumns_port_state_out_14_3_3;
    roundReg_14_3_4 <= mixColumns_port_state_out_14_3_4;
    roundReg_14_3_5 <= mixColumns_port_state_out_14_3_5;
    roundReg_14_3_6 <= mixColumns_port_state_out_14_3_6;
    roundReg_14_3_7 <= mixColumns_port_state_out_14_3_7;
    roundReg_15_0_0 <= mixColumns_port_state_out_15_0_0;
    roundReg_15_0_1 <= mixColumns_port_state_out_15_0_1;
    roundReg_15_0_2 <= mixColumns_port_state_out_15_0_2;
    roundReg_15_0_3 <= mixColumns_port_state_out_15_0_3;
    roundReg_15_0_4 <= mixColumns_port_state_out_15_0_4;
    roundReg_15_0_5 <= mixColumns_port_state_out_15_0_5;
    roundReg_15_0_6 <= mixColumns_port_state_out_15_0_6;
    roundReg_15_0_7 <= mixColumns_port_state_out_15_0_7;
    roundReg_15_1_0 <= mixColumns_port_state_out_15_1_0;
    roundReg_15_1_1 <= mixColumns_port_state_out_15_1_1;
    roundReg_15_1_2 <= mixColumns_port_state_out_15_1_2;
    roundReg_15_1_3 <= mixColumns_port_state_out_15_1_3;
    roundReg_15_1_4 <= mixColumns_port_state_out_15_1_4;
    roundReg_15_1_5 <= mixColumns_port_state_out_15_1_5;
    roundReg_15_1_6 <= mixColumns_port_state_out_15_1_6;
    roundReg_15_1_7 <= mixColumns_port_state_out_15_1_7;
    roundReg_15_2_0 <= mixColumns_port_state_out_15_2_0;
    roundReg_15_2_1 <= mixColumns_port_state_out_15_2_1;
    roundReg_15_2_2 <= mixColumns_port_state_out_15_2_2;
    roundReg_15_2_3 <= mixColumns_port_state_out_15_2_3;
    roundReg_15_2_4 <= mixColumns_port_state_out_15_2_4;
    roundReg_15_2_5 <= mixColumns_port_state_out_15_2_5;
    roundReg_15_2_6 <= mixColumns_port_state_out_15_2_6;
    roundReg_15_2_7 <= mixColumns_port_state_out_15_2_7;
    roundReg_15_3_0 <= mixColumns_port_state_out_15_3_0;
    roundReg_15_3_1 <= mixColumns_port_state_out_15_3_1;
    roundReg_15_3_2 <= mixColumns_port_state_out_15_3_2;
    roundReg_15_3_3 <= mixColumns_port_state_out_15_3_3;
    roundReg_15_3_4 <= mixColumns_port_state_out_15_3_4;
    roundReg_15_3_5 <= mixColumns_port_state_out_15_3_5;
    roundReg_15_3_6 <= mixColumns_port_state_out_15_3_6;
    roundReg_15_3_7 <= mixColumns_port_state_out_15_3_7;
  end


endmodule

module Aes_MixColumn (
  input      [0:0]    port_state_in_0_0_0,
  input      [0:0]    port_state_in_0_0_1,
  input      [0:0]    port_state_in_0_0_2,
  input      [0:0]    port_state_in_0_0_3,
  input      [0:0]    port_state_in_0_0_4,
  input      [0:0]    port_state_in_0_0_5,
  input      [0:0]    port_state_in_0_0_6,
  input      [0:0]    port_state_in_0_0_7,
  input      [0:0]    port_state_in_0_1_0,
  input      [0:0]    port_state_in_0_1_1,
  input      [0:0]    port_state_in_0_1_2,
  input      [0:0]    port_state_in_0_1_3,
  input      [0:0]    port_state_in_0_1_4,
  input      [0:0]    port_state_in_0_1_5,
  input      [0:0]    port_state_in_0_1_6,
  input      [0:0]    port_state_in_0_1_7,
  input      [0:0]    port_state_in_0_2_0,
  input      [0:0]    port_state_in_0_2_1,
  input      [0:0]    port_state_in_0_2_2,
  input      [0:0]    port_state_in_0_2_3,
  input      [0:0]    port_state_in_0_2_4,
  input      [0:0]    port_state_in_0_2_5,
  input      [0:0]    port_state_in_0_2_6,
  input      [0:0]    port_state_in_0_2_7,
  input      [0:0]    port_state_in_0_3_0,
  input      [0:0]    port_state_in_0_3_1,
  input      [0:0]    port_state_in_0_3_2,
  input      [0:0]    port_state_in_0_3_3,
  input      [0:0]    port_state_in_0_3_4,
  input      [0:0]    port_state_in_0_3_5,
  input      [0:0]    port_state_in_0_3_6,
  input      [0:0]    port_state_in_0_3_7,
  input      [0:0]    port_state_in_1_0_0,
  input      [0:0]    port_state_in_1_0_1,
  input      [0:0]    port_state_in_1_0_2,
  input      [0:0]    port_state_in_1_0_3,
  input      [0:0]    port_state_in_1_0_4,
  input      [0:0]    port_state_in_1_0_5,
  input      [0:0]    port_state_in_1_0_6,
  input      [0:0]    port_state_in_1_0_7,
  input      [0:0]    port_state_in_1_1_0,
  input      [0:0]    port_state_in_1_1_1,
  input      [0:0]    port_state_in_1_1_2,
  input      [0:0]    port_state_in_1_1_3,
  input      [0:0]    port_state_in_1_1_4,
  input      [0:0]    port_state_in_1_1_5,
  input      [0:0]    port_state_in_1_1_6,
  input      [0:0]    port_state_in_1_1_7,
  input      [0:0]    port_state_in_1_2_0,
  input      [0:0]    port_state_in_1_2_1,
  input      [0:0]    port_state_in_1_2_2,
  input      [0:0]    port_state_in_1_2_3,
  input      [0:0]    port_state_in_1_2_4,
  input      [0:0]    port_state_in_1_2_5,
  input      [0:0]    port_state_in_1_2_6,
  input      [0:0]    port_state_in_1_2_7,
  input      [0:0]    port_state_in_1_3_0,
  input      [0:0]    port_state_in_1_3_1,
  input      [0:0]    port_state_in_1_3_2,
  input      [0:0]    port_state_in_1_3_3,
  input      [0:0]    port_state_in_1_3_4,
  input      [0:0]    port_state_in_1_3_5,
  input      [0:0]    port_state_in_1_3_6,
  input      [0:0]    port_state_in_1_3_7,
  input      [0:0]    port_state_in_2_0_0,
  input      [0:0]    port_state_in_2_0_1,
  input      [0:0]    port_state_in_2_0_2,
  input      [0:0]    port_state_in_2_0_3,
  input      [0:0]    port_state_in_2_0_4,
  input      [0:0]    port_state_in_2_0_5,
  input      [0:0]    port_state_in_2_0_6,
  input      [0:0]    port_state_in_2_0_7,
  input      [0:0]    port_state_in_2_1_0,
  input      [0:0]    port_state_in_2_1_1,
  input      [0:0]    port_state_in_2_1_2,
  input      [0:0]    port_state_in_2_1_3,
  input      [0:0]    port_state_in_2_1_4,
  input      [0:0]    port_state_in_2_1_5,
  input      [0:0]    port_state_in_2_1_6,
  input      [0:0]    port_state_in_2_1_7,
  input      [0:0]    port_state_in_2_2_0,
  input      [0:0]    port_state_in_2_2_1,
  input      [0:0]    port_state_in_2_2_2,
  input      [0:0]    port_state_in_2_2_3,
  input      [0:0]    port_state_in_2_2_4,
  input      [0:0]    port_state_in_2_2_5,
  input      [0:0]    port_state_in_2_2_6,
  input      [0:0]    port_state_in_2_2_7,
  input      [0:0]    port_state_in_2_3_0,
  input      [0:0]    port_state_in_2_3_1,
  input      [0:0]    port_state_in_2_3_2,
  input      [0:0]    port_state_in_2_3_3,
  input      [0:0]    port_state_in_2_3_4,
  input      [0:0]    port_state_in_2_3_5,
  input      [0:0]    port_state_in_2_3_6,
  input      [0:0]    port_state_in_2_3_7,
  input      [0:0]    port_state_in_3_0_0,
  input      [0:0]    port_state_in_3_0_1,
  input      [0:0]    port_state_in_3_0_2,
  input      [0:0]    port_state_in_3_0_3,
  input      [0:0]    port_state_in_3_0_4,
  input      [0:0]    port_state_in_3_0_5,
  input      [0:0]    port_state_in_3_0_6,
  input      [0:0]    port_state_in_3_0_7,
  input      [0:0]    port_state_in_3_1_0,
  input      [0:0]    port_state_in_3_1_1,
  input      [0:0]    port_state_in_3_1_2,
  input      [0:0]    port_state_in_3_1_3,
  input      [0:0]    port_state_in_3_1_4,
  input      [0:0]    port_state_in_3_1_5,
  input      [0:0]    port_state_in_3_1_6,
  input      [0:0]    port_state_in_3_1_7,
  input      [0:0]    port_state_in_3_2_0,
  input      [0:0]    port_state_in_3_2_1,
  input      [0:0]    port_state_in_3_2_2,
  input      [0:0]    port_state_in_3_2_3,
  input      [0:0]    port_state_in_3_2_4,
  input      [0:0]    port_state_in_3_2_5,
  input      [0:0]    port_state_in_3_2_6,
  input      [0:0]    port_state_in_3_2_7,
  input      [0:0]    port_state_in_3_3_0,
  input      [0:0]    port_state_in_3_3_1,
  input      [0:0]    port_state_in_3_3_2,
  input      [0:0]    port_state_in_3_3_3,
  input      [0:0]    port_state_in_3_3_4,
  input      [0:0]    port_state_in_3_3_5,
  input      [0:0]    port_state_in_3_3_6,
  input      [0:0]    port_state_in_3_3_7,
  input      [0:0]    port_state_in_4_0_0,
  input      [0:0]    port_state_in_4_0_1,
  input      [0:0]    port_state_in_4_0_2,
  input      [0:0]    port_state_in_4_0_3,
  input      [0:0]    port_state_in_4_0_4,
  input      [0:0]    port_state_in_4_0_5,
  input      [0:0]    port_state_in_4_0_6,
  input      [0:0]    port_state_in_4_0_7,
  input      [0:0]    port_state_in_4_1_0,
  input      [0:0]    port_state_in_4_1_1,
  input      [0:0]    port_state_in_4_1_2,
  input      [0:0]    port_state_in_4_1_3,
  input      [0:0]    port_state_in_4_1_4,
  input      [0:0]    port_state_in_4_1_5,
  input      [0:0]    port_state_in_4_1_6,
  input      [0:0]    port_state_in_4_1_7,
  input      [0:0]    port_state_in_4_2_0,
  input      [0:0]    port_state_in_4_2_1,
  input      [0:0]    port_state_in_4_2_2,
  input      [0:0]    port_state_in_4_2_3,
  input      [0:0]    port_state_in_4_2_4,
  input      [0:0]    port_state_in_4_2_5,
  input      [0:0]    port_state_in_4_2_6,
  input      [0:0]    port_state_in_4_2_7,
  input      [0:0]    port_state_in_4_3_0,
  input      [0:0]    port_state_in_4_3_1,
  input      [0:0]    port_state_in_4_3_2,
  input      [0:0]    port_state_in_4_3_3,
  input      [0:0]    port_state_in_4_3_4,
  input      [0:0]    port_state_in_4_3_5,
  input      [0:0]    port_state_in_4_3_6,
  input      [0:0]    port_state_in_4_3_7,
  input      [0:0]    port_state_in_5_0_0,
  input      [0:0]    port_state_in_5_0_1,
  input      [0:0]    port_state_in_5_0_2,
  input      [0:0]    port_state_in_5_0_3,
  input      [0:0]    port_state_in_5_0_4,
  input      [0:0]    port_state_in_5_0_5,
  input      [0:0]    port_state_in_5_0_6,
  input      [0:0]    port_state_in_5_0_7,
  input      [0:0]    port_state_in_5_1_0,
  input      [0:0]    port_state_in_5_1_1,
  input      [0:0]    port_state_in_5_1_2,
  input      [0:0]    port_state_in_5_1_3,
  input      [0:0]    port_state_in_5_1_4,
  input      [0:0]    port_state_in_5_1_5,
  input      [0:0]    port_state_in_5_1_6,
  input      [0:0]    port_state_in_5_1_7,
  input      [0:0]    port_state_in_5_2_0,
  input      [0:0]    port_state_in_5_2_1,
  input      [0:0]    port_state_in_5_2_2,
  input      [0:0]    port_state_in_5_2_3,
  input      [0:0]    port_state_in_5_2_4,
  input      [0:0]    port_state_in_5_2_5,
  input      [0:0]    port_state_in_5_2_6,
  input      [0:0]    port_state_in_5_2_7,
  input      [0:0]    port_state_in_5_3_0,
  input      [0:0]    port_state_in_5_3_1,
  input      [0:0]    port_state_in_5_3_2,
  input      [0:0]    port_state_in_5_3_3,
  input      [0:0]    port_state_in_5_3_4,
  input      [0:0]    port_state_in_5_3_5,
  input      [0:0]    port_state_in_5_3_6,
  input      [0:0]    port_state_in_5_3_7,
  input      [0:0]    port_state_in_6_0_0,
  input      [0:0]    port_state_in_6_0_1,
  input      [0:0]    port_state_in_6_0_2,
  input      [0:0]    port_state_in_6_0_3,
  input      [0:0]    port_state_in_6_0_4,
  input      [0:0]    port_state_in_6_0_5,
  input      [0:0]    port_state_in_6_0_6,
  input      [0:0]    port_state_in_6_0_7,
  input      [0:0]    port_state_in_6_1_0,
  input      [0:0]    port_state_in_6_1_1,
  input      [0:0]    port_state_in_6_1_2,
  input      [0:0]    port_state_in_6_1_3,
  input      [0:0]    port_state_in_6_1_4,
  input      [0:0]    port_state_in_6_1_5,
  input      [0:0]    port_state_in_6_1_6,
  input      [0:0]    port_state_in_6_1_7,
  input      [0:0]    port_state_in_6_2_0,
  input      [0:0]    port_state_in_6_2_1,
  input      [0:0]    port_state_in_6_2_2,
  input      [0:0]    port_state_in_6_2_3,
  input      [0:0]    port_state_in_6_2_4,
  input      [0:0]    port_state_in_6_2_5,
  input      [0:0]    port_state_in_6_2_6,
  input      [0:0]    port_state_in_6_2_7,
  input      [0:0]    port_state_in_6_3_0,
  input      [0:0]    port_state_in_6_3_1,
  input      [0:0]    port_state_in_6_3_2,
  input      [0:0]    port_state_in_6_3_3,
  input      [0:0]    port_state_in_6_3_4,
  input      [0:0]    port_state_in_6_3_5,
  input      [0:0]    port_state_in_6_3_6,
  input      [0:0]    port_state_in_6_3_7,
  input      [0:0]    port_state_in_7_0_0,
  input      [0:0]    port_state_in_7_0_1,
  input      [0:0]    port_state_in_7_0_2,
  input      [0:0]    port_state_in_7_0_3,
  input      [0:0]    port_state_in_7_0_4,
  input      [0:0]    port_state_in_7_0_5,
  input      [0:0]    port_state_in_7_0_6,
  input      [0:0]    port_state_in_7_0_7,
  input      [0:0]    port_state_in_7_1_0,
  input      [0:0]    port_state_in_7_1_1,
  input      [0:0]    port_state_in_7_1_2,
  input      [0:0]    port_state_in_7_1_3,
  input      [0:0]    port_state_in_7_1_4,
  input      [0:0]    port_state_in_7_1_5,
  input      [0:0]    port_state_in_7_1_6,
  input      [0:0]    port_state_in_7_1_7,
  input      [0:0]    port_state_in_7_2_0,
  input      [0:0]    port_state_in_7_2_1,
  input      [0:0]    port_state_in_7_2_2,
  input      [0:0]    port_state_in_7_2_3,
  input      [0:0]    port_state_in_7_2_4,
  input      [0:0]    port_state_in_7_2_5,
  input      [0:0]    port_state_in_7_2_6,
  input      [0:0]    port_state_in_7_2_7,
  input      [0:0]    port_state_in_7_3_0,
  input      [0:0]    port_state_in_7_3_1,
  input      [0:0]    port_state_in_7_3_2,
  input      [0:0]    port_state_in_7_3_3,
  input      [0:0]    port_state_in_7_3_4,
  input      [0:0]    port_state_in_7_3_5,
  input      [0:0]    port_state_in_7_3_6,
  input      [0:0]    port_state_in_7_3_7,
  input      [0:0]    port_state_in_8_0_0,
  input      [0:0]    port_state_in_8_0_1,
  input      [0:0]    port_state_in_8_0_2,
  input      [0:0]    port_state_in_8_0_3,
  input      [0:0]    port_state_in_8_0_4,
  input      [0:0]    port_state_in_8_0_5,
  input      [0:0]    port_state_in_8_0_6,
  input      [0:0]    port_state_in_8_0_7,
  input      [0:0]    port_state_in_8_1_0,
  input      [0:0]    port_state_in_8_1_1,
  input      [0:0]    port_state_in_8_1_2,
  input      [0:0]    port_state_in_8_1_3,
  input      [0:0]    port_state_in_8_1_4,
  input      [0:0]    port_state_in_8_1_5,
  input      [0:0]    port_state_in_8_1_6,
  input      [0:0]    port_state_in_8_1_7,
  input      [0:0]    port_state_in_8_2_0,
  input      [0:0]    port_state_in_8_2_1,
  input      [0:0]    port_state_in_8_2_2,
  input      [0:0]    port_state_in_8_2_3,
  input      [0:0]    port_state_in_8_2_4,
  input      [0:0]    port_state_in_8_2_5,
  input      [0:0]    port_state_in_8_2_6,
  input      [0:0]    port_state_in_8_2_7,
  input      [0:0]    port_state_in_8_3_0,
  input      [0:0]    port_state_in_8_3_1,
  input      [0:0]    port_state_in_8_3_2,
  input      [0:0]    port_state_in_8_3_3,
  input      [0:0]    port_state_in_8_3_4,
  input      [0:0]    port_state_in_8_3_5,
  input      [0:0]    port_state_in_8_3_6,
  input      [0:0]    port_state_in_8_3_7,
  input      [0:0]    port_state_in_9_0_0,
  input      [0:0]    port_state_in_9_0_1,
  input      [0:0]    port_state_in_9_0_2,
  input      [0:0]    port_state_in_9_0_3,
  input      [0:0]    port_state_in_9_0_4,
  input      [0:0]    port_state_in_9_0_5,
  input      [0:0]    port_state_in_9_0_6,
  input      [0:0]    port_state_in_9_0_7,
  input      [0:0]    port_state_in_9_1_0,
  input      [0:0]    port_state_in_9_1_1,
  input      [0:0]    port_state_in_9_1_2,
  input      [0:0]    port_state_in_9_1_3,
  input      [0:0]    port_state_in_9_1_4,
  input      [0:0]    port_state_in_9_1_5,
  input      [0:0]    port_state_in_9_1_6,
  input      [0:0]    port_state_in_9_1_7,
  input      [0:0]    port_state_in_9_2_0,
  input      [0:0]    port_state_in_9_2_1,
  input      [0:0]    port_state_in_9_2_2,
  input      [0:0]    port_state_in_9_2_3,
  input      [0:0]    port_state_in_9_2_4,
  input      [0:0]    port_state_in_9_2_5,
  input      [0:0]    port_state_in_9_2_6,
  input      [0:0]    port_state_in_9_2_7,
  input      [0:0]    port_state_in_9_3_0,
  input      [0:0]    port_state_in_9_3_1,
  input      [0:0]    port_state_in_9_3_2,
  input      [0:0]    port_state_in_9_3_3,
  input      [0:0]    port_state_in_9_3_4,
  input      [0:0]    port_state_in_9_3_5,
  input      [0:0]    port_state_in_9_3_6,
  input      [0:0]    port_state_in_9_3_7,
  input      [0:0]    port_state_in_10_0_0,
  input      [0:0]    port_state_in_10_0_1,
  input      [0:0]    port_state_in_10_0_2,
  input      [0:0]    port_state_in_10_0_3,
  input      [0:0]    port_state_in_10_0_4,
  input      [0:0]    port_state_in_10_0_5,
  input      [0:0]    port_state_in_10_0_6,
  input      [0:0]    port_state_in_10_0_7,
  input      [0:0]    port_state_in_10_1_0,
  input      [0:0]    port_state_in_10_1_1,
  input      [0:0]    port_state_in_10_1_2,
  input      [0:0]    port_state_in_10_1_3,
  input      [0:0]    port_state_in_10_1_4,
  input      [0:0]    port_state_in_10_1_5,
  input      [0:0]    port_state_in_10_1_6,
  input      [0:0]    port_state_in_10_1_7,
  input      [0:0]    port_state_in_10_2_0,
  input      [0:0]    port_state_in_10_2_1,
  input      [0:0]    port_state_in_10_2_2,
  input      [0:0]    port_state_in_10_2_3,
  input      [0:0]    port_state_in_10_2_4,
  input      [0:0]    port_state_in_10_2_5,
  input      [0:0]    port_state_in_10_2_6,
  input      [0:0]    port_state_in_10_2_7,
  input      [0:0]    port_state_in_10_3_0,
  input      [0:0]    port_state_in_10_3_1,
  input      [0:0]    port_state_in_10_3_2,
  input      [0:0]    port_state_in_10_3_3,
  input      [0:0]    port_state_in_10_3_4,
  input      [0:0]    port_state_in_10_3_5,
  input      [0:0]    port_state_in_10_3_6,
  input      [0:0]    port_state_in_10_3_7,
  input      [0:0]    port_state_in_11_0_0,
  input      [0:0]    port_state_in_11_0_1,
  input      [0:0]    port_state_in_11_0_2,
  input      [0:0]    port_state_in_11_0_3,
  input      [0:0]    port_state_in_11_0_4,
  input      [0:0]    port_state_in_11_0_5,
  input      [0:0]    port_state_in_11_0_6,
  input      [0:0]    port_state_in_11_0_7,
  input      [0:0]    port_state_in_11_1_0,
  input      [0:0]    port_state_in_11_1_1,
  input      [0:0]    port_state_in_11_1_2,
  input      [0:0]    port_state_in_11_1_3,
  input      [0:0]    port_state_in_11_1_4,
  input      [0:0]    port_state_in_11_1_5,
  input      [0:0]    port_state_in_11_1_6,
  input      [0:0]    port_state_in_11_1_7,
  input      [0:0]    port_state_in_11_2_0,
  input      [0:0]    port_state_in_11_2_1,
  input      [0:0]    port_state_in_11_2_2,
  input      [0:0]    port_state_in_11_2_3,
  input      [0:0]    port_state_in_11_2_4,
  input      [0:0]    port_state_in_11_2_5,
  input      [0:0]    port_state_in_11_2_6,
  input      [0:0]    port_state_in_11_2_7,
  input      [0:0]    port_state_in_11_3_0,
  input      [0:0]    port_state_in_11_3_1,
  input      [0:0]    port_state_in_11_3_2,
  input      [0:0]    port_state_in_11_3_3,
  input      [0:0]    port_state_in_11_3_4,
  input      [0:0]    port_state_in_11_3_5,
  input      [0:0]    port_state_in_11_3_6,
  input      [0:0]    port_state_in_11_3_7,
  input      [0:0]    port_state_in_12_0_0,
  input      [0:0]    port_state_in_12_0_1,
  input      [0:0]    port_state_in_12_0_2,
  input      [0:0]    port_state_in_12_0_3,
  input      [0:0]    port_state_in_12_0_4,
  input      [0:0]    port_state_in_12_0_5,
  input      [0:0]    port_state_in_12_0_6,
  input      [0:0]    port_state_in_12_0_7,
  input      [0:0]    port_state_in_12_1_0,
  input      [0:0]    port_state_in_12_1_1,
  input      [0:0]    port_state_in_12_1_2,
  input      [0:0]    port_state_in_12_1_3,
  input      [0:0]    port_state_in_12_1_4,
  input      [0:0]    port_state_in_12_1_5,
  input      [0:0]    port_state_in_12_1_6,
  input      [0:0]    port_state_in_12_1_7,
  input      [0:0]    port_state_in_12_2_0,
  input      [0:0]    port_state_in_12_2_1,
  input      [0:0]    port_state_in_12_2_2,
  input      [0:0]    port_state_in_12_2_3,
  input      [0:0]    port_state_in_12_2_4,
  input      [0:0]    port_state_in_12_2_5,
  input      [0:0]    port_state_in_12_2_6,
  input      [0:0]    port_state_in_12_2_7,
  input      [0:0]    port_state_in_12_3_0,
  input      [0:0]    port_state_in_12_3_1,
  input      [0:0]    port_state_in_12_3_2,
  input      [0:0]    port_state_in_12_3_3,
  input      [0:0]    port_state_in_12_3_4,
  input      [0:0]    port_state_in_12_3_5,
  input      [0:0]    port_state_in_12_3_6,
  input      [0:0]    port_state_in_12_3_7,
  input      [0:0]    port_state_in_13_0_0,
  input      [0:0]    port_state_in_13_0_1,
  input      [0:0]    port_state_in_13_0_2,
  input      [0:0]    port_state_in_13_0_3,
  input      [0:0]    port_state_in_13_0_4,
  input      [0:0]    port_state_in_13_0_5,
  input      [0:0]    port_state_in_13_0_6,
  input      [0:0]    port_state_in_13_0_7,
  input      [0:0]    port_state_in_13_1_0,
  input      [0:0]    port_state_in_13_1_1,
  input      [0:0]    port_state_in_13_1_2,
  input      [0:0]    port_state_in_13_1_3,
  input      [0:0]    port_state_in_13_1_4,
  input      [0:0]    port_state_in_13_1_5,
  input      [0:0]    port_state_in_13_1_6,
  input      [0:0]    port_state_in_13_1_7,
  input      [0:0]    port_state_in_13_2_0,
  input      [0:0]    port_state_in_13_2_1,
  input      [0:0]    port_state_in_13_2_2,
  input      [0:0]    port_state_in_13_2_3,
  input      [0:0]    port_state_in_13_2_4,
  input      [0:0]    port_state_in_13_2_5,
  input      [0:0]    port_state_in_13_2_6,
  input      [0:0]    port_state_in_13_2_7,
  input      [0:0]    port_state_in_13_3_0,
  input      [0:0]    port_state_in_13_3_1,
  input      [0:0]    port_state_in_13_3_2,
  input      [0:0]    port_state_in_13_3_3,
  input      [0:0]    port_state_in_13_3_4,
  input      [0:0]    port_state_in_13_3_5,
  input      [0:0]    port_state_in_13_3_6,
  input      [0:0]    port_state_in_13_3_7,
  input      [0:0]    port_state_in_14_0_0,
  input      [0:0]    port_state_in_14_0_1,
  input      [0:0]    port_state_in_14_0_2,
  input      [0:0]    port_state_in_14_0_3,
  input      [0:0]    port_state_in_14_0_4,
  input      [0:0]    port_state_in_14_0_5,
  input      [0:0]    port_state_in_14_0_6,
  input      [0:0]    port_state_in_14_0_7,
  input      [0:0]    port_state_in_14_1_0,
  input      [0:0]    port_state_in_14_1_1,
  input      [0:0]    port_state_in_14_1_2,
  input      [0:0]    port_state_in_14_1_3,
  input      [0:0]    port_state_in_14_1_4,
  input      [0:0]    port_state_in_14_1_5,
  input      [0:0]    port_state_in_14_1_6,
  input      [0:0]    port_state_in_14_1_7,
  input      [0:0]    port_state_in_14_2_0,
  input      [0:0]    port_state_in_14_2_1,
  input      [0:0]    port_state_in_14_2_2,
  input      [0:0]    port_state_in_14_2_3,
  input      [0:0]    port_state_in_14_2_4,
  input      [0:0]    port_state_in_14_2_5,
  input      [0:0]    port_state_in_14_2_6,
  input      [0:0]    port_state_in_14_2_7,
  input      [0:0]    port_state_in_14_3_0,
  input      [0:0]    port_state_in_14_3_1,
  input      [0:0]    port_state_in_14_3_2,
  input      [0:0]    port_state_in_14_3_3,
  input      [0:0]    port_state_in_14_3_4,
  input      [0:0]    port_state_in_14_3_5,
  input      [0:0]    port_state_in_14_3_6,
  input      [0:0]    port_state_in_14_3_7,
  input      [0:0]    port_state_in_15_0_0,
  input      [0:0]    port_state_in_15_0_1,
  input      [0:0]    port_state_in_15_0_2,
  input      [0:0]    port_state_in_15_0_3,
  input      [0:0]    port_state_in_15_0_4,
  input      [0:0]    port_state_in_15_0_5,
  input      [0:0]    port_state_in_15_0_6,
  input      [0:0]    port_state_in_15_0_7,
  input      [0:0]    port_state_in_15_1_0,
  input      [0:0]    port_state_in_15_1_1,
  input      [0:0]    port_state_in_15_1_2,
  input      [0:0]    port_state_in_15_1_3,
  input      [0:0]    port_state_in_15_1_4,
  input      [0:0]    port_state_in_15_1_5,
  input      [0:0]    port_state_in_15_1_6,
  input      [0:0]    port_state_in_15_1_7,
  input      [0:0]    port_state_in_15_2_0,
  input      [0:0]    port_state_in_15_2_1,
  input      [0:0]    port_state_in_15_2_2,
  input      [0:0]    port_state_in_15_2_3,
  input      [0:0]    port_state_in_15_2_4,
  input      [0:0]    port_state_in_15_2_5,
  input      [0:0]    port_state_in_15_2_6,
  input      [0:0]    port_state_in_15_2_7,
  input      [0:0]    port_state_in_15_3_0,
  input      [0:0]    port_state_in_15_3_1,
  input      [0:0]    port_state_in_15_3_2,
  input      [0:0]    port_state_in_15_3_3,
  input      [0:0]    port_state_in_15_3_4,
  input      [0:0]    port_state_in_15_3_5,
  input      [0:0]    port_state_in_15_3_6,
  input      [0:0]    port_state_in_15_3_7,
  output     [0:0]    port_state_out_0_0_0,
  output     [0:0]    port_state_out_0_0_1,
  output     [0:0]    port_state_out_0_0_2,
  output     [0:0]    port_state_out_0_0_3,
  output     [0:0]    port_state_out_0_0_4,
  output     [0:0]    port_state_out_0_0_5,
  output     [0:0]    port_state_out_0_0_6,
  output     [0:0]    port_state_out_0_0_7,
  output     [0:0]    port_state_out_0_1_0,
  output     [0:0]    port_state_out_0_1_1,
  output     [0:0]    port_state_out_0_1_2,
  output     [0:0]    port_state_out_0_1_3,
  output     [0:0]    port_state_out_0_1_4,
  output     [0:0]    port_state_out_0_1_5,
  output     [0:0]    port_state_out_0_1_6,
  output     [0:0]    port_state_out_0_1_7,
  output     [0:0]    port_state_out_0_2_0,
  output     [0:0]    port_state_out_0_2_1,
  output     [0:0]    port_state_out_0_2_2,
  output     [0:0]    port_state_out_0_2_3,
  output     [0:0]    port_state_out_0_2_4,
  output     [0:0]    port_state_out_0_2_5,
  output     [0:0]    port_state_out_0_2_6,
  output     [0:0]    port_state_out_0_2_7,
  output     [0:0]    port_state_out_0_3_0,
  output     [0:0]    port_state_out_0_3_1,
  output     [0:0]    port_state_out_0_3_2,
  output     [0:0]    port_state_out_0_3_3,
  output     [0:0]    port_state_out_0_3_4,
  output     [0:0]    port_state_out_0_3_5,
  output     [0:0]    port_state_out_0_3_6,
  output     [0:0]    port_state_out_0_3_7,
  output     [0:0]    port_state_out_1_0_0,
  output     [0:0]    port_state_out_1_0_1,
  output     [0:0]    port_state_out_1_0_2,
  output     [0:0]    port_state_out_1_0_3,
  output     [0:0]    port_state_out_1_0_4,
  output     [0:0]    port_state_out_1_0_5,
  output     [0:0]    port_state_out_1_0_6,
  output     [0:0]    port_state_out_1_0_7,
  output     [0:0]    port_state_out_1_1_0,
  output     [0:0]    port_state_out_1_1_1,
  output     [0:0]    port_state_out_1_1_2,
  output     [0:0]    port_state_out_1_1_3,
  output     [0:0]    port_state_out_1_1_4,
  output     [0:0]    port_state_out_1_1_5,
  output     [0:0]    port_state_out_1_1_6,
  output     [0:0]    port_state_out_1_1_7,
  output     [0:0]    port_state_out_1_2_0,
  output     [0:0]    port_state_out_1_2_1,
  output     [0:0]    port_state_out_1_2_2,
  output     [0:0]    port_state_out_1_2_3,
  output     [0:0]    port_state_out_1_2_4,
  output     [0:0]    port_state_out_1_2_5,
  output     [0:0]    port_state_out_1_2_6,
  output     [0:0]    port_state_out_1_2_7,
  output     [0:0]    port_state_out_1_3_0,
  output     [0:0]    port_state_out_1_3_1,
  output     [0:0]    port_state_out_1_3_2,
  output     [0:0]    port_state_out_1_3_3,
  output     [0:0]    port_state_out_1_3_4,
  output     [0:0]    port_state_out_1_3_5,
  output     [0:0]    port_state_out_1_3_6,
  output     [0:0]    port_state_out_1_3_7,
  output     [0:0]    port_state_out_2_0_0,
  output     [0:0]    port_state_out_2_0_1,
  output     [0:0]    port_state_out_2_0_2,
  output     [0:0]    port_state_out_2_0_3,
  output     [0:0]    port_state_out_2_0_4,
  output     [0:0]    port_state_out_2_0_5,
  output     [0:0]    port_state_out_2_0_6,
  output     [0:0]    port_state_out_2_0_7,
  output     [0:0]    port_state_out_2_1_0,
  output     [0:0]    port_state_out_2_1_1,
  output     [0:0]    port_state_out_2_1_2,
  output     [0:0]    port_state_out_2_1_3,
  output     [0:0]    port_state_out_2_1_4,
  output     [0:0]    port_state_out_2_1_5,
  output     [0:0]    port_state_out_2_1_6,
  output     [0:0]    port_state_out_2_1_7,
  output     [0:0]    port_state_out_2_2_0,
  output     [0:0]    port_state_out_2_2_1,
  output     [0:0]    port_state_out_2_2_2,
  output     [0:0]    port_state_out_2_2_3,
  output     [0:0]    port_state_out_2_2_4,
  output     [0:0]    port_state_out_2_2_5,
  output     [0:0]    port_state_out_2_2_6,
  output     [0:0]    port_state_out_2_2_7,
  output     [0:0]    port_state_out_2_3_0,
  output     [0:0]    port_state_out_2_3_1,
  output     [0:0]    port_state_out_2_3_2,
  output     [0:0]    port_state_out_2_3_3,
  output     [0:0]    port_state_out_2_3_4,
  output     [0:0]    port_state_out_2_3_5,
  output     [0:0]    port_state_out_2_3_6,
  output     [0:0]    port_state_out_2_3_7,
  output     [0:0]    port_state_out_3_0_0,
  output     [0:0]    port_state_out_3_0_1,
  output     [0:0]    port_state_out_3_0_2,
  output     [0:0]    port_state_out_3_0_3,
  output     [0:0]    port_state_out_3_0_4,
  output     [0:0]    port_state_out_3_0_5,
  output     [0:0]    port_state_out_3_0_6,
  output     [0:0]    port_state_out_3_0_7,
  output     [0:0]    port_state_out_3_1_0,
  output     [0:0]    port_state_out_3_1_1,
  output     [0:0]    port_state_out_3_1_2,
  output     [0:0]    port_state_out_3_1_3,
  output     [0:0]    port_state_out_3_1_4,
  output     [0:0]    port_state_out_3_1_5,
  output     [0:0]    port_state_out_3_1_6,
  output     [0:0]    port_state_out_3_1_7,
  output     [0:0]    port_state_out_3_2_0,
  output     [0:0]    port_state_out_3_2_1,
  output     [0:0]    port_state_out_3_2_2,
  output     [0:0]    port_state_out_3_2_3,
  output     [0:0]    port_state_out_3_2_4,
  output     [0:0]    port_state_out_3_2_5,
  output     [0:0]    port_state_out_3_2_6,
  output     [0:0]    port_state_out_3_2_7,
  output     [0:0]    port_state_out_3_3_0,
  output     [0:0]    port_state_out_3_3_1,
  output     [0:0]    port_state_out_3_3_2,
  output     [0:0]    port_state_out_3_3_3,
  output     [0:0]    port_state_out_3_3_4,
  output     [0:0]    port_state_out_3_3_5,
  output     [0:0]    port_state_out_3_3_6,
  output     [0:0]    port_state_out_3_3_7,
  output     [0:0]    port_state_out_4_0_0,
  output     [0:0]    port_state_out_4_0_1,
  output     [0:0]    port_state_out_4_0_2,
  output     [0:0]    port_state_out_4_0_3,
  output     [0:0]    port_state_out_4_0_4,
  output     [0:0]    port_state_out_4_0_5,
  output     [0:0]    port_state_out_4_0_6,
  output     [0:0]    port_state_out_4_0_7,
  output     [0:0]    port_state_out_4_1_0,
  output     [0:0]    port_state_out_4_1_1,
  output     [0:0]    port_state_out_4_1_2,
  output     [0:0]    port_state_out_4_1_3,
  output     [0:0]    port_state_out_4_1_4,
  output     [0:0]    port_state_out_4_1_5,
  output     [0:0]    port_state_out_4_1_6,
  output     [0:0]    port_state_out_4_1_7,
  output     [0:0]    port_state_out_4_2_0,
  output     [0:0]    port_state_out_4_2_1,
  output     [0:0]    port_state_out_4_2_2,
  output     [0:0]    port_state_out_4_2_3,
  output     [0:0]    port_state_out_4_2_4,
  output     [0:0]    port_state_out_4_2_5,
  output     [0:0]    port_state_out_4_2_6,
  output     [0:0]    port_state_out_4_2_7,
  output     [0:0]    port_state_out_4_3_0,
  output     [0:0]    port_state_out_4_3_1,
  output     [0:0]    port_state_out_4_3_2,
  output     [0:0]    port_state_out_4_3_3,
  output     [0:0]    port_state_out_4_3_4,
  output     [0:0]    port_state_out_4_3_5,
  output     [0:0]    port_state_out_4_3_6,
  output     [0:0]    port_state_out_4_3_7,
  output     [0:0]    port_state_out_5_0_0,
  output     [0:0]    port_state_out_5_0_1,
  output     [0:0]    port_state_out_5_0_2,
  output     [0:0]    port_state_out_5_0_3,
  output     [0:0]    port_state_out_5_0_4,
  output     [0:0]    port_state_out_5_0_5,
  output     [0:0]    port_state_out_5_0_6,
  output     [0:0]    port_state_out_5_0_7,
  output     [0:0]    port_state_out_5_1_0,
  output     [0:0]    port_state_out_5_1_1,
  output     [0:0]    port_state_out_5_1_2,
  output     [0:0]    port_state_out_5_1_3,
  output     [0:0]    port_state_out_5_1_4,
  output     [0:0]    port_state_out_5_1_5,
  output     [0:0]    port_state_out_5_1_6,
  output     [0:0]    port_state_out_5_1_7,
  output     [0:0]    port_state_out_5_2_0,
  output     [0:0]    port_state_out_5_2_1,
  output     [0:0]    port_state_out_5_2_2,
  output     [0:0]    port_state_out_5_2_3,
  output     [0:0]    port_state_out_5_2_4,
  output     [0:0]    port_state_out_5_2_5,
  output     [0:0]    port_state_out_5_2_6,
  output     [0:0]    port_state_out_5_2_7,
  output     [0:0]    port_state_out_5_3_0,
  output     [0:0]    port_state_out_5_3_1,
  output     [0:0]    port_state_out_5_3_2,
  output     [0:0]    port_state_out_5_3_3,
  output     [0:0]    port_state_out_5_3_4,
  output     [0:0]    port_state_out_5_3_5,
  output     [0:0]    port_state_out_5_3_6,
  output     [0:0]    port_state_out_5_3_7,
  output     [0:0]    port_state_out_6_0_0,
  output     [0:0]    port_state_out_6_0_1,
  output     [0:0]    port_state_out_6_0_2,
  output     [0:0]    port_state_out_6_0_3,
  output     [0:0]    port_state_out_6_0_4,
  output     [0:0]    port_state_out_6_0_5,
  output     [0:0]    port_state_out_6_0_6,
  output     [0:0]    port_state_out_6_0_7,
  output     [0:0]    port_state_out_6_1_0,
  output     [0:0]    port_state_out_6_1_1,
  output     [0:0]    port_state_out_6_1_2,
  output     [0:0]    port_state_out_6_1_3,
  output     [0:0]    port_state_out_6_1_4,
  output     [0:0]    port_state_out_6_1_5,
  output     [0:0]    port_state_out_6_1_6,
  output     [0:0]    port_state_out_6_1_7,
  output     [0:0]    port_state_out_6_2_0,
  output     [0:0]    port_state_out_6_2_1,
  output     [0:0]    port_state_out_6_2_2,
  output     [0:0]    port_state_out_6_2_3,
  output     [0:0]    port_state_out_6_2_4,
  output     [0:0]    port_state_out_6_2_5,
  output     [0:0]    port_state_out_6_2_6,
  output     [0:0]    port_state_out_6_2_7,
  output     [0:0]    port_state_out_6_3_0,
  output     [0:0]    port_state_out_6_3_1,
  output     [0:0]    port_state_out_6_3_2,
  output     [0:0]    port_state_out_6_3_3,
  output     [0:0]    port_state_out_6_3_4,
  output     [0:0]    port_state_out_6_3_5,
  output     [0:0]    port_state_out_6_3_6,
  output     [0:0]    port_state_out_6_3_7,
  output     [0:0]    port_state_out_7_0_0,
  output     [0:0]    port_state_out_7_0_1,
  output     [0:0]    port_state_out_7_0_2,
  output     [0:0]    port_state_out_7_0_3,
  output     [0:0]    port_state_out_7_0_4,
  output     [0:0]    port_state_out_7_0_5,
  output     [0:0]    port_state_out_7_0_6,
  output     [0:0]    port_state_out_7_0_7,
  output     [0:0]    port_state_out_7_1_0,
  output     [0:0]    port_state_out_7_1_1,
  output     [0:0]    port_state_out_7_1_2,
  output     [0:0]    port_state_out_7_1_3,
  output     [0:0]    port_state_out_7_1_4,
  output     [0:0]    port_state_out_7_1_5,
  output     [0:0]    port_state_out_7_1_6,
  output     [0:0]    port_state_out_7_1_7,
  output     [0:0]    port_state_out_7_2_0,
  output     [0:0]    port_state_out_7_2_1,
  output     [0:0]    port_state_out_7_2_2,
  output     [0:0]    port_state_out_7_2_3,
  output     [0:0]    port_state_out_7_2_4,
  output     [0:0]    port_state_out_7_2_5,
  output     [0:0]    port_state_out_7_2_6,
  output     [0:0]    port_state_out_7_2_7,
  output     [0:0]    port_state_out_7_3_0,
  output     [0:0]    port_state_out_7_3_1,
  output     [0:0]    port_state_out_7_3_2,
  output     [0:0]    port_state_out_7_3_3,
  output     [0:0]    port_state_out_7_3_4,
  output     [0:0]    port_state_out_7_3_5,
  output     [0:0]    port_state_out_7_3_6,
  output     [0:0]    port_state_out_7_3_7,
  output     [0:0]    port_state_out_8_0_0,
  output     [0:0]    port_state_out_8_0_1,
  output     [0:0]    port_state_out_8_0_2,
  output     [0:0]    port_state_out_8_0_3,
  output     [0:0]    port_state_out_8_0_4,
  output     [0:0]    port_state_out_8_0_5,
  output     [0:0]    port_state_out_8_0_6,
  output     [0:0]    port_state_out_8_0_7,
  output     [0:0]    port_state_out_8_1_0,
  output     [0:0]    port_state_out_8_1_1,
  output     [0:0]    port_state_out_8_1_2,
  output     [0:0]    port_state_out_8_1_3,
  output     [0:0]    port_state_out_8_1_4,
  output     [0:0]    port_state_out_8_1_5,
  output     [0:0]    port_state_out_8_1_6,
  output     [0:0]    port_state_out_8_1_7,
  output     [0:0]    port_state_out_8_2_0,
  output     [0:0]    port_state_out_8_2_1,
  output     [0:0]    port_state_out_8_2_2,
  output     [0:0]    port_state_out_8_2_3,
  output     [0:0]    port_state_out_8_2_4,
  output     [0:0]    port_state_out_8_2_5,
  output     [0:0]    port_state_out_8_2_6,
  output     [0:0]    port_state_out_8_2_7,
  output     [0:0]    port_state_out_8_3_0,
  output     [0:0]    port_state_out_8_3_1,
  output     [0:0]    port_state_out_8_3_2,
  output     [0:0]    port_state_out_8_3_3,
  output     [0:0]    port_state_out_8_3_4,
  output     [0:0]    port_state_out_8_3_5,
  output     [0:0]    port_state_out_8_3_6,
  output     [0:0]    port_state_out_8_3_7,
  output     [0:0]    port_state_out_9_0_0,
  output     [0:0]    port_state_out_9_0_1,
  output     [0:0]    port_state_out_9_0_2,
  output     [0:0]    port_state_out_9_0_3,
  output     [0:0]    port_state_out_9_0_4,
  output     [0:0]    port_state_out_9_0_5,
  output     [0:0]    port_state_out_9_0_6,
  output     [0:0]    port_state_out_9_0_7,
  output     [0:0]    port_state_out_9_1_0,
  output     [0:0]    port_state_out_9_1_1,
  output     [0:0]    port_state_out_9_1_2,
  output     [0:0]    port_state_out_9_1_3,
  output     [0:0]    port_state_out_9_1_4,
  output     [0:0]    port_state_out_9_1_5,
  output     [0:0]    port_state_out_9_1_6,
  output     [0:0]    port_state_out_9_1_7,
  output     [0:0]    port_state_out_9_2_0,
  output     [0:0]    port_state_out_9_2_1,
  output     [0:0]    port_state_out_9_2_2,
  output     [0:0]    port_state_out_9_2_3,
  output     [0:0]    port_state_out_9_2_4,
  output     [0:0]    port_state_out_9_2_5,
  output     [0:0]    port_state_out_9_2_6,
  output     [0:0]    port_state_out_9_2_7,
  output     [0:0]    port_state_out_9_3_0,
  output     [0:0]    port_state_out_9_3_1,
  output     [0:0]    port_state_out_9_3_2,
  output     [0:0]    port_state_out_9_3_3,
  output     [0:0]    port_state_out_9_3_4,
  output     [0:0]    port_state_out_9_3_5,
  output     [0:0]    port_state_out_9_3_6,
  output     [0:0]    port_state_out_9_3_7,
  output     [0:0]    port_state_out_10_0_0,
  output     [0:0]    port_state_out_10_0_1,
  output     [0:0]    port_state_out_10_0_2,
  output     [0:0]    port_state_out_10_0_3,
  output     [0:0]    port_state_out_10_0_4,
  output     [0:0]    port_state_out_10_0_5,
  output     [0:0]    port_state_out_10_0_6,
  output     [0:0]    port_state_out_10_0_7,
  output     [0:0]    port_state_out_10_1_0,
  output     [0:0]    port_state_out_10_1_1,
  output     [0:0]    port_state_out_10_1_2,
  output     [0:0]    port_state_out_10_1_3,
  output     [0:0]    port_state_out_10_1_4,
  output     [0:0]    port_state_out_10_1_5,
  output     [0:0]    port_state_out_10_1_6,
  output     [0:0]    port_state_out_10_1_7,
  output     [0:0]    port_state_out_10_2_0,
  output     [0:0]    port_state_out_10_2_1,
  output     [0:0]    port_state_out_10_2_2,
  output     [0:0]    port_state_out_10_2_3,
  output     [0:0]    port_state_out_10_2_4,
  output     [0:0]    port_state_out_10_2_5,
  output     [0:0]    port_state_out_10_2_6,
  output     [0:0]    port_state_out_10_2_7,
  output     [0:0]    port_state_out_10_3_0,
  output     [0:0]    port_state_out_10_3_1,
  output     [0:0]    port_state_out_10_3_2,
  output     [0:0]    port_state_out_10_3_3,
  output     [0:0]    port_state_out_10_3_4,
  output     [0:0]    port_state_out_10_3_5,
  output     [0:0]    port_state_out_10_3_6,
  output     [0:0]    port_state_out_10_3_7,
  output     [0:0]    port_state_out_11_0_0,
  output     [0:0]    port_state_out_11_0_1,
  output     [0:0]    port_state_out_11_0_2,
  output     [0:0]    port_state_out_11_0_3,
  output     [0:0]    port_state_out_11_0_4,
  output     [0:0]    port_state_out_11_0_5,
  output     [0:0]    port_state_out_11_0_6,
  output     [0:0]    port_state_out_11_0_7,
  output     [0:0]    port_state_out_11_1_0,
  output     [0:0]    port_state_out_11_1_1,
  output     [0:0]    port_state_out_11_1_2,
  output     [0:0]    port_state_out_11_1_3,
  output     [0:0]    port_state_out_11_1_4,
  output     [0:0]    port_state_out_11_1_5,
  output     [0:0]    port_state_out_11_1_6,
  output     [0:0]    port_state_out_11_1_7,
  output     [0:0]    port_state_out_11_2_0,
  output     [0:0]    port_state_out_11_2_1,
  output     [0:0]    port_state_out_11_2_2,
  output     [0:0]    port_state_out_11_2_3,
  output     [0:0]    port_state_out_11_2_4,
  output     [0:0]    port_state_out_11_2_5,
  output     [0:0]    port_state_out_11_2_6,
  output     [0:0]    port_state_out_11_2_7,
  output     [0:0]    port_state_out_11_3_0,
  output     [0:0]    port_state_out_11_3_1,
  output     [0:0]    port_state_out_11_3_2,
  output     [0:0]    port_state_out_11_3_3,
  output     [0:0]    port_state_out_11_3_4,
  output     [0:0]    port_state_out_11_3_5,
  output     [0:0]    port_state_out_11_3_6,
  output     [0:0]    port_state_out_11_3_7,
  output     [0:0]    port_state_out_12_0_0,
  output     [0:0]    port_state_out_12_0_1,
  output     [0:0]    port_state_out_12_0_2,
  output     [0:0]    port_state_out_12_0_3,
  output     [0:0]    port_state_out_12_0_4,
  output     [0:0]    port_state_out_12_0_5,
  output     [0:0]    port_state_out_12_0_6,
  output     [0:0]    port_state_out_12_0_7,
  output     [0:0]    port_state_out_12_1_0,
  output     [0:0]    port_state_out_12_1_1,
  output     [0:0]    port_state_out_12_1_2,
  output     [0:0]    port_state_out_12_1_3,
  output     [0:0]    port_state_out_12_1_4,
  output     [0:0]    port_state_out_12_1_5,
  output     [0:0]    port_state_out_12_1_6,
  output     [0:0]    port_state_out_12_1_7,
  output     [0:0]    port_state_out_12_2_0,
  output     [0:0]    port_state_out_12_2_1,
  output     [0:0]    port_state_out_12_2_2,
  output     [0:0]    port_state_out_12_2_3,
  output     [0:0]    port_state_out_12_2_4,
  output     [0:0]    port_state_out_12_2_5,
  output     [0:0]    port_state_out_12_2_6,
  output     [0:0]    port_state_out_12_2_7,
  output     [0:0]    port_state_out_12_3_0,
  output     [0:0]    port_state_out_12_3_1,
  output     [0:0]    port_state_out_12_3_2,
  output     [0:0]    port_state_out_12_3_3,
  output     [0:0]    port_state_out_12_3_4,
  output     [0:0]    port_state_out_12_3_5,
  output     [0:0]    port_state_out_12_3_6,
  output     [0:0]    port_state_out_12_3_7,
  output     [0:0]    port_state_out_13_0_0,
  output     [0:0]    port_state_out_13_0_1,
  output     [0:0]    port_state_out_13_0_2,
  output     [0:0]    port_state_out_13_0_3,
  output     [0:0]    port_state_out_13_0_4,
  output     [0:0]    port_state_out_13_0_5,
  output     [0:0]    port_state_out_13_0_6,
  output     [0:0]    port_state_out_13_0_7,
  output     [0:0]    port_state_out_13_1_0,
  output     [0:0]    port_state_out_13_1_1,
  output     [0:0]    port_state_out_13_1_2,
  output     [0:0]    port_state_out_13_1_3,
  output     [0:0]    port_state_out_13_1_4,
  output     [0:0]    port_state_out_13_1_5,
  output     [0:0]    port_state_out_13_1_6,
  output     [0:0]    port_state_out_13_1_7,
  output     [0:0]    port_state_out_13_2_0,
  output     [0:0]    port_state_out_13_2_1,
  output     [0:0]    port_state_out_13_2_2,
  output     [0:0]    port_state_out_13_2_3,
  output     [0:0]    port_state_out_13_2_4,
  output     [0:0]    port_state_out_13_2_5,
  output     [0:0]    port_state_out_13_2_6,
  output     [0:0]    port_state_out_13_2_7,
  output     [0:0]    port_state_out_13_3_0,
  output     [0:0]    port_state_out_13_3_1,
  output     [0:0]    port_state_out_13_3_2,
  output     [0:0]    port_state_out_13_3_3,
  output     [0:0]    port_state_out_13_3_4,
  output     [0:0]    port_state_out_13_3_5,
  output     [0:0]    port_state_out_13_3_6,
  output     [0:0]    port_state_out_13_3_7,
  output     [0:0]    port_state_out_14_0_0,
  output     [0:0]    port_state_out_14_0_1,
  output     [0:0]    port_state_out_14_0_2,
  output     [0:0]    port_state_out_14_0_3,
  output     [0:0]    port_state_out_14_0_4,
  output     [0:0]    port_state_out_14_0_5,
  output     [0:0]    port_state_out_14_0_6,
  output     [0:0]    port_state_out_14_0_7,
  output     [0:0]    port_state_out_14_1_0,
  output     [0:0]    port_state_out_14_1_1,
  output     [0:0]    port_state_out_14_1_2,
  output     [0:0]    port_state_out_14_1_3,
  output     [0:0]    port_state_out_14_1_4,
  output     [0:0]    port_state_out_14_1_5,
  output     [0:0]    port_state_out_14_1_6,
  output     [0:0]    port_state_out_14_1_7,
  output     [0:0]    port_state_out_14_2_0,
  output     [0:0]    port_state_out_14_2_1,
  output     [0:0]    port_state_out_14_2_2,
  output     [0:0]    port_state_out_14_2_3,
  output     [0:0]    port_state_out_14_2_4,
  output     [0:0]    port_state_out_14_2_5,
  output     [0:0]    port_state_out_14_2_6,
  output     [0:0]    port_state_out_14_2_7,
  output     [0:0]    port_state_out_14_3_0,
  output     [0:0]    port_state_out_14_3_1,
  output     [0:0]    port_state_out_14_3_2,
  output     [0:0]    port_state_out_14_3_3,
  output     [0:0]    port_state_out_14_3_4,
  output     [0:0]    port_state_out_14_3_5,
  output     [0:0]    port_state_out_14_3_6,
  output     [0:0]    port_state_out_14_3_7,
  output     [0:0]    port_state_out_15_0_0,
  output     [0:0]    port_state_out_15_0_1,
  output     [0:0]    port_state_out_15_0_2,
  output     [0:0]    port_state_out_15_0_3,
  output     [0:0]    port_state_out_15_0_4,
  output     [0:0]    port_state_out_15_0_5,
  output     [0:0]    port_state_out_15_0_6,
  output     [0:0]    port_state_out_15_0_7,
  output     [0:0]    port_state_out_15_1_0,
  output     [0:0]    port_state_out_15_1_1,
  output     [0:0]    port_state_out_15_1_2,
  output     [0:0]    port_state_out_15_1_3,
  output     [0:0]    port_state_out_15_1_4,
  output     [0:0]    port_state_out_15_1_5,
  output     [0:0]    port_state_out_15_1_6,
  output     [0:0]    port_state_out_15_1_7,
  output     [0:0]    port_state_out_15_2_0,
  output     [0:0]    port_state_out_15_2_1,
  output     [0:0]    port_state_out_15_2_2,
  output     [0:0]    port_state_out_15_2_3,
  output     [0:0]    port_state_out_15_2_4,
  output     [0:0]    port_state_out_15_2_5,
  output     [0:0]    port_state_out_15_2_6,
  output     [0:0]    port_state_out_15_2_7,
  output     [0:0]    port_state_out_15_3_0,
  output     [0:0]    port_state_out_15_3_1,
  output     [0:0]    port_state_out_15_3_2,
  output     [0:0]    port_state_out_15_3_3,
  output     [0:0]    port_state_out_15_3_4,
  output     [0:0]    port_state_out_15_3_5,
  output     [0:0]    port_state_out_15_3_6,
  output     [0:0]    port_state_out_15_3_7
);

  wire       [0:0]    mul2_64_port_byte_out_0;
  wire       [0:0]    mul2_64_port_byte_out_1;
  wire       [0:0]    mul2_64_port_byte_out_2;
  wire       [0:0]    mul2_64_port_byte_out_3;
  wire       [0:0]    mul2_64_port_byte_out_4;
  wire       [0:0]    mul2_64_port_byte_out_5;
  wire       [0:0]    mul2_64_port_byte_out_6;
  wire       [0:0]    mul2_64_port_byte_out_7;
  wire       [0:0]    mul3_64_port_byte_out_0;
  wire       [0:0]    mul3_64_port_byte_out_1;
  wire       [0:0]    mul3_64_port_byte_out_2;
  wire       [0:0]    mul3_64_port_byte_out_3;
  wire       [0:0]    mul3_64_port_byte_out_4;
  wire       [0:0]    mul3_64_port_byte_out_5;
  wire       [0:0]    mul3_64_port_byte_out_6;
  wire       [0:0]    mul3_64_port_byte_out_7;
  wire       [0:0]    mul2_65_port_byte_out_0;
  wire       [0:0]    mul2_65_port_byte_out_1;
  wire       [0:0]    mul2_65_port_byte_out_2;
  wire       [0:0]    mul2_65_port_byte_out_3;
  wire       [0:0]    mul2_65_port_byte_out_4;
  wire       [0:0]    mul2_65_port_byte_out_5;
  wire       [0:0]    mul2_65_port_byte_out_6;
  wire       [0:0]    mul2_65_port_byte_out_7;
  wire       [0:0]    mul3_65_port_byte_out_0;
  wire       [0:0]    mul3_65_port_byte_out_1;
  wire       [0:0]    mul3_65_port_byte_out_2;
  wire       [0:0]    mul3_65_port_byte_out_3;
  wire       [0:0]    mul3_65_port_byte_out_4;
  wire       [0:0]    mul3_65_port_byte_out_5;
  wire       [0:0]    mul3_65_port_byte_out_6;
  wire       [0:0]    mul3_65_port_byte_out_7;
  wire       [0:0]    mul2_66_port_byte_out_0;
  wire       [0:0]    mul2_66_port_byte_out_1;
  wire       [0:0]    mul2_66_port_byte_out_2;
  wire       [0:0]    mul2_66_port_byte_out_3;
  wire       [0:0]    mul2_66_port_byte_out_4;
  wire       [0:0]    mul2_66_port_byte_out_5;
  wire       [0:0]    mul2_66_port_byte_out_6;
  wire       [0:0]    mul2_66_port_byte_out_7;
  wire       [0:0]    mul3_66_port_byte_out_0;
  wire       [0:0]    mul3_66_port_byte_out_1;
  wire       [0:0]    mul3_66_port_byte_out_2;
  wire       [0:0]    mul3_66_port_byte_out_3;
  wire       [0:0]    mul3_66_port_byte_out_4;
  wire       [0:0]    mul3_66_port_byte_out_5;
  wire       [0:0]    mul3_66_port_byte_out_6;
  wire       [0:0]    mul3_66_port_byte_out_7;
  wire       [0:0]    mul2_67_port_byte_out_0;
  wire       [0:0]    mul2_67_port_byte_out_1;
  wire       [0:0]    mul2_67_port_byte_out_2;
  wire       [0:0]    mul2_67_port_byte_out_3;
  wire       [0:0]    mul2_67_port_byte_out_4;
  wire       [0:0]    mul2_67_port_byte_out_5;
  wire       [0:0]    mul2_67_port_byte_out_6;
  wire       [0:0]    mul2_67_port_byte_out_7;
  wire       [0:0]    mul3_67_port_byte_out_0;
  wire       [0:0]    mul3_67_port_byte_out_1;
  wire       [0:0]    mul3_67_port_byte_out_2;
  wire       [0:0]    mul3_67_port_byte_out_3;
  wire       [0:0]    mul3_67_port_byte_out_4;
  wire       [0:0]    mul3_67_port_byte_out_5;
  wire       [0:0]    mul3_67_port_byte_out_6;
  wire       [0:0]    mul3_67_port_byte_out_7;
  wire       [0:0]    mul2_68_port_byte_out_0;
  wire       [0:0]    mul2_68_port_byte_out_1;
  wire       [0:0]    mul2_68_port_byte_out_2;
  wire       [0:0]    mul2_68_port_byte_out_3;
  wire       [0:0]    mul2_68_port_byte_out_4;
  wire       [0:0]    mul2_68_port_byte_out_5;
  wire       [0:0]    mul2_68_port_byte_out_6;
  wire       [0:0]    mul2_68_port_byte_out_7;
  wire       [0:0]    mul3_68_port_byte_out_0;
  wire       [0:0]    mul3_68_port_byte_out_1;
  wire       [0:0]    mul3_68_port_byte_out_2;
  wire       [0:0]    mul3_68_port_byte_out_3;
  wire       [0:0]    mul3_68_port_byte_out_4;
  wire       [0:0]    mul3_68_port_byte_out_5;
  wire       [0:0]    mul3_68_port_byte_out_6;
  wire       [0:0]    mul3_68_port_byte_out_7;
  wire       [0:0]    mul2_69_port_byte_out_0;
  wire       [0:0]    mul2_69_port_byte_out_1;
  wire       [0:0]    mul2_69_port_byte_out_2;
  wire       [0:0]    mul2_69_port_byte_out_3;
  wire       [0:0]    mul2_69_port_byte_out_4;
  wire       [0:0]    mul2_69_port_byte_out_5;
  wire       [0:0]    mul2_69_port_byte_out_6;
  wire       [0:0]    mul2_69_port_byte_out_7;
  wire       [0:0]    mul3_69_port_byte_out_0;
  wire       [0:0]    mul3_69_port_byte_out_1;
  wire       [0:0]    mul3_69_port_byte_out_2;
  wire       [0:0]    mul3_69_port_byte_out_3;
  wire       [0:0]    mul3_69_port_byte_out_4;
  wire       [0:0]    mul3_69_port_byte_out_5;
  wire       [0:0]    mul3_69_port_byte_out_6;
  wire       [0:0]    mul3_69_port_byte_out_7;
  wire       [0:0]    mul2_70_port_byte_out_0;
  wire       [0:0]    mul2_70_port_byte_out_1;
  wire       [0:0]    mul2_70_port_byte_out_2;
  wire       [0:0]    mul2_70_port_byte_out_3;
  wire       [0:0]    mul2_70_port_byte_out_4;
  wire       [0:0]    mul2_70_port_byte_out_5;
  wire       [0:0]    mul2_70_port_byte_out_6;
  wire       [0:0]    mul2_70_port_byte_out_7;
  wire       [0:0]    mul3_70_port_byte_out_0;
  wire       [0:0]    mul3_70_port_byte_out_1;
  wire       [0:0]    mul3_70_port_byte_out_2;
  wire       [0:0]    mul3_70_port_byte_out_3;
  wire       [0:0]    mul3_70_port_byte_out_4;
  wire       [0:0]    mul3_70_port_byte_out_5;
  wire       [0:0]    mul3_70_port_byte_out_6;
  wire       [0:0]    mul3_70_port_byte_out_7;
  wire       [0:0]    mul2_71_port_byte_out_0;
  wire       [0:0]    mul2_71_port_byte_out_1;
  wire       [0:0]    mul2_71_port_byte_out_2;
  wire       [0:0]    mul2_71_port_byte_out_3;
  wire       [0:0]    mul2_71_port_byte_out_4;
  wire       [0:0]    mul2_71_port_byte_out_5;
  wire       [0:0]    mul2_71_port_byte_out_6;
  wire       [0:0]    mul2_71_port_byte_out_7;
  wire       [0:0]    mul3_71_port_byte_out_0;
  wire       [0:0]    mul3_71_port_byte_out_1;
  wire       [0:0]    mul3_71_port_byte_out_2;
  wire       [0:0]    mul3_71_port_byte_out_3;
  wire       [0:0]    mul3_71_port_byte_out_4;
  wire       [0:0]    mul3_71_port_byte_out_5;
  wire       [0:0]    mul3_71_port_byte_out_6;
  wire       [0:0]    mul3_71_port_byte_out_7;
  wire       [0:0]    mul2_72_port_byte_out_0;
  wire       [0:0]    mul2_72_port_byte_out_1;
  wire       [0:0]    mul2_72_port_byte_out_2;
  wire       [0:0]    mul2_72_port_byte_out_3;
  wire       [0:0]    mul2_72_port_byte_out_4;
  wire       [0:0]    mul2_72_port_byte_out_5;
  wire       [0:0]    mul2_72_port_byte_out_6;
  wire       [0:0]    mul2_72_port_byte_out_7;
  wire       [0:0]    mul3_72_port_byte_out_0;
  wire       [0:0]    mul3_72_port_byte_out_1;
  wire       [0:0]    mul3_72_port_byte_out_2;
  wire       [0:0]    mul3_72_port_byte_out_3;
  wire       [0:0]    mul3_72_port_byte_out_4;
  wire       [0:0]    mul3_72_port_byte_out_5;
  wire       [0:0]    mul3_72_port_byte_out_6;
  wire       [0:0]    mul3_72_port_byte_out_7;
  wire       [0:0]    mul2_73_port_byte_out_0;
  wire       [0:0]    mul2_73_port_byte_out_1;
  wire       [0:0]    mul2_73_port_byte_out_2;
  wire       [0:0]    mul2_73_port_byte_out_3;
  wire       [0:0]    mul2_73_port_byte_out_4;
  wire       [0:0]    mul2_73_port_byte_out_5;
  wire       [0:0]    mul2_73_port_byte_out_6;
  wire       [0:0]    mul2_73_port_byte_out_7;
  wire       [0:0]    mul3_73_port_byte_out_0;
  wire       [0:0]    mul3_73_port_byte_out_1;
  wire       [0:0]    mul3_73_port_byte_out_2;
  wire       [0:0]    mul3_73_port_byte_out_3;
  wire       [0:0]    mul3_73_port_byte_out_4;
  wire       [0:0]    mul3_73_port_byte_out_5;
  wire       [0:0]    mul3_73_port_byte_out_6;
  wire       [0:0]    mul3_73_port_byte_out_7;
  wire       [0:0]    mul2_74_port_byte_out_0;
  wire       [0:0]    mul2_74_port_byte_out_1;
  wire       [0:0]    mul2_74_port_byte_out_2;
  wire       [0:0]    mul2_74_port_byte_out_3;
  wire       [0:0]    mul2_74_port_byte_out_4;
  wire       [0:0]    mul2_74_port_byte_out_5;
  wire       [0:0]    mul2_74_port_byte_out_6;
  wire       [0:0]    mul2_74_port_byte_out_7;
  wire       [0:0]    mul3_74_port_byte_out_0;
  wire       [0:0]    mul3_74_port_byte_out_1;
  wire       [0:0]    mul3_74_port_byte_out_2;
  wire       [0:0]    mul3_74_port_byte_out_3;
  wire       [0:0]    mul3_74_port_byte_out_4;
  wire       [0:0]    mul3_74_port_byte_out_5;
  wire       [0:0]    mul3_74_port_byte_out_6;
  wire       [0:0]    mul3_74_port_byte_out_7;
  wire       [0:0]    mul2_75_port_byte_out_0;
  wire       [0:0]    mul2_75_port_byte_out_1;
  wire       [0:0]    mul2_75_port_byte_out_2;
  wire       [0:0]    mul2_75_port_byte_out_3;
  wire       [0:0]    mul2_75_port_byte_out_4;
  wire       [0:0]    mul2_75_port_byte_out_5;
  wire       [0:0]    mul2_75_port_byte_out_6;
  wire       [0:0]    mul2_75_port_byte_out_7;
  wire       [0:0]    mul3_75_port_byte_out_0;
  wire       [0:0]    mul3_75_port_byte_out_1;
  wire       [0:0]    mul3_75_port_byte_out_2;
  wire       [0:0]    mul3_75_port_byte_out_3;
  wire       [0:0]    mul3_75_port_byte_out_4;
  wire       [0:0]    mul3_75_port_byte_out_5;
  wire       [0:0]    mul3_75_port_byte_out_6;
  wire       [0:0]    mul3_75_port_byte_out_7;
  wire       [0:0]    mul2_76_port_byte_out_0;
  wire       [0:0]    mul2_76_port_byte_out_1;
  wire       [0:0]    mul2_76_port_byte_out_2;
  wire       [0:0]    mul2_76_port_byte_out_3;
  wire       [0:0]    mul2_76_port_byte_out_4;
  wire       [0:0]    mul2_76_port_byte_out_5;
  wire       [0:0]    mul2_76_port_byte_out_6;
  wire       [0:0]    mul2_76_port_byte_out_7;
  wire       [0:0]    mul3_76_port_byte_out_0;
  wire       [0:0]    mul3_76_port_byte_out_1;
  wire       [0:0]    mul3_76_port_byte_out_2;
  wire       [0:0]    mul3_76_port_byte_out_3;
  wire       [0:0]    mul3_76_port_byte_out_4;
  wire       [0:0]    mul3_76_port_byte_out_5;
  wire       [0:0]    mul3_76_port_byte_out_6;
  wire       [0:0]    mul3_76_port_byte_out_7;
  wire       [0:0]    mul2_77_port_byte_out_0;
  wire       [0:0]    mul2_77_port_byte_out_1;
  wire       [0:0]    mul2_77_port_byte_out_2;
  wire       [0:0]    mul2_77_port_byte_out_3;
  wire       [0:0]    mul2_77_port_byte_out_4;
  wire       [0:0]    mul2_77_port_byte_out_5;
  wire       [0:0]    mul2_77_port_byte_out_6;
  wire       [0:0]    mul2_77_port_byte_out_7;
  wire       [0:0]    mul3_77_port_byte_out_0;
  wire       [0:0]    mul3_77_port_byte_out_1;
  wire       [0:0]    mul3_77_port_byte_out_2;
  wire       [0:0]    mul3_77_port_byte_out_3;
  wire       [0:0]    mul3_77_port_byte_out_4;
  wire       [0:0]    mul3_77_port_byte_out_5;
  wire       [0:0]    mul3_77_port_byte_out_6;
  wire       [0:0]    mul3_77_port_byte_out_7;
  wire       [0:0]    mul2_78_port_byte_out_0;
  wire       [0:0]    mul2_78_port_byte_out_1;
  wire       [0:0]    mul2_78_port_byte_out_2;
  wire       [0:0]    mul2_78_port_byte_out_3;
  wire       [0:0]    mul2_78_port_byte_out_4;
  wire       [0:0]    mul2_78_port_byte_out_5;
  wire       [0:0]    mul2_78_port_byte_out_6;
  wire       [0:0]    mul2_78_port_byte_out_7;
  wire       [0:0]    mul3_78_port_byte_out_0;
  wire       [0:0]    mul3_78_port_byte_out_1;
  wire       [0:0]    mul3_78_port_byte_out_2;
  wire       [0:0]    mul3_78_port_byte_out_3;
  wire       [0:0]    mul3_78_port_byte_out_4;
  wire       [0:0]    mul3_78_port_byte_out_5;
  wire       [0:0]    mul3_78_port_byte_out_6;
  wire       [0:0]    mul3_78_port_byte_out_7;
  wire       [0:0]    mul2_79_port_byte_out_0;
  wire       [0:0]    mul2_79_port_byte_out_1;
  wire       [0:0]    mul2_79_port_byte_out_2;
  wire       [0:0]    mul2_79_port_byte_out_3;
  wire       [0:0]    mul2_79_port_byte_out_4;
  wire       [0:0]    mul2_79_port_byte_out_5;
  wire       [0:0]    mul2_79_port_byte_out_6;
  wire       [0:0]    mul2_79_port_byte_out_7;
  wire       [0:0]    mul3_79_port_byte_out_0;
  wire       [0:0]    mul3_79_port_byte_out_1;
  wire       [0:0]    mul3_79_port_byte_out_2;
  wire       [0:0]    mul3_79_port_byte_out_3;
  wire       [0:0]    mul3_79_port_byte_out_4;
  wire       [0:0]    mul3_79_port_byte_out_5;
  wire       [0:0]    mul3_79_port_byte_out_6;
  wire       [0:0]    mul3_79_port_byte_out_7;
  wire       [0:0]    mul2_80_port_byte_out_0;
  wire       [0:0]    mul2_80_port_byte_out_1;
  wire       [0:0]    mul2_80_port_byte_out_2;
  wire       [0:0]    mul2_80_port_byte_out_3;
  wire       [0:0]    mul2_80_port_byte_out_4;
  wire       [0:0]    mul2_80_port_byte_out_5;
  wire       [0:0]    mul2_80_port_byte_out_6;
  wire       [0:0]    mul2_80_port_byte_out_7;
  wire       [0:0]    mul3_80_port_byte_out_0;
  wire       [0:0]    mul3_80_port_byte_out_1;
  wire       [0:0]    mul3_80_port_byte_out_2;
  wire       [0:0]    mul3_80_port_byte_out_3;
  wire       [0:0]    mul3_80_port_byte_out_4;
  wire       [0:0]    mul3_80_port_byte_out_5;
  wire       [0:0]    mul3_80_port_byte_out_6;
  wire       [0:0]    mul3_80_port_byte_out_7;
  wire       [0:0]    mul2_81_port_byte_out_0;
  wire       [0:0]    mul2_81_port_byte_out_1;
  wire       [0:0]    mul2_81_port_byte_out_2;
  wire       [0:0]    mul2_81_port_byte_out_3;
  wire       [0:0]    mul2_81_port_byte_out_4;
  wire       [0:0]    mul2_81_port_byte_out_5;
  wire       [0:0]    mul2_81_port_byte_out_6;
  wire       [0:0]    mul2_81_port_byte_out_7;
  wire       [0:0]    mul3_81_port_byte_out_0;
  wire       [0:0]    mul3_81_port_byte_out_1;
  wire       [0:0]    mul3_81_port_byte_out_2;
  wire       [0:0]    mul3_81_port_byte_out_3;
  wire       [0:0]    mul3_81_port_byte_out_4;
  wire       [0:0]    mul3_81_port_byte_out_5;
  wire       [0:0]    mul3_81_port_byte_out_6;
  wire       [0:0]    mul3_81_port_byte_out_7;
  wire       [0:0]    mul2_82_port_byte_out_0;
  wire       [0:0]    mul2_82_port_byte_out_1;
  wire       [0:0]    mul2_82_port_byte_out_2;
  wire       [0:0]    mul2_82_port_byte_out_3;
  wire       [0:0]    mul2_82_port_byte_out_4;
  wire       [0:0]    mul2_82_port_byte_out_5;
  wire       [0:0]    mul2_82_port_byte_out_6;
  wire       [0:0]    mul2_82_port_byte_out_7;
  wire       [0:0]    mul3_82_port_byte_out_0;
  wire       [0:0]    mul3_82_port_byte_out_1;
  wire       [0:0]    mul3_82_port_byte_out_2;
  wire       [0:0]    mul3_82_port_byte_out_3;
  wire       [0:0]    mul3_82_port_byte_out_4;
  wire       [0:0]    mul3_82_port_byte_out_5;
  wire       [0:0]    mul3_82_port_byte_out_6;
  wire       [0:0]    mul3_82_port_byte_out_7;
  wire       [0:0]    mul2_83_port_byte_out_0;
  wire       [0:0]    mul2_83_port_byte_out_1;
  wire       [0:0]    mul2_83_port_byte_out_2;
  wire       [0:0]    mul2_83_port_byte_out_3;
  wire       [0:0]    mul2_83_port_byte_out_4;
  wire       [0:0]    mul2_83_port_byte_out_5;
  wire       [0:0]    mul2_83_port_byte_out_6;
  wire       [0:0]    mul2_83_port_byte_out_7;
  wire       [0:0]    mul3_83_port_byte_out_0;
  wire       [0:0]    mul3_83_port_byte_out_1;
  wire       [0:0]    mul3_83_port_byte_out_2;
  wire       [0:0]    mul3_83_port_byte_out_3;
  wire       [0:0]    mul3_83_port_byte_out_4;
  wire       [0:0]    mul3_83_port_byte_out_5;
  wire       [0:0]    mul3_83_port_byte_out_6;
  wire       [0:0]    mul3_83_port_byte_out_7;
  wire       [0:0]    mul2_84_port_byte_out_0;
  wire       [0:0]    mul2_84_port_byte_out_1;
  wire       [0:0]    mul2_84_port_byte_out_2;
  wire       [0:0]    mul2_84_port_byte_out_3;
  wire       [0:0]    mul2_84_port_byte_out_4;
  wire       [0:0]    mul2_84_port_byte_out_5;
  wire       [0:0]    mul2_84_port_byte_out_6;
  wire       [0:0]    mul2_84_port_byte_out_7;
  wire       [0:0]    mul3_84_port_byte_out_0;
  wire       [0:0]    mul3_84_port_byte_out_1;
  wire       [0:0]    mul3_84_port_byte_out_2;
  wire       [0:0]    mul3_84_port_byte_out_3;
  wire       [0:0]    mul3_84_port_byte_out_4;
  wire       [0:0]    mul3_84_port_byte_out_5;
  wire       [0:0]    mul3_84_port_byte_out_6;
  wire       [0:0]    mul3_84_port_byte_out_7;
  wire       [0:0]    mul2_85_port_byte_out_0;
  wire       [0:0]    mul2_85_port_byte_out_1;
  wire       [0:0]    mul2_85_port_byte_out_2;
  wire       [0:0]    mul2_85_port_byte_out_3;
  wire       [0:0]    mul2_85_port_byte_out_4;
  wire       [0:0]    mul2_85_port_byte_out_5;
  wire       [0:0]    mul2_85_port_byte_out_6;
  wire       [0:0]    mul2_85_port_byte_out_7;
  wire       [0:0]    mul3_85_port_byte_out_0;
  wire       [0:0]    mul3_85_port_byte_out_1;
  wire       [0:0]    mul3_85_port_byte_out_2;
  wire       [0:0]    mul3_85_port_byte_out_3;
  wire       [0:0]    mul3_85_port_byte_out_4;
  wire       [0:0]    mul3_85_port_byte_out_5;
  wire       [0:0]    mul3_85_port_byte_out_6;
  wire       [0:0]    mul3_85_port_byte_out_7;
  wire       [0:0]    mul2_86_port_byte_out_0;
  wire       [0:0]    mul2_86_port_byte_out_1;
  wire       [0:0]    mul2_86_port_byte_out_2;
  wire       [0:0]    mul2_86_port_byte_out_3;
  wire       [0:0]    mul2_86_port_byte_out_4;
  wire       [0:0]    mul2_86_port_byte_out_5;
  wire       [0:0]    mul2_86_port_byte_out_6;
  wire       [0:0]    mul2_86_port_byte_out_7;
  wire       [0:0]    mul3_86_port_byte_out_0;
  wire       [0:0]    mul3_86_port_byte_out_1;
  wire       [0:0]    mul3_86_port_byte_out_2;
  wire       [0:0]    mul3_86_port_byte_out_3;
  wire       [0:0]    mul3_86_port_byte_out_4;
  wire       [0:0]    mul3_86_port_byte_out_5;
  wire       [0:0]    mul3_86_port_byte_out_6;
  wire       [0:0]    mul3_86_port_byte_out_7;
  wire       [0:0]    mul2_87_port_byte_out_0;
  wire       [0:0]    mul2_87_port_byte_out_1;
  wire       [0:0]    mul2_87_port_byte_out_2;
  wire       [0:0]    mul2_87_port_byte_out_3;
  wire       [0:0]    mul2_87_port_byte_out_4;
  wire       [0:0]    mul2_87_port_byte_out_5;
  wire       [0:0]    mul2_87_port_byte_out_6;
  wire       [0:0]    mul2_87_port_byte_out_7;
  wire       [0:0]    mul3_87_port_byte_out_0;
  wire       [0:0]    mul3_87_port_byte_out_1;
  wire       [0:0]    mul3_87_port_byte_out_2;
  wire       [0:0]    mul3_87_port_byte_out_3;
  wire       [0:0]    mul3_87_port_byte_out_4;
  wire       [0:0]    mul3_87_port_byte_out_5;
  wire       [0:0]    mul3_87_port_byte_out_6;
  wire       [0:0]    mul3_87_port_byte_out_7;
  wire       [0:0]    mul2_88_port_byte_out_0;
  wire       [0:0]    mul2_88_port_byte_out_1;
  wire       [0:0]    mul2_88_port_byte_out_2;
  wire       [0:0]    mul2_88_port_byte_out_3;
  wire       [0:0]    mul2_88_port_byte_out_4;
  wire       [0:0]    mul2_88_port_byte_out_5;
  wire       [0:0]    mul2_88_port_byte_out_6;
  wire       [0:0]    mul2_88_port_byte_out_7;
  wire       [0:0]    mul3_88_port_byte_out_0;
  wire       [0:0]    mul3_88_port_byte_out_1;
  wire       [0:0]    mul3_88_port_byte_out_2;
  wire       [0:0]    mul3_88_port_byte_out_3;
  wire       [0:0]    mul3_88_port_byte_out_4;
  wire       [0:0]    mul3_88_port_byte_out_5;
  wire       [0:0]    mul3_88_port_byte_out_6;
  wire       [0:0]    mul3_88_port_byte_out_7;
  wire       [0:0]    mul2_89_port_byte_out_0;
  wire       [0:0]    mul2_89_port_byte_out_1;
  wire       [0:0]    mul2_89_port_byte_out_2;
  wire       [0:0]    mul2_89_port_byte_out_3;
  wire       [0:0]    mul2_89_port_byte_out_4;
  wire       [0:0]    mul2_89_port_byte_out_5;
  wire       [0:0]    mul2_89_port_byte_out_6;
  wire       [0:0]    mul2_89_port_byte_out_7;
  wire       [0:0]    mul3_89_port_byte_out_0;
  wire       [0:0]    mul3_89_port_byte_out_1;
  wire       [0:0]    mul3_89_port_byte_out_2;
  wire       [0:0]    mul3_89_port_byte_out_3;
  wire       [0:0]    mul3_89_port_byte_out_4;
  wire       [0:0]    mul3_89_port_byte_out_5;
  wire       [0:0]    mul3_89_port_byte_out_6;
  wire       [0:0]    mul3_89_port_byte_out_7;
  wire       [0:0]    mul2_90_port_byte_out_0;
  wire       [0:0]    mul2_90_port_byte_out_1;
  wire       [0:0]    mul2_90_port_byte_out_2;
  wire       [0:0]    mul2_90_port_byte_out_3;
  wire       [0:0]    mul2_90_port_byte_out_4;
  wire       [0:0]    mul2_90_port_byte_out_5;
  wire       [0:0]    mul2_90_port_byte_out_6;
  wire       [0:0]    mul2_90_port_byte_out_7;
  wire       [0:0]    mul3_90_port_byte_out_0;
  wire       [0:0]    mul3_90_port_byte_out_1;
  wire       [0:0]    mul3_90_port_byte_out_2;
  wire       [0:0]    mul3_90_port_byte_out_3;
  wire       [0:0]    mul3_90_port_byte_out_4;
  wire       [0:0]    mul3_90_port_byte_out_5;
  wire       [0:0]    mul3_90_port_byte_out_6;
  wire       [0:0]    mul3_90_port_byte_out_7;
  wire       [0:0]    mul2_91_port_byte_out_0;
  wire       [0:0]    mul2_91_port_byte_out_1;
  wire       [0:0]    mul2_91_port_byte_out_2;
  wire       [0:0]    mul2_91_port_byte_out_3;
  wire       [0:0]    mul2_91_port_byte_out_4;
  wire       [0:0]    mul2_91_port_byte_out_5;
  wire       [0:0]    mul2_91_port_byte_out_6;
  wire       [0:0]    mul2_91_port_byte_out_7;
  wire       [0:0]    mul3_91_port_byte_out_0;
  wire       [0:0]    mul3_91_port_byte_out_1;
  wire       [0:0]    mul3_91_port_byte_out_2;
  wire       [0:0]    mul3_91_port_byte_out_3;
  wire       [0:0]    mul3_91_port_byte_out_4;
  wire       [0:0]    mul3_91_port_byte_out_5;
  wire       [0:0]    mul3_91_port_byte_out_6;
  wire       [0:0]    mul3_91_port_byte_out_7;
  wire       [0:0]    mul2_92_port_byte_out_0;
  wire       [0:0]    mul2_92_port_byte_out_1;
  wire       [0:0]    mul2_92_port_byte_out_2;
  wire       [0:0]    mul2_92_port_byte_out_3;
  wire       [0:0]    mul2_92_port_byte_out_4;
  wire       [0:0]    mul2_92_port_byte_out_5;
  wire       [0:0]    mul2_92_port_byte_out_6;
  wire       [0:0]    mul2_92_port_byte_out_7;
  wire       [0:0]    mul3_92_port_byte_out_0;
  wire       [0:0]    mul3_92_port_byte_out_1;
  wire       [0:0]    mul3_92_port_byte_out_2;
  wire       [0:0]    mul3_92_port_byte_out_3;
  wire       [0:0]    mul3_92_port_byte_out_4;
  wire       [0:0]    mul3_92_port_byte_out_5;
  wire       [0:0]    mul3_92_port_byte_out_6;
  wire       [0:0]    mul3_92_port_byte_out_7;
  wire       [0:0]    mul2_93_port_byte_out_0;
  wire       [0:0]    mul2_93_port_byte_out_1;
  wire       [0:0]    mul2_93_port_byte_out_2;
  wire       [0:0]    mul2_93_port_byte_out_3;
  wire       [0:0]    mul2_93_port_byte_out_4;
  wire       [0:0]    mul2_93_port_byte_out_5;
  wire       [0:0]    mul2_93_port_byte_out_6;
  wire       [0:0]    mul2_93_port_byte_out_7;
  wire       [0:0]    mul3_93_port_byte_out_0;
  wire       [0:0]    mul3_93_port_byte_out_1;
  wire       [0:0]    mul3_93_port_byte_out_2;
  wire       [0:0]    mul3_93_port_byte_out_3;
  wire       [0:0]    mul3_93_port_byte_out_4;
  wire       [0:0]    mul3_93_port_byte_out_5;
  wire       [0:0]    mul3_93_port_byte_out_6;
  wire       [0:0]    mul3_93_port_byte_out_7;
  wire       [0:0]    mul2_94_port_byte_out_0;
  wire       [0:0]    mul2_94_port_byte_out_1;
  wire       [0:0]    mul2_94_port_byte_out_2;
  wire       [0:0]    mul2_94_port_byte_out_3;
  wire       [0:0]    mul2_94_port_byte_out_4;
  wire       [0:0]    mul2_94_port_byte_out_5;
  wire       [0:0]    mul2_94_port_byte_out_6;
  wire       [0:0]    mul2_94_port_byte_out_7;
  wire       [0:0]    mul3_94_port_byte_out_0;
  wire       [0:0]    mul3_94_port_byte_out_1;
  wire       [0:0]    mul3_94_port_byte_out_2;
  wire       [0:0]    mul3_94_port_byte_out_3;
  wire       [0:0]    mul3_94_port_byte_out_4;
  wire       [0:0]    mul3_94_port_byte_out_5;
  wire       [0:0]    mul3_94_port_byte_out_6;
  wire       [0:0]    mul3_94_port_byte_out_7;
  wire       [0:0]    mul2_95_port_byte_out_0;
  wire       [0:0]    mul2_95_port_byte_out_1;
  wire       [0:0]    mul2_95_port_byte_out_2;
  wire       [0:0]    mul2_95_port_byte_out_3;
  wire       [0:0]    mul2_95_port_byte_out_4;
  wire       [0:0]    mul2_95_port_byte_out_5;
  wire       [0:0]    mul2_95_port_byte_out_6;
  wire       [0:0]    mul2_95_port_byte_out_7;
  wire       [0:0]    mul3_95_port_byte_out_0;
  wire       [0:0]    mul3_95_port_byte_out_1;
  wire       [0:0]    mul3_95_port_byte_out_2;
  wire       [0:0]    mul3_95_port_byte_out_3;
  wire       [0:0]    mul3_95_port_byte_out_4;
  wire       [0:0]    mul3_95_port_byte_out_5;
  wire       [0:0]    mul3_95_port_byte_out_6;
  wire       [0:0]    mul3_95_port_byte_out_7;
  wire       [0:0]    mul2_96_port_byte_out_0;
  wire       [0:0]    mul2_96_port_byte_out_1;
  wire       [0:0]    mul2_96_port_byte_out_2;
  wire       [0:0]    mul2_96_port_byte_out_3;
  wire       [0:0]    mul2_96_port_byte_out_4;
  wire       [0:0]    mul2_96_port_byte_out_5;
  wire       [0:0]    mul2_96_port_byte_out_6;
  wire       [0:0]    mul2_96_port_byte_out_7;
  wire       [0:0]    mul3_96_port_byte_out_0;
  wire       [0:0]    mul3_96_port_byte_out_1;
  wire       [0:0]    mul3_96_port_byte_out_2;
  wire       [0:0]    mul3_96_port_byte_out_3;
  wire       [0:0]    mul3_96_port_byte_out_4;
  wire       [0:0]    mul3_96_port_byte_out_5;
  wire       [0:0]    mul3_96_port_byte_out_6;
  wire       [0:0]    mul3_96_port_byte_out_7;
  wire       [0:0]    mul2_97_port_byte_out_0;
  wire       [0:0]    mul2_97_port_byte_out_1;
  wire       [0:0]    mul2_97_port_byte_out_2;
  wire       [0:0]    mul2_97_port_byte_out_3;
  wire       [0:0]    mul2_97_port_byte_out_4;
  wire       [0:0]    mul2_97_port_byte_out_5;
  wire       [0:0]    mul2_97_port_byte_out_6;
  wire       [0:0]    mul2_97_port_byte_out_7;
  wire       [0:0]    mul3_97_port_byte_out_0;
  wire       [0:0]    mul3_97_port_byte_out_1;
  wire       [0:0]    mul3_97_port_byte_out_2;
  wire       [0:0]    mul3_97_port_byte_out_3;
  wire       [0:0]    mul3_97_port_byte_out_4;
  wire       [0:0]    mul3_97_port_byte_out_5;
  wire       [0:0]    mul3_97_port_byte_out_6;
  wire       [0:0]    mul3_97_port_byte_out_7;
  wire       [0:0]    mul2_98_port_byte_out_0;
  wire       [0:0]    mul2_98_port_byte_out_1;
  wire       [0:0]    mul2_98_port_byte_out_2;
  wire       [0:0]    mul2_98_port_byte_out_3;
  wire       [0:0]    mul2_98_port_byte_out_4;
  wire       [0:0]    mul2_98_port_byte_out_5;
  wire       [0:0]    mul2_98_port_byte_out_6;
  wire       [0:0]    mul2_98_port_byte_out_7;
  wire       [0:0]    mul3_98_port_byte_out_0;
  wire       [0:0]    mul3_98_port_byte_out_1;
  wire       [0:0]    mul3_98_port_byte_out_2;
  wire       [0:0]    mul3_98_port_byte_out_3;
  wire       [0:0]    mul3_98_port_byte_out_4;
  wire       [0:0]    mul3_98_port_byte_out_5;
  wire       [0:0]    mul3_98_port_byte_out_6;
  wire       [0:0]    mul3_98_port_byte_out_7;
  wire       [0:0]    mul2_99_port_byte_out_0;
  wire       [0:0]    mul2_99_port_byte_out_1;
  wire       [0:0]    mul2_99_port_byte_out_2;
  wire       [0:0]    mul2_99_port_byte_out_3;
  wire       [0:0]    mul2_99_port_byte_out_4;
  wire       [0:0]    mul2_99_port_byte_out_5;
  wire       [0:0]    mul2_99_port_byte_out_6;
  wire       [0:0]    mul2_99_port_byte_out_7;
  wire       [0:0]    mul3_99_port_byte_out_0;
  wire       [0:0]    mul3_99_port_byte_out_1;
  wire       [0:0]    mul3_99_port_byte_out_2;
  wire       [0:0]    mul3_99_port_byte_out_3;
  wire       [0:0]    mul3_99_port_byte_out_4;
  wire       [0:0]    mul3_99_port_byte_out_5;
  wire       [0:0]    mul3_99_port_byte_out_6;
  wire       [0:0]    mul3_99_port_byte_out_7;
  wire       [0:0]    mul2_100_port_byte_out_0;
  wire       [0:0]    mul2_100_port_byte_out_1;
  wire       [0:0]    mul2_100_port_byte_out_2;
  wire       [0:0]    mul2_100_port_byte_out_3;
  wire       [0:0]    mul2_100_port_byte_out_4;
  wire       [0:0]    mul2_100_port_byte_out_5;
  wire       [0:0]    mul2_100_port_byte_out_6;
  wire       [0:0]    mul2_100_port_byte_out_7;
  wire       [0:0]    mul3_100_port_byte_out_0;
  wire       [0:0]    mul3_100_port_byte_out_1;
  wire       [0:0]    mul3_100_port_byte_out_2;
  wire       [0:0]    mul3_100_port_byte_out_3;
  wire       [0:0]    mul3_100_port_byte_out_4;
  wire       [0:0]    mul3_100_port_byte_out_5;
  wire       [0:0]    mul3_100_port_byte_out_6;
  wire       [0:0]    mul3_100_port_byte_out_7;
  wire       [0:0]    mul2_101_port_byte_out_0;
  wire       [0:0]    mul2_101_port_byte_out_1;
  wire       [0:0]    mul2_101_port_byte_out_2;
  wire       [0:0]    mul2_101_port_byte_out_3;
  wire       [0:0]    mul2_101_port_byte_out_4;
  wire       [0:0]    mul2_101_port_byte_out_5;
  wire       [0:0]    mul2_101_port_byte_out_6;
  wire       [0:0]    mul2_101_port_byte_out_7;
  wire       [0:0]    mul3_101_port_byte_out_0;
  wire       [0:0]    mul3_101_port_byte_out_1;
  wire       [0:0]    mul3_101_port_byte_out_2;
  wire       [0:0]    mul3_101_port_byte_out_3;
  wire       [0:0]    mul3_101_port_byte_out_4;
  wire       [0:0]    mul3_101_port_byte_out_5;
  wire       [0:0]    mul3_101_port_byte_out_6;
  wire       [0:0]    mul3_101_port_byte_out_7;
  wire       [0:0]    mul2_102_port_byte_out_0;
  wire       [0:0]    mul2_102_port_byte_out_1;
  wire       [0:0]    mul2_102_port_byte_out_2;
  wire       [0:0]    mul2_102_port_byte_out_3;
  wire       [0:0]    mul2_102_port_byte_out_4;
  wire       [0:0]    mul2_102_port_byte_out_5;
  wire       [0:0]    mul2_102_port_byte_out_6;
  wire       [0:0]    mul2_102_port_byte_out_7;
  wire       [0:0]    mul3_102_port_byte_out_0;
  wire       [0:0]    mul3_102_port_byte_out_1;
  wire       [0:0]    mul3_102_port_byte_out_2;
  wire       [0:0]    mul3_102_port_byte_out_3;
  wire       [0:0]    mul3_102_port_byte_out_4;
  wire       [0:0]    mul3_102_port_byte_out_5;
  wire       [0:0]    mul3_102_port_byte_out_6;
  wire       [0:0]    mul3_102_port_byte_out_7;
  wire       [0:0]    mul2_103_port_byte_out_0;
  wire       [0:0]    mul2_103_port_byte_out_1;
  wire       [0:0]    mul2_103_port_byte_out_2;
  wire       [0:0]    mul2_103_port_byte_out_3;
  wire       [0:0]    mul2_103_port_byte_out_4;
  wire       [0:0]    mul2_103_port_byte_out_5;
  wire       [0:0]    mul2_103_port_byte_out_6;
  wire       [0:0]    mul2_103_port_byte_out_7;
  wire       [0:0]    mul3_103_port_byte_out_0;
  wire       [0:0]    mul3_103_port_byte_out_1;
  wire       [0:0]    mul3_103_port_byte_out_2;
  wire       [0:0]    mul3_103_port_byte_out_3;
  wire       [0:0]    mul3_103_port_byte_out_4;
  wire       [0:0]    mul3_103_port_byte_out_5;
  wire       [0:0]    mul3_103_port_byte_out_6;
  wire       [0:0]    mul3_103_port_byte_out_7;
  wire       [0:0]    mul2_104_port_byte_out_0;
  wire       [0:0]    mul2_104_port_byte_out_1;
  wire       [0:0]    mul2_104_port_byte_out_2;
  wire       [0:0]    mul2_104_port_byte_out_3;
  wire       [0:0]    mul2_104_port_byte_out_4;
  wire       [0:0]    mul2_104_port_byte_out_5;
  wire       [0:0]    mul2_104_port_byte_out_6;
  wire       [0:0]    mul2_104_port_byte_out_7;
  wire       [0:0]    mul3_104_port_byte_out_0;
  wire       [0:0]    mul3_104_port_byte_out_1;
  wire       [0:0]    mul3_104_port_byte_out_2;
  wire       [0:0]    mul3_104_port_byte_out_3;
  wire       [0:0]    mul3_104_port_byte_out_4;
  wire       [0:0]    mul3_104_port_byte_out_5;
  wire       [0:0]    mul3_104_port_byte_out_6;
  wire       [0:0]    mul3_104_port_byte_out_7;
  wire       [0:0]    mul2_105_port_byte_out_0;
  wire       [0:0]    mul2_105_port_byte_out_1;
  wire       [0:0]    mul2_105_port_byte_out_2;
  wire       [0:0]    mul2_105_port_byte_out_3;
  wire       [0:0]    mul2_105_port_byte_out_4;
  wire       [0:0]    mul2_105_port_byte_out_5;
  wire       [0:0]    mul2_105_port_byte_out_6;
  wire       [0:0]    mul2_105_port_byte_out_7;
  wire       [0:0]    mul3_105_port_byte_out_0;
  wire       [0:0]    mul3_105_port_byte_out_1;
  wire       [0:0]    mul3_105_port_byte_out_2;
  wire       [0:0]    mul3_105_port_byte_out_3;
  wire       [0:0]    mul3_105_port_byte_out_4;
  wire       [0:0]    mul3_105_port_byte_out_5;
  wire       [0:0]    mul3_105_port_byte_out_6;
  wire       [0:0]    mul3_105_port_byte_out_7;
  wire       [0:0]    mul2_106_port_byte_out_0;
  wire       [0:0]    mul2_106_port_byte_out_1;
  wire       [0:0]    mul2_106_port_byte_out_2;
  wire       [0:0]    mul2_106_port_byte_out_3;
  wire       [0:0]    mul2_106_port_byte_out_4;
  wire       [0:0]    mul2_106_port_byte_out_5;
  wire       [0:0]    mul2_106_port_byte_out_6;
  wire       [0:0]    mul2_106_port_byte_out_7;
  wire       [0:0]    mul3_106_port_byte_out_0;
  wire       [0:0]    mul3_106_port_byte_out_1;
  wire       [0:0]    mul3_106_port_byte_out_2;
  wire       [0:0]    mul3_106_port_byte_out_3;
  wire       [0:0]    mul3_106_port_byte_out_4;
  wire       [0:0]    mul3_106_port_byte_out_5;
  wire       [0:0]    mul3_106_port_byte_out_6;
  wire       [0:0]    mul3_106_port_byte_out_7;
  wire       [0:0]    mul2_107_port_byte_out_0;
  wire       [0:0]    mul2_107_port_byte_out_1;
  wire       [0:0]    mul2_107_port_byte_out_2;
  wire       [0:0]    mul2_107_port_byte_out_3;
  wire       [0:0]    mul2_107_port_byte_out_4;
  wire       [0:0]    mul2_107_port_byte_out_5;
  wire       [0:0]    mul2_107_port_byte_out_6;
  wire       [0:0]    mul2_107_port_byte_out_7;
  wire       [0:0]    mul3_107_port_byte_out_0;
  wire       [0:0]    mul3_107_port_byte_out_1;
  wire       [0:0]    mul3_107_port_byte_out_2;
  wire       [0:0]    mul3_107_port_byte_out_3;
  wire       [0:0]    mul3_107_port_byte_out_4;
  wire       [0:0]    mul3_107_port_byte_out_5;
  wire       [0:0]    mul3_107_port_byte_out_6;
  wire       [0:0]    mul3_107_port_byte_out_7;
  wire       [0:0]    mul2_108_port_byte_out_0;
  wire       [0:0]    mul2_108_port_byte_out_1;
  wire       [0:0]    mul2_108_port_byte_out_2;
  wire       [0:0]    mul2_108_port_byte_out_3;
  wire       [0:0]    mul2_108_port_byte_out_4;
  wire       [0:0]    mul2_108_port_byte_out_5;
  wire       [0:0]    mul2_108_port_byte_out_6;
  wire       [0:0]    mul2_108_port_byte_out_7;
  wire       [0:0]    mul3_108_port_byte_out_0;
  wire       [0:0]    mul3_108_port_byte_out_1;
  wire       [0:0]    mul3_108_port_byte_out_2;
  wire       [0:0]    mul3_108_port_byte_out_3;
  wire       [0:0]    mul3_108_port_byte_out_4;
  wire       [0:0]    mul3_108_port_byte_out_5;
  wire       [0:0]    mul3_108_port_byte_out_6;
  wire       [0:0]    mul3_108_port_byte_out_7;
  wire       [0:0]    mul2_109_port_byte_out_0;
  wire       [0:0]    mul2_109_port_byte_out_1;
  wire       [0:0]    mul2_109_port_byte_out_2;
  wire       [0:0]    mul2_109_port_byte_out_3;
  wire       [0:0]    mul2_109_port_byte_out_4;
  wire       [0:0]    mul2_109_port_byte_out_5;
  wire       [0:0]    mul2_109_port_byte_out_6;
  wire       [0:0]    mul2_109_port_byte_out_7;
  wire       [0:0]    mul3_109_port_byte_out_0;
  wire       [0:0]    mul3_109_port_byte_out_1;
  wire       [0:0]    mul3_109_port_byte_out_2;
  wire       [0:0]    mul3_109_port_byte_out_3;
  wire       [0:0]    mul3_109_port_byte_out_4;
  wire       [0:0]    mul3_109_port_byte_out_5;
  wire       [0:0]    mul3_109_port_byte_out_6;
  wire       [0:0]    mul3_109_port_byte_out_7;
  wire       [0:0]    mul2_110_port_byte_out_0;
  wire       [0:0]    mul2_110_port_byte_out_1;
  wire       [0:0]    mul2_110_port_byte_out_2;
  wire       [0:0]    mul2_110_port_byte_out_3;
  wire       [0:0]    mul2_110_port_byte_out_4;
  wire       [0:0]    mul2_110_port_byte_out_5;
  wire       [0:0]    mul2_110_port_byte_out_6;
  wire       [0:0]    mul2_110_port_byte_out_7;
  wire       [0:0]    mul3_110_port_byte_out_0;
  wire       [0:0]    mul3_110_port_byte_out_1;
  wire       [0:0]    mul3_110_port_byte_out_2;
  wire       [0:0]    mul3_110_port_byte_out_3;
  wire       [0:0]    mul3_110_port_byte_out_4;
  wire       [0:0]    mul3_110_port_byte_out_5;
  wire       [0:0]    mul3_110_port_byte_out_6;
  wire       [0:0]    mul3_110_port_byte_out_7;
  wire       [0:0]    mul2_111_port_byte_out_0;
  wire       [0:0]    mul2_111_port_byte_out_1;
  wire       [0:0]    mul2_111_port_byte_out_2;
  wire       [0:0]    mul2_111_port_byte_out_3;
  wire       [0:0]    mul2_111_port_byte_out_4;
  wire       [0:0]    mul2_111_port_byte_out_5;
  wire       [0:0]    mul2_111_port_byte_out_6;
  wire       [0:0]    mul2_111_port_byte_out_7;
  wire       [0:0]    mul3_111_port_byte_out_0;
  wire       [0:0]    mul3_111_port_byte_out_1;
  wire       [0:0]    mul3_111_port_byte_out_2;
  wire       [0:0]    mul3_111_port_byte_out_3;
  wire       [0:0]    mul3_111_port_byte_out_4;
  wire       [0:0]    mul3_111_port_byte_out_5;
  wire       [0:0]    mul3_111_port_byte_out_6;
  wire       [0:0]    mul3_111_port_byte_out_7;
  wire       [0:0]    mul2_112_port_byte_out_0;
  wire       [0:0]    mul2_112_port_byte_out_1;
  wire       [0:0]    mul2_112_port_byte_out_2;
  wire       [0:0]    mul2_112_port_byte_out_3;
  wire       [0:0]    mul2_112_port_byte_out_4;
  wire       [0:0]    mul2_112_port_byte_out_5;
  wire       [0:0]    mul2_112_port_byte_out_6;
  wire       [0:0]    mul2_112_port_byte_out_7;
  wire       [0:0]    mul3_112_port_byte_out_0;
  wire       [0:0]    mul3_112_port_byte_out_1;
  wire       [0:0]    mul3_112_port_byte_out_2;
  wire       [0:0]    mul3_112_port_byte_out_3;
  wire       [0:0]    mul3_112_port_byte_out_4;
  wire       [0:0]    mul3_112_port_byte_out_5;
  wire       [0:0]    mul3_112_port_byte_out_6;
  wire       [0:0]    mul3_112_port_byte_out_7;
  wire       [0:0]    mul2_113_port_byte_out_0;
  wire       [0:0]    mul2_113_port_byte_out_1;
  wire       [0:0]    mul2_113_port_byte_out_2;
  wire       [0:0]    mul2_113_port_byte_out_3;
  wire       [0:0]    mul2_113_port_byte_out_4;
  wire       [0:0]    mul2_113_port_byte_out_5;
  wire       [0:0]    mul2_113_port_byte_out_6;
  wire       [0:0]    mul2_113_port_byte_out_7;
  wire       [0:0]    mul3_113_port_byte_out_0;
  wire       [0:0]    mul3_113_port_byte_out_1;
  wire       [0:0]    mul3_113_port_byte_out_2;
  wire       [0:0]    mul3_113_port_byte_out_3;
  wire       [0:0]    mul3_113_port_byte_out_4;
  wire       [0:0]    mul3_113_port_byte_out_5;
  wire       [0:0]    mul3_113_port_byte_out_6;
  wire       [0:0]    mul3_113_port_byte_out_7;
  wire       [0:0]    mul2_114_port_byte_out_0;
  wire       [0:0]    mul2_114_port_byte_out_1;
  wire       [0:0]    mul2_114_port_byte_out_2;
  wire       [0:0]    mul2_114_port_byte_out_3;
  wire       [0:0]    mul2_114_port_byte_out_4;
  wire       [0:0]    mul2_114_port_byte_out_5;
  wire       [0:0]    mul2_114_port_byte_out_6;
  wire       [0:0]    mul2_114_port_byte_out_7;
  wire       [0:0]    mul3_114_port_byte_out_0;
  wire       [0:0]    mul3_114_port_byte_out_1;
  wire       [0:0]    mul3_114_port_byte_out_2;
  wire       [0:0]    mul3_114_port_byte_out_3;
  wire       [0:0]    mul3_114_port_byte_out_4;
  wire       [0:0]    mul3_114_port_byte_out_5;
  wire       [0:0]    mul3_114_port_byte_out_6;
  wire       [0:0]    mul3_114_port_byte_out_7;
  wire       [0:0]    mul2_115_port_byte_out_0;
  wire       [0:0]    mul2_115_port_byte_out_1;
  wire       [0:0]    mul2_115_port_byte_out_2;
  wire       [0:0]    mul2_115_port_byte_out_3;
  wire       [0:0]    mul2_115_port_byte_out_4;
  wire       [0:0]    mul2_115_port_byte_out_5;
  wire       [0:0]    mul2_115_port_byte_out_6;
  wire       [0:0]    mul2_115_port_byte_out_7;
  wire       [0:0]    mul3_115_port_byte_out_0;
  wire       [0:0]    mul3_115_port_byte_out_1;
  wire       [0:0]    mul3_115_port_byte_out_2;
  wire       [0:0]    mul3_115_port_byte_out_3;
  wire       [0:0]    mul3_115_port_byte_out_4;
  wire       [0:0]    mul3_115_port_byte_out_5;
  wire       [0:0]    mul3_115_port_byte_out_6;
  wire       [0:0]    mul3_115_port_byte_out_7;
  wire       [0:0]    mul2_116_port_byte_out_0;
  wire       [0:0]    mul2_116_port_byte_out_1;
  wire       [0:0]    mul2_116_port_byte_out_2;
  wire       [0:0]    mul2_116_port_byte_out_3;
  wire       [0:0]    mul2_116_port_byte_out_4;
  wire       [0:0]    mul2_116_port_byte_out_5;
  wire       [0:0]    mul2_116_port_byte_out_6;
  wire       [0:0]    mul2_116_port_byte_out_7;
  wire       [0:0]    mul3_116_port_byte_out_0;
  wire       [0:0]    mul3_116_port_byte_out_1;
  wire       [0:0]    mul3_116_port_byte_out_2;
  wire       [0:0]    mul3_116_port_byte_out_3;
  wire       [0:0]    mul3_116_port_byte_out_4;
  wire       [0:0]    mul3_116_port_byte_out_5;
  wire       [0:0]    mul3_116_port_byte_out_6;
  wire       [0:0]    mul3_116_port_byte_out_7;
  wire       [0:0]    mul2_117_port_byte_out_0;
  wire       [0:0]    mul2_117_port_byte_out_1;
  wire       [0:0]    mul2_117_port_byte_out_2;
  wire       [0:0]    mul2_117_port_byte_out_3;
  wire       [0:0]    mul2_117_port_byte_out_4;
  wire       [0:0]    mul2_117_port_byte_out_5;
  wire       [0:0]    mul2_117_port_byte_out_6;
  wire       [0:0]    mul2_117_port_byte_out_7;
  wire       [0:0]    mul3_117_port_byte_out_0;
  wire       [0:0]    mul3_117_port_byte_out_1;
  wire       [0:0]    mul3_117_port_byte_out_2;
  wire       [0:0]    mul3_117_port_byte_out_3;
  wire       [0:0]    mul3_117_port_byte_out_4;
  wire       [0:0]    mul3_117_port_byte_out_5;
  wire       [0:0]    mul3_117_port_byte_out_6;
  wire       [0:0]    mul3_117_port_byte_out_7;
  wire       [0:0]    mul2_118_port_byte_out_0;
  wire       [0:0]    mul2_118_port_byte_out_1;
  wire       [0:0]    mul2_118_port_byte_out_2;
  wire       [0:0]    mul2_118_port_byte_out_3;
  wire       [0:0]    mul2_118_port_byte_out_4;
  wire       [0:0]    mul2_118_port_byte_out_5;
  wire       [0:0]    mul2_118_port_byte_out_6;
  wire       [0:0]    mul2_118_port_byte_out_7;
  wire       [0:0]    mul3_118_port_byte_out_0;
  wire       [0:0]    mul3_118_port_byte_out_1;
  wire       [0:0]    mul3_118_port_byte_out_2;
  wire       [0:0]    mul3_118_port_byte_out_3;
  wire       [0:0]    mul3_118_port_byte_out_4;
  wire       [0:0]    mul3_118_port_byte_out_5;
  wire       [0:0]    mul3_118_port_byte_out_6;
  wire       [0:0]    mul3_118_port_byte_out_7;
  wire       [0:0]    mul2_119_port_byte_out_0;
  wire       [0:0]    mul2_119_port_byte_out_1;
  wire       [0:0]    mul2_119_port_byte_out_2;
  wire       [0:0]    mul2_119_port_byte_out_3;
  wire       [0:0]    mul2_119_port_byte_out_4;
  wire       [0:0]    mul2_119_port_byte_out_5;
  wire       [0:0]    mul2_119_port_byte_out_6;
  wire       [0:0]    mul2_119_port_byte_out_7;
  wire       [0:0]    mul3_119_port_byte_out_0;
  wire       [0:0]    mul3_119_port_byte_out_1;
  wire       [0:0]    mul3_119_port_byte_out_2;
  wire       [0:0]    mul3_119_port_byte_out_3;
  wire       [0:0]    mul3_119_port_byte_out_4;
  wire       [0:0]    mul3_119_port_byte_out_5;
  wire       [0:0]    mul3_119_port_byte_out_6;
  wire       [0:0]    mul3_119_port_byte_out_7;
  wire       [0:0]    mul2_120_port_byte_out_0;
  wire       [0:0]    mul2_120_port_byte_out_1;
  wire       [0:0]    mul2_120_port_byte_out_2;
  wire       [0:0]    mul2_120_port_byte_out_3;
  wire       [0:0]    mul2_120_port_byte_out_4;
  wire       [0:0]    mul2_120_port_byte_out_5;
  wire       [0:0]    mul2_120_port_byte_out_6;
  wire       [0:0]    mul2_120_port_byte_out_7;
  wire       [0:0]    mul3_120_port_byte_out_0;
  wire       [0:0]    mul3_120_port_byte_out_1;
  wire       [0:0]    mul3_120_port_byte_out_2;
  wire       [0:0]    mul3_120_port_byte_out_3;
  wire       [0:0]    mul3_120_port_byte_out_4;
  wire       [0:0]    mul3_120_port_byte_out_5;
  wire       [0:0]    mul3_120_port_byte_out_6;
  wire       [0:0]    mul3_120_port_byte_out_7;
  wire       [0:0]    mul2_121_port_byte_out_0;
  wire       [0:0]    mul2_121_port_byte_out_1;
  wire       [0:0]    mul2_121_port_byte_out_2;
  wire       [0:0]    mul2_121_port_byte_out_3;
  wire       [0:0]    mul2_121_port_byte_out_4;
  wire       [0:0]    mul2_121_port_byte_out_5;
  wire       [0:0]    mul2_121_port_byte_out_6;
  wire       [0:0]    mul2_121_port_byte_out_7;
  wire       [0:0]    mul3_121_port_byte_out_0;
  wire       [0:0]    mul3_121_port_byte_out_1;
  wire       [0:0]    mul3_121_port_byte_out_2;
  wire       [0:0]    mul3_121_port_byte_out_3;
  wire       [0:0]    mul3_121_port_byte_out_4;
  wire       [0:0]    mul3_121_port_byte_out_5;
  wire       [0:0]    mul3_121_port_byte_out_6;
  wire       [0:0]    mul3_121_port_byte_out_7;
  wire       [0:0]    mul2_122_port_byte_out_0;
  wire       [0:0]    mul2_122_port_byte_out_1;
  wire       [0:0]    mul2_122_port_byte_out_2;
  wire       [0:0]    mul2_122_port_byte_out_3;
  wire       [0:0]    mul2_122_port_byte_out_4;
  wire       [0:0]    mul2_122_port_byte_out_5;
  wire       [0:0]    mul2_122_port_byte_out_6;
  wire       [0:0]    mul2_122_port_byte_out_7;
  wire       [0:0]    mul3_122_port_byte_out_0;
  wire       [0:0]    mul3_122_port_byte_out_1;
  wire       [0:0]    mul3_122_port_byte_out_2;
  wire       [0:0]    mul3_122_port_byte_out_3;
  wire       [0:0]    mul3_122_port_byte_out_4;
  wire       [0:0]    mul3_122_port_byte_out_5;
  wire       [0:0]    mul3_122_port_byte_out_6;
  wire       [0:0]    mul3_122_port_byte_out_7;
  wire       [0:0]    mul2_123_port_byte_out_0;
  wire       [0:0]    mul2_123_port_byte_out_1;
  wire       [0:0]    mul2_123_port_byte_out_2;
  wire       [0:0]    mul2_123_port_byte_out_3;
  wire       [0:0]    mul2_123_port_byte_out_4;
  wire       [0:0]    mul2_123_port_byte_out_5;
  wire       [0:0]    mul2_123_port_byte_out_6;
  wire       [0:0]    mul2_123_port_byte_out_7;
  wire       [0:0]    mul3_123_port_byte_out_0;
  wire       [0:0]    mul3_123_port_byte_out_1;
  wire       [0:0]    mul3_123_port_byte_out_2;
  wire       [0:0]    mul3_123_port_byte_out_3;
  wire       [0:0]    mul3_123_port_byte_out_4;
  wire       [0:0]    mul3_123_port_byte_out_5;
  wire       [0:0]    mul3_123_port_byte_out_6;
  wire       [0:0]    mul3_123_port_byte_out_7;
  wire       [0:0]    mul2_124_port_byte_out_0;
  wire       [0:0]    mul2_124_port_byte_out_1;
  wire       [0:0]    mul2_124_port_byte_out_2;
  wire       [0:0]    mul2_124_port_byte_out_3;
  wire       [0:0]    mul2_124_port_byte_out_4;
  wire       [0:0]    mul2_124_port_byte_out_5;
  wire       [0:0]    mul2_124_port_byte_out_6;
  wire       [0:0]    mul2_124_port_byte_out_7;
  wire       [0:0]    mul3_124_port_byte_out_0;
  wire       [0:0]    mul3_124_port_byte_out_1;
  wire       [0:0]    mul3_124_port_byte_out_2;
  wire       [0:0]    mul3_124_port_byte_out_3;
  wire       [0:0]    mul3_124_port_byte_out_4;
  wire       [0:0]    mul3_124_port_byte_out_5;
  wire       [0:0]    mul3_124_port_byte_out_6;
  wire       [0:0]    mul3_124_port_byte_out_7;
  wire       [0:0]    mul2_125_port_byte_out_0;
  wire       [0:0]    mul2_125_port_byte_out_1;
  wire       [0:0]    mul2_125_port_byte_out_2;
  wire       [0:0]    mul2_125_port_byte_out_3;
  wire       [0:0]    mul2_125_port_byte_out_4;
  wire       [0:0]    mul2_125_port_byte_out_5;
  wire       [0:0]    mul2_125_port_byte_out_6;
  wire       [0:0]    mul2_125_port_byte_out_7;
  wire       [0:0]    mul3_125_port_byte_out_0;
  wire       [0:0]    mul3_125_port_byte_out_1;
  wire       [0:0]    mul3_125_port_byte_out_2;
  wire       [0:0]    mul3_125_port_byte_out_3;
  wire       [0:0]    mul3_125_port_byte_out_4;
  wire       [0:0]    mul3_125_port_byte_out_5;
  wire       [0:0]    mul3_125_port_byte_out_6;
  wire       [0:0]    mul3_125_port_byte_out_7;
  wire       [0:0]    mul2_126_port_byte_out_0;
  wire       [0:0]    mul2_126_port_byte_out_1;
  wire       [0:0]    mul2_126_port_byte_out_2;
  wire       [0:0]    mul2_126_port_byte_out_3;
  wire       [0:0]    mul2_126_port_byte_out_4;
  wire       [0:0]    mul2_126_port_byte_out_5;
  wire       [0:0]    mul2_126_port_byte_out_6;
  wire       [0:0]    mul2_126_port_byte_out_7;
  wire       [0:0]    mul3_126_port_byte_out_0;
  wire       [0:0]    mul3_126_port_byte_out_1;
  wire       [0:0]    mul3_126_port_byte_out_2;
  wire       [0:0]    mul3_126_port_byte_out_3;
  wire       [0:0]    mul3_126_port_byte_out_4;
  wire       [0:0]    mul3_126_port_byte_out_5;
  wire       [0:0]    mul3_126_port_byte_out_6;
  wire       [0:0]    mul3_126_port_byte_out_7;
  wire       [0:0]    mul2_127_port_byte_out_0;
  wire       [0:0]    mul2_127_port_byte_out_1;
  wire       [0:0]    mul2_127_port_byte_out_2;
  wire       [0:0]    mul2_127_port_byte_out_3;
  wire       [0:0]    mul2_127_port_byte_out_4;
  wire       [0:0]    mul2_127_port_byte_out_5;
  wire       [0:0]    mul2_127_port_byte_out_6;
  wire       [0:0]    mul2_127_port_byte_out_7;
  wire       [0:0]    mul3_127_port_byte_out_0;
  wire       [0:0]    mul3_127_port_byte_out_1;
  wire       [0:0]    mul3_127_port_byte_out_2;
  wire       [0:0]    mul3_127_port_byte_out_3;
  wire       [0:0]    mul3_127_port_byte_out_4;
  wire       [0:0]    mul3_127_port_byte_out_5;
  wire       [0:0]    mul3_127_port_byte_out_6;
  wire       [0:0]    mul3_127_port_byte_out_7;
  wire       [0:0]    state_out_0_0_0;
  wire       [0:0]    state_out_0_0_1;
  wire       [0:0]    state_out_0_0_2;
  wire       [0:0]    state_out_0_0_3;
  wire       [0:0]    state_out_0_0_4;
  wire       [0:0]    state_out_0_0_5;
  wire       [0:0]    state_out_0_0_6;
  wire       [0:0]    state_out_0_0_7;
  wire       [0:0]    state_out_0_1_0;
  wire       [0:0]    state_out_0_1_1;
  wire       [0:0]    state_out_0_1_2;
  wire       [0:0]    state_out_0_1_3;
  wire       [0:0]    state_out_0_1_4;
  wire       [0:0]    state_out_0_1_5;
  wire       [0:0]    state_out_0_1_6;
  wire       [0:0]    state_out_0_1_7;
  wire       [0:0]    state_out_0_2_0;
  wire       [0:0]    state_out_0_2_1;
  wire       [0:0]    state_out_0_2_2;
  wire       [0:0]    state_out_0_2_3;
  wire       [0:0]    state_out_0_2_4;
  wire       [0:0]    state_out_0_2_5;
  wire       [0:0]    state_out_0_2_6;
  wire       [0:0]    state_out_0_2_7;
  wire       [0:0]    state_out_0_3_0;
  wire       [0:0]    state_out_0_3_1;
  wire       [0:0]    state_out_0_3_2;
  wire       [0:0]    state_out_0_3_3;
  wire       [0:0]    state_out_0_3_4;
  wire       [0:0]    state_out_0_3_5;
  wire       [0:0]    state_out_0_3_6;
  wire       [0:0]    state_out_0_3_7;
  wire       [0:0]    state_out_1_0_0;
  wire       [0:0]    state_out_1_0_1;
  wire       [0:0]    state_out_1_0_2;
  wire       [0:0]    state_out_1_0_3;
  wire       [0:0]    state_out_1_0_4;
  wire       [0:0]    state_out_1_0_5;
  wire       [0:0]    state_out_1_0_6;
  wire       [0:0]    state_out_1_0_7;
  wire       [0:0]    state_out_1_1_0;
  wire       [0:0]    state_out_1_1_1;
  wire       [0:0]    state_out_1_1_2;
  wire       [0:0]    state_out_1_1_3;
  wire       [0:0]    state_out_1_1_4;
  wire       [0:0]    state_out_1_1_5;
  wire       [0:0]    state_out_1_1_6;
  wire       [0:0]    state_out_1_1_7;
  wire       [0:0]    state_out_1_2_0;
  wire       [0:0]    state_out_1_2_1;
  wire       [0:0]    state_out_1_2_2;
  wire       [0:0]    state_out_1_2_3;
  wire       [0:0]    state_out_1_2_4;
  wire       [0:0]    state_out_1_2_5;
  wire       [0:0]    state_out_1_2_6;
  wire       [0:0]    state_out_1_2_7;
  wire       [0:0]    state_out_1_3_0;
  wire       [0:0]    state_out_1_3_1;
  wire       [0:0]    state_out_1_3_2;
  wire       [0:0]    state_out_1_3_3;
  wire       [0:0]    state_out_1_3_4;
  wire       [0:0]    state_out_1_3_5;
  wire       [0:0]    state_out_1_3_6;
  wire       [0:0]    state_out_1_3_7;
  wire       [0:0]    state_out_2_0_0;
  wire       [0:0]    state_out_2_0_1;
  wire       [0:0]    state_out_2_0_2;
  wire       [0:0]    state_out_2_0_3;
  wire       [0:0]    state_out_2_0_4;
  wire       [0:0]    state_out_2_0_5;
  wire       [0:0]    state_out_2_0_6;
  wire       [0:0]    state_out_2_0_7;
  wire       [0:0]    state_out_2_1_0;
  wire       [0:0]    state_out_2_1_1;
  wire       [0:0]    state_out_2_1_2;
  wire       [0:0]    state_out_2_1_3;
  wire       [0:0]    state_out_2_1_4;
  wire       [0:0]    state_out_2_1_5;
  wire       [0:0]    state_out_2_1_6;
  wire       [0:0]    state_out_2_1_7;
  wire       [0:0]    state_out_2_2_0;
  wire       [0:0]    state_out_2_2_1;
  wire       [0:0]    state_out_2_2_2;
  wire       [0:0]    state_out_2_2_3;
  wire       [0:0]    state_out_2_2_4;
  wire       [0:0]    state_out_2_2_5;
  wire       [0:0]    state_out_2_2_6;
  wire       [0:0]    state_out_2_2_7;
  wire       [0:0]    state_out_2_3_0;
  wire       [0:0]    state_out_2_3_1;
  wire       [0:0]    state_out_2_3_2;
  wire       [0:0]    state_out_2_3_3;
  wire       [0:0]    state_out_2_3_4;
  wire       [0:0]    state_out_2_3_5;
  wire       [0:0]    state_out_2_3_6;
  wire       [0:0]    state_out_2_3_7;
  wire       [0:0]    state_out_3_0_0;
  wire       [0:0]    state_out_3_0_1;
  wire       [0:0]    state_out_3_0_2;
  wire       [0:0]    state_out_3_0_3;
  wire       [0:0]    state_out_3_0_4;
  wire       [0:0]    state_out_3_0_5;
  wire       [0:0]    state_out_3_0_6;
  wire       [0:0]    state_out_3_0_7;
  wire       [0:0]    state_out_3_1_0;
  wire       [0:0]    state_out_3_1_1;
  wire       [0:0]    state_out_3_1_2;
  wire       [0:0]    state_out_3_1_3;
  wire       [0:0]    state_out_3_1_4;
  wire       [0:0]    state_out_3_1_5;
  wire       [0:0]    state_out_3_1_6;
  wire       [0:0]    state_out_3_1_7;
  wire       [0:0]    state_out_3_2_0;
  wire       [0:0]    state_out_3_2_1;
  wire       [0:0]    state_out_3_2_2;
  wire       [0:0]    state_out_3_2_3;
  wire       [0:0]    state_out_3_2_4;
  wire       [0:0]    state_out_3_2_5;
  wire       [0:0]    state_out_3_2_6;
  wire       [0:0]    state_out_3_2_7;
  wire       [0:0]    state_out_3_3_0;
  wire       [0:0]    state_out_3_3_1;
  wire       [0:0]    state_out_3_3_2;
  wire       [0:0]    state_out_3_3_3;
  wire       [0:0]    state_out_3_3_4;
  wire       [0:0]    state_out_3_3_5;
  wire       [0:0]    state_out_3_3_6;
  wire       [0:0]    state_out_3_3_7;
  wire       [0:0]    state_out_4_0_0;
  wire       [0:0]    state_out_4_0_1;
  wire       [0:0]    state_out_4_0_2;
  wire       [0:0]    state_out_4_0_3;
  wire       [0:0]    state_out_4_0_4;
  wire       [0:0]    state_out_4_0_5;
  wire       [0:0]    state_out_4_0_6;
  wire       [0:0]    state_out_4_0_7;
  wire       [0:0]    state_out_4_1_0;
  wire       [0:0]    state_out_4_1_1;
  wire       [0:0]    state_out_4_1_2;
  wire       [0:0]    state_out_4_1_3;
  wire       [0:0]    state_out_4_1_4;
  wire       [0:0]    state_out_4_1_5;
  wire       [0:0]    state_out_4_1_6;
  wire       [0:0]    state_out_4_1_7;
  wire       [0:0]    state_out_4_2_0;
  wire       [0:0]    state_out_4_2_1;
  wire       [0:0]    state_out_4_2_2;
  wire       [0:0]    state_out_4_2_3;
  wire       [0:0]    state_out_4_2_4;
  wire       [0:0]    state_out_4_2_5;
  wire       [0:0]    state_out_4_2_6;
  wire       [0:0]    state_out_4_2_7;
  wire       [0:0]    state_out_4_3_0;
  wire       [0:0]    state_out_4_3_1;
  wire       [0:0]    state_out_4_3_2;
  wire       [0:0]    state_out_4_3_3;
  wire       [0:0]    state_out_4_3_4;
  wire       [0:0]    state_out_4_3_5;
  wire       [0:0]    state_out_4_3_6;
  wire       [0:0]    state_out_4_3_7;
  wire       [0:0]    state_out_5_0_0;
  wire       [0:0]    state_out_5_0_1;
  wire       [0:0]    state_out_5_0_2;
  wire       [0:0]    state_out_5_0_3;
  wire       [0:0]    state_out_5_0_4;
  wire       [0:0]    state_out_5_0_5;
  wire       [0:0]    state_out_5_0_6;
  wire       [0:0]    state_out_5_0_7;
  wire       [0:0]    state_out_5_1_0;
  wire       [0:0]    state_out_5_1_1;
  wire       [0:0]    state_out_5_1_2;
  wire       [0:0]    state_out_5_1_3;
  wire       [0:0]    state_out_5_1_4;
  wire       [0:0]    state_out_5_1_5;
  wire       [0:0]    state_out_5_1_6;
  wire       [0:0]    state_out_5_1_7;
  wire       [0:0]    state_out_5_2_0;
  wire       [0:0]    state_out_5_2_1;
  wire       [0:0]    state_out_5_2_2;
  wire       [0:0]    state_out_5_2_3;
  wire       [0:0]    state_out_5_2_4;
  wire       [0:0]    state_out_5_2_5;
  wire       [0:0]    state_out_5_2_6;
  wire       [0:0]    state_out_5_2_7;
  wire       [0:0]    state_out_5_3_0;
  wire       [0:0]    state_out_5_3_1;
  wire       [0:0]    state_out_5_3_2;
  wire       [0:0]    state_out_5_3_3;
  wire       [0:0]    state_out_5_3_4;
  wire       [0:0]    state_out_5_3_5;
  wire       [0:0]    state_out_5_3_6;
  wire       [0:0]    state_out_5_3_7;
  wire       [0:0]    state_out_6_0_0;
  wire       [0:0]    state_out_6_0_1;
  wire       [0:0]    state_out_6_0_2;
  wire       [0:0]    state_out_6_0_3;
  wire       [0:0]    state_out_6_0_4;
  wire       [0:0]    state_out_6_0_5;
  wire       [0:0]    state_out_6_0_6;
  wire       [0:0]    state_out_6_0_7;
  wire       [0:0]    state_out_6_1_0;
  wire       [0:0]    state_out_6_1_1;
  wire       [0:0]    state_out_6_1_2;
  wire       [0:0]    state_out_6_1_3;
  wire       [0:0]    state_out_6_1_4;
  wire       [0:0]    state_out_6_1_5;
  wire       [0:0]    state_out_6_1_6;
  wire       [0:0]    state_out_6_1_7;
  wire       [0:0]    state_out_6_2_0;
  wire       [0:0]    state_out_6_2_1;
  wire       [0:0]    state_out_6_2_2;
  wire       [0:0]    state_out_6_2_3;
  wire       [0:0]    state_out_6_2_4;
  wire       [0:0]    state_out_6_2_5;
  wire       [0:0]    state_out_6_2_6;
  wire       [0:0]    state_out_6_2_7;
  wire       [0:0]    state_out_6_3_0;
  wire       [0:0]    state_out_6_3_1;
  wire       [0:0]    state_out_6_3_2;
  wire       [0:0]    state_out_6_3_3;
  wire       [0:0]    state_out_6_3_4;
  wire       [0:0]    state_out_6_3_5;
  wire       [0:0]    state_out_6_3_6;
  wire       [0:0]    state_out_6_3_7;
  wire       [0:0]    state_out_7_0_0;
  wire       [0:0]    state_out_7_0_1;
  wire       [0:0]    state_out_7_0_2;
  wire       [0:0]    state_out_7_0_3;
  wire       [0:0]    state_out_7_0_4;
  wire       [0:0]    state_out_7_0_5;
  wire       [0:0]    state_out_7_0_6;
  wire       [0:0]    state_out_7_0_7;
  wire       [0:0]    state_out_7_1_0;
  wire       [0:0]    state_out_7_1_1;
  wire       [0:0]    state_out_7_1_2;
  wire       [0:0]    state_out_7_1_3;
  wire       [0:0]    state_out_7_1_4;
  wire       [0:0]    state_out_7_1_5;
  wire       [0:0]    state_out_7_1_6;
  wire       [0:0]    state_out_7_1_7;
  wire       [0:0]    state_out_7_2_0;
  wire       [0:0]    state_out_7_2_1;
  wire       [0:0]    state_out_7_2_2;
  wire       [0:0]    state_out_7_2_3;
  wire       [0:0]    state_out_7_2_4;
  wire       [0:0]    state_out_7_2_5;
  wire       [0:0]    state_out_7_2_6;
  wire       [0:0]    state_out_7_2_7;
  wire       [0:0]    state_out_7_3_0;
  wire       [0:0]    state_out_7_3_1;
  wire       [0:0]    state_out_7_3_2;
  wire       [0:0]    state_out_7_3_3;
  wire       [0:0]    state_out_7_3_4;
  wire       [0:0]    state_out_7_3_5;
  wire       [0:0]    state_out_7_3_6;
  wire       [0:0]    state_out_7_3_7;
  wire       [0:0]    state_out_8_0_0;
  wire       [0:0]    state_out_8_0_1;
  wire       [0:0]    state_out_8_0_2;
  wire       [0:0]    state_out_8_0_3;
  wire       [0:0]    state_out_8_0_4;
  wire       [0:0]    state_out_8_0_5;
  wire       [0:0]    state_out_8_0_6;
  wire       [0:0]    state_out_8_0_7;
  wire       [0:0]    state_out_8_1_0;
  wire       [0:0]    state_out_8_1_1;
  wire       [0:0]    state_out_8_1_2;
  wire       [0:0]    state_out_8_1_3;
  wire       [0:0]    state_out_8_1_4;
  wire       [0:0]    state_out_8_1_5;
  wire       [0:0]    state_out_8_1_6;
  wire       [0:0]    state_out_8_1_7;
  wire       [0:0]    state_out_8_2_0;
  wire       [0:0]    state_out_8_2_1;
  wire       [0:0]    state_out_8_2_2;
  wire       [0:0]    state_out_8_2_3;
  wire       [0:0]    state_out_8_2_4;
  wire       [0:0]    state_out_8_2_5;
  wire       [0:0]    state_out_8_2_6;
  wire       [0:0]    state_out_8_2_7;
  wire       [0:0]    state_out_8_3_0;
  wire       [0:0]    state_out_8_3_1;
  wire       [0:0]    state_out_8_3_2;
  wire       [0:0]    state_out_8_3_3;
  wire       [0:0]    state_out_8_3_4;
  wire       [0:0]    state_out_8_3_5;
  wire       [0:0]    state_out_8_3_6;
  wire       [0:0]    state_out_8_3_7;
  wire       [0:0]    state_out_9_0_0;
  wire       [0:0]    state_out_9_0_1;
  wire       [0:0]    state_out_9_0_2;
  wire       [0:0]    state_out_9_0_3;
  wire       [0:0]    state_out_9_0_4;
  wire       [0:0]    state_out_9_0_5;
  wire       [0:0]    state_out_9_0_6;
  wire       [0:0]    state_out_9_0_7;
  wire       [0:0]    state_out_9_1_0;
  wire       [0:0]    state_out_9_1_1;
  wire       [0:0]    state_out_9_1_2;
  wire       [0:0]    state_out_9_1_3;
  wire       [0:0]    state_out_9_1_4;
  wire       [0:0]    state_out_9_1_5;
  wire       [0:0]    state_out_9_1_6;
  wire       [0:0]    state_out_9_1_7;
  wire       [0:0]    state_out_9_2_0;
  wire       [0:0]    state_out_9_2_1;
  wire       [0:0]    state_out_9_2_2;
  wire       [0:0]    state_out_9_2_3;
  wire       [0:0]    state_out_9_2_4;
  wire       [0:0]    state_out_9_2_5;
  wire       [0:0]    state_out_9_2_6;
  wire       [0:0]    state_out_9_2_7;
  wire       [0:0]    state_out_9_3_0;
  wire       [0:0]    state_out_9_3_1;
  wire       [0:0]    state_out_9_3_2;
  wire       [0:0]    state_out_9_3_3;
  wire       [0:0]    state_out_9_3_4;
  wire       [0:0]    state_out_9_3_5;
  wire       [0:0]    state_out_9_3_6;
  wire       [0:0]    state_out_9_3_7;
  wire       [0:0]    state_out_10_0_0;
  wire       [0:0]    state_out_10_0_1;
  wire       [0:0]    state_out_10_0_2;
  wire       [0:0]    state_out_10_0_3;
  wire       [0:0]    state_out_10_0_4;
  wire       [0:0]    state_out_10_0_5;
  wire       [0:0]    state_out_10_0_6;
  wire       [0:0]    state_out_10_0_7;
  wire       [0:0]    state_out_10_1_0;
  wire       [0:0]    state_out_10_1_1;
  wire       [0:0]    state_out_10_1_2;
  wire       [0:0]    state_out_10_1_3;
  wire       [0:0]    state_out_10_1_4;
  wire       [0:0]    state_out_10_1_5;
  wire       [0:0]    state_out_10_1_6;
  wire       [0:0]    state_out_10_1_7;
  wire       [0:0]    state_out_10_2_0;
  wire       [0:0]    state_out_10_2_1;
  wire       [0:0]    state_out_10_2_2;
  wire       [0:0]    state_out_10_2_3;
  wire       [0:0]    state_out_10_2_4;
  wire       [0:0]    state_out_10_2_5;
  wire       [0:0]    state_out_10_2_6;
  wire       [0:0]    state_out_10_2_7;
  wire       [0:0]    state_out_10_3_0;
  wire       [0:0]    state_out_10_3_1;
  wire       [0:0]    state_out_10_3_2;
  wire       [0:0]    state_out_10_3_3;
  wire       [0:0]    state_out_10_3_4;
  wire       [0:0]    state_out_10_3_5;
  wire       [0:0]    state_out_10_3_6;
  wire       [0:0]    state_out_10_3_7;
  wire       [0:0]    state_out_11_0_0;
  wire       [0:0]    state_out_11_0_1;
  wire       [0:0]    state_out_11_0_2;
  wire       [0:0]    state_out_11_0_3;
  wire       [0:0]    state_out_11_0_4;
  wire       [0:0]    state_out_11_0_5;
  wire       [0:0]    state_out_11_0_6;
  wire       [0:0]    state_out_11_0_7;
  wire       [0:0]    state_out_11_1_0;
  wire       [0:0]    state_out_11_1_1;
  wire       [0:0]    state_out_11_1_2;
  wire       [0:0]    state_out_11_1_3;
  wire       [0:0]    state_out_11_1_4;
  wire       [0:0]    state_out_11_1_5;
  wire       [0:0]    state_out_11_1_6;
  wire       [0:0]    state_out_11_1_7;
  wire       [0:0]    state_out_11_2_0;
  wire       [0:0]    state_out_11_2_1;
  wire       [0:0]    state_out_11_2_2;
  wire       [0:0]    state_out_11_2_3;
  wire       [0:0]    state_out_11_2_4;
  wire       [0:0]    state_out_11_2_5;
  wire       [0:0]    state_out_11_2_6;
  wire       [0:0]    state_out_11_2_7;
  wire       [0:0]    state_out_11_3_0;
  wire       [0:0]    state_out_11_3_1;
  wire       [0:0]    state_out_11_3_2;
  wire       [0:0]    state_out_11_3_3;
  wire       [0:0]    state_out_11_3_4;
  wire       [0:0]    state_out_11_3_5;
  wire       [0:0]    state_out_11_3_6;
  wire       [0:0]    state_out_11_3_7;
  wire       [0:0]    state_out_12_0_0;
  wire       [0:0]    state_out_12_0_1;
  wire       [0:0]    state_out_12_0_2;
  wire       [0:0]    state_out_12_0_3;
  wire       [0:0]    state_out_12_0_4;
  wire       [0:0]    state_out_12_0_5;
  wire       [0:0]    state_out_12_0_6;
  wire       [0:0]    state_out_12_0_7;
  wire       [0:0]    state_out_12_1_0;
  wire       [0:0]    state_out_12_1_1;
  wire       [0:0]    state_out_12_1_2;
  wire       [0:0]    state_out_12_1_3;
  wire       [0:0]    state_out_12_1_4;
  wire       [0:0]    state_out_12_1_5;
  wire       [0:0]    state_out_12_1_6;
  wire       [0:0]    state_out_12_1_7;
  wire       [0:0]    state_out_12_2_0;
  wire       [0:0]    state_out_12_2_1;
  wire       [0:0]    state_out_12_2_2;
  wire       [0:0]    state_out_12_2_3;
  wire       [0:0]    state_out_12_2_4;
  wire       [0:0]    state_out_12_2_5;
  wire       [0:0]    state_out_12_2_6;
  wire       [0:0]    state_out_12_2_7;
  wire       [0:0]    state_out_12_3_0;
  wire       [0:0]    state_out_12_3_1;
  wire       [0:0]    state_out_12_3_2;
  wire       [0:0]    state_out_12_3_3;
  wire       [0:0]    state_out_12_3_4;
  wire       [0:0]    state_out_12_3_5;
  wire       [0:0]    state_out_12_3_6;
  wire       [0:0]    state_out_12_3_7;
  wire       [0:0]    state_out_13_0_0;
  wire       [0:0]    state_out_13_0_1;
  wire       [0:0]    state_out_13_0_2;
  wire       [0:0]    state_out_13_0_3;
  wire       [0:0]    state_out_13_0_4;
  wire       [0:0]    state_out_13_0_5;
  wire       [0:0]    state_out_13_0_6;
  wire       [0:0]    state_out_13_0_7;
  wire       [0:0]    state_out_13_1_0;
  wire       [0:0]    state_out_13_1_1;
  wire       [0:0]    state_out_13_1_2;
  wire       [0:0]    state_out_13_1_3;
  wire       [0:0]    state_out_13_1_4;
  wire       [0:0]    state_out_13_1_5;
  wire       [0:0]    state_out_13_1_6;
  wire       [0:0]    state_out_13_1_7;
  wire       [0:0]    state_out_13_2_0;
  wire       [0:0]    state_out_13_2_1;
  wire       [0:0]    state_out_13_2_2;
  wire       [0:0]    state_out_13_2_3;
  wire       [0:0]    state_out_13_2_4;
  wire       [0:0]    state_out_13_2_5;
  wire       [0:0]    state_out_13_2_6;
  wire       [0:0]    state_out_13_2_7;
  wire       [0:0]    state_out_13_3_0;
  wire       [0:0]    state_out_13_3_1;
  wire       [0:0]    state_out_13_3_2;
  wire       [0:0]    state_out_13_3_3;
  wire       [0:0]    state_out_13_3_4;
  wire       [0:0]    state_out_13_3_5;
  wire       [0:0]    state_out_13_3_6;
  wire       [0:0]    state_out_13_3_7;
  wire       [0:0]    state_out_14_0_0;
  wire       [0:0]    state_out_14_0_1;
  wire       [0:0]    state_out_14_0_2;
  wire       [0:0]    state_out_14_0_3;
  wire       [0:0]    state_out_14_0_4;
  wire       [0:0]    state_out_14_0_5;
  wire       [0:0]    state_out_14_0_6;
  wire       [0:0]    state_out_14_0_7;
  wire       [0:0]    state_out_14_1_0;
  wire       [0:0]    state_out_14_1_1;
  wire       [0:0]    state_out_14_1_2;
  wire       [0:0]    state_out_14_1_3;
  wire       [0:0]    state_out_14_1_4;
  wire       [0:0]    state_out_14_1_5;
  wire       [0:0]    state_out_14_1_6;
  wire       [0:0]    state_out_14_1_7;
  wire       [0:0]    state_out_14_2_0;
  wire       [0:0]    state_out_14_2_1;
  wire       [0:0]    state_out_14_2_2;
  wire       [0:0]    state_out_14_2_3;
  wire       [0:0]    state_out_14_2_4;
  wire       [0:0]    state_out_14_2_5;
  wire       [0:0]    state_out_14_2_6;
  wire       [0:0]    state_out_14_2_7;
  wire       [0:0]    state_out_14_3_0;
  wire       [0:0]    state_out_14_3_1;
  wire       [0:0]    state_out_14_3_2;
  wire       [0:0]    state_out_14_3_3;
  wire       [0:0]    state_out_14_3_4;
  wire       [0:0]    state_out_14_3_5;
  wire       [0:0]    state_out_14_3_6;
  wire       [0:0]    state_out_14_3_7;
  wire       [0:0]    state_out_15_0_0;
  wire       [0:0]    state_out_15_0_1;
  wire       [0:0]    state_out_15_0_2;
  wire       [0:0]    state_out_15_0_3;
  wire       [0:0]    state_out_15_0_4;
  wire       [0:0]    state_out_15_0_5;
  wire       [0:0]    state_out_15_0_6;
  wire       [0:0]    state_out_15_0_7;
  wire       [0:0]    state_out_15_1_0;
  wire       [0:0]    state_out_15_1_1;
  wire       [0:0]    state_out_15_1_2;
  wire       [0:0]    state_out_15_1_3;
  wire       [0:0]    state_out_15_1_4;
  wire       [0:0]    state_out_15_1_5;
  wire       [0:0]    state_out_15_1_6;
  wire       [0:0]    state_out_15_1_7;
  wire       [0:0]    state_out_15_2_0;
  wire       [0:0]    state_out_15_2_1;
  wire       [0:0]    state_out_15_2_2;
  wire       [0:0]    state_out_15_2_3;
  wire       [0:0]    state_out_15_2_4;
  wire       [0:0]    state_out_15_2_5;
  wire       [0:0]    state_out_15_2_6;
  wire       [0:0]    state_out_15_2_7;
  wire       [0:0]    state_out_15_3_0;
  wire       [0:0]    state_out_15_3_1;
  wire       [0:0]    state_out_15_3_2;
  wire       [0:0]    state_out_15_3_3;
  wire       [0:0]    state_out_15_3_4;
  wire       [0:0]    state_out_15_3_5;
  wire       [0:0]    state_out_15_3_6;
  wire       [0:0]    state_out_15_3_7;

  Mul2 mul2_64 (
    .port_byte_in_0  (port_state_in_0_0_0    ), //i
    .port_byte_in_1  (port_state_in_0_0_1    ), //i
    .port_byte_in_2  (port_state_in_0_0_2    ), //i
    .port_byte_in_3  (port_state_in_0_0_3    ), //i
    .port_byte_in_4  (port_state_in_0_0_4    ), //i
    .port_byte_in_5  (port_state_in_0_0_5    ), //i
    .port_byte_in_6  (port_state_in_0_0_6    ), //i
    .port_byte_in_7  (port_state_in_0_0_7    ), //i
    .port_byte_out_0 (mul2_64_port_byte_out_0), //o
    .port_byte_out_1 (mul2_64_port_byte_out_1), //o
    .port_byte_out_2 (mul2_64_port_byte_out_2), //o
    .port_byte_out_3 (mul2_64_port_byte_out_3), //o
    .port_byte_out_4 (mul2_64_port_byte_out_4), //o
    .port_byte_out_5 (mul2_64_port_byte_out_5), //o
    .port_byte_out_6 (mul2_64_port_byte_out_6), //o
    .port_byte_out_7 (mul2_64_port_byte_out_7)  //o
  );
  Mul3 mul3_64 (
    .port_byte_in_0  (port_state_in_1_0_0    ), //i
    .port_byte_in_1  (port_state_in_1_0_1    ), //i
    .port_byte_in_2  (port_state_in_1_0_2    ), //i
    .port_byte_in_3  (port_state_in_1_0_3    ), //i
    .port_byte_in_4  (port_state_in_1_0_4    ), //i
    .port_byte_in_5  (port_state_in_1_0_5    ), //i
    .port_byte_in_6  (port_state_in_1_0_6    ), //i
    .port_byte_in_7  (port_state_in_1_0_7    ), //i
    .port_byte_out_0 (mul3_64_port_byte_out_0), //o
    .port_byte_out_1 (mul3_64_port_byte_out_1), //o
    .port_byte_out_2 (mul3_64_port_byte_out_2), //o
    .port_byte_out_3 (mul3_64_port_byte_out_3), //o
    .port_byte_out_4 (mul3_64_port_byte_out_4), //o
    .port_byte_out_5 (mul3_64_port_byte_out_5), //o
    .port_byte_out_6 (mul3_64_port_byte_out_6), //o
    .port_byte_out_7 (mul3_64_port_byte_out_7)  //o
  );
  Mul2 mul2_65 (
    .port_byte_in_0  (port_state_in_1_0_0    ), //i
    .port_byte_in_1  (port_state_in_1_0_1    ), //i
    .port_byte_in_2  (port_state_in_1_0_2    ), //i
    .port_byte_in_3  (port_state_in_1_0_3    ), //i
    .port_byte_in_4  (port_state_in_1_0_4    ), //i
    .port_byte_in_5  (port_state_in_1_0_5    ), //i
    .port_byte_in_6  (port_state_in_1_0_6    ), //i
    .port_byte_in_7  (port_state_in_1_0_7    ), //i
    .port_byte_out_0 (mul2_65_port_byte_out_0), //o
    .port_byte_out_1 (mul2_65_port_byte_out_1), //o
    .port_byte_out_2 (mul2_65_port_byte_out_2), //o
    .port_byte_out_3 (mul2_65_port_byte_out_3), //o
    .port_byte_out_4 (mul2_65_port_byte_out_4), //o
    .port_byte_out_5 (mul2_65_port_byte_out_5), //o
    .port_byte_out_6 (mul2_65_port_byte_out_6), //o
    .port_byte_out_7 (mul2_65_port_byte_out_7)  //o
  );
  Mul3 mul3_65 (
    .port_byte_in_0  (port_state_in_2_0_0    ), //i
    .port_byte_in_1  (port_state_in_2_0_1    ), //i
    .port_byte_in_2  (port_state_in_2_0_2    ), //i
    .port_byte_in_3  (port_state_in_2_0_3    ), //i
    .port_byte_in_4  (port_state_in_2_0_4    ), //i
    .port_byte_in_5  (port_state_in_2_0_5    ), //i
    .port_byte_in_6  (port_state_in_2_0_6    ), //i
    .port_byte_in_7  (port_state_in_2_0_7    ), //i
    .port_byte_out_0 (mul3_65_port_byte_out_0), //o
    .port_byte_out_1 (mul3_65_port_byte_out_1), //o
    .port_byte_out_2 (mul3_65_port_byte_out_2), //o
    .port_byte_out_3 (mul3_65_port_byte_out_3), //o
    .port_byte_out_4 (mul3_65_port_byte_out_4), //o
    .port_byte_out_5 (mul3_65_port_byte_out_5), //o
    .port_byte_out_6 (mul3_65_port_byte_out_6), //o
    .port_byte_out_7 (mul3_65_port_byte_out_7)  //o
  );
  Mul2 mul2_66 (
    .port_byte_in_0  (port_state_in_2_0_0    ), //i
    .port_byte_in_1  (port_state_in_2_0_1    ), //i
    .port_byte_in_2  (port_state_in_2_0_2    ), //i
    .port_byte_in_3  (port_state_in_2_0_3    ), //i
    .port_byte_in_4  (port_state_in_2_0_4    ), //i
    .port_byte_in_5  (port_state_in_2_0_5    ), //i
    .port_byte_in_6  (port_state_in_2_0_6    ), //i
    .port_byte_in_7  (port_state_in_2_0_7    ), //i
    .port_byte_out_0 (mul2_66_port_byte_out_0), //o
    .port_byte_out_1 (mul2_66_port_byte_out_1), //o
    .port_byte_out_2 (mul2_66_port_byte_out_2), //o
    .port_byte_out_3 (mul2_66_port_byte_out_3), //o
    .port_byte_out_4 (mul2_66_port_byte_out_4), //o
    .port_byte_out_5 (mul2_66_port_byte_out_5), //o
    .port_byte_out_6 (mul2_66_port_byte_out_6), //o
    .port_byte_out_7 (mul2_66_port_byte_out_7)  //o
  );
  Mul3 mul3_66 (
    .port_byte_in_0  (port_state_in_3_0_0    ), //i
    .port_byte_in_1  (port_state_in_3_0_1    ), //i
    .port_byte_in_2  (port_state_in_3_0_2    ), //i
    .port_byte_in_3  (port_state_in_3_0_3    ), //i
    .port_byte_in_4  (port_state_in_3_0_4    ), //i
    .port_byte_in_5  (port_state_in_3_0_5    ), //i
    .port_byte_in_6  (port_state_in_3_0_6    ), //i
    .port_byte_in_7  (port_state_in_3_0_7    ), //i
    .port_byte_out_0 (mul3_66_port_byte_out_0), //o
    .port_byte_out_1 (mul3_66_port_byte_out_1), //o
    .port_byte_out_2 (mul3_66_port_byte_out_2), //o
    .port_byte_out_3 (mul3_66_port_byte_out_3), //o
    .port_byte_out_4 (mul3_66_port_byte_out_4), //o
    .port_byte_out_5 (mul3_66_port_byte_out_5), //o
    .port_byte_out_6 (mul3_66_port_byte_out_6), //o
    .port_byte_out_7 (mul3_66_port_byte_out_7)  //o
  );
  Mul2 mul2_67 (
    .port_byte_in_0  (port_state_in_3_0_0    ), //i
    .port_byte_in_1  (port_state_in_3_0_1    ), //i
    .port_byte_in_2  (port_state_in_3_0_2    ), //i
    .port_byte_in_3  (port_state_in_3_0_3    ), //i
    .port_byte_in_4  (port_state_in_3_0_4    ), //i
    .port_byte_in_5  (port_state_in_3_0_5    ), //i
    .port_byte_in_6  (port_state_in_3_0_6    ), //i
    .port_byte_in_7  (port_state_in_3_0_7    ), //i
    .port_byte_out_0 (mul2_67_port_byte_out_0), //o
    .port_byte_out_1 (mul2_67_port_byte_out_1), //o
    .port_byte_out_2 (mul2_67_port_byte_out_2), //o
    .port_byte_out_3 (mul2_67_port_byte_out_3), //o
    .port_byte_out_4 (mul2_67_port_byte_out_4), //o
    .port_byte_out_5 (mul2_67_port_byte_out_5), //o
    .port_byte_out_6 (mul2_67_port_byte_out_6), //o
    .port_byte_out_7 (mul2_67_port_byte_out_7)  //o
  );
  Mul3 mul3_67 (
    .port_byte_in_0  (port_state_in_0_0_0    ), //i
    .port_byte_in_1  (port_state_in_0_0_1    ), //i
    .port_byte_in_2  (port_state_in_0_0_2    ), //i
    .port_byte_in_3  (port_state_in_0_0_3    ), //i
    .port_byte_in_4  (port_state_in_0_0_4    ), //i
    .port_byte_in_5  (port_state_in_0_0_5    ), //i
    .port_byte_in_6  (port_state_in_0_0_6    ), //i
    .port_byte_in_7  (port_state_in_0_0_7    ), //i
    .port_byte_out_0 (mul3_67_port_byte_out_0), //o
    .port_byte_out_1 (mul3_67_port_byte_out_1), //o
    .port_byte_out_2 (mul3_67_port_byte_out_2), //o
    .port_byte_out_3 (mul3_67_port_byte_out_3), //o
    .port_byte_out_4 (mul3_67_port_byte_out_4), //o
    .port_byte_out_5 (mul3_67_port_byte_out_5), //o
    .port_byte_out_6 (mul3_67_port_byte_out_6), //o
    .port_byte_out_7 (mul3_67_port_byte_out_7)  //o
  );
  Mul2 mul2_68 (
    .port_byte_in_0  (port_state_in_0_1_0    ), //i
    .port_byte_in_1  (port_state_in_0_1_1    ), //i
    .port_byte_in_2  (port_state_in_0_1_2    ), //i
    .port_byte_in_3  (port_state_in_0_1_3    ), //i
    .port_byte_in_4  (port_state_in_0_1_4    ), //i
    .port_byte_in_5  (port_state_in_0_1_5    ), //i
    .port_byte_in_6  (port_state_in_0_1_6    ), //i
    .port_byte_in_7  (port_state_in_0_1_7    ), //i
    .port_byte_out_0 (mul2_68_port_byte_out_0), //o
    .port_byte_out_1 (mul2_68_port_byte_out_1), //o
    .port_byte_out_2 (mul2_68_port_byte_out_2), //o
    .port_byte_out_3 (mul2_68_port_byte_out_3), //o
    .port_byte_out_4 (mul2_68_port_byte_out_4), //o
    .port_byte_out_5 (mul2_68_port_byte_out_5), //o
    .port_byte_out_6 (mul2_68_port_byte_out_6), //o
    .port_byte_out_7 (mul2_68_port_byte_out_7)  //o
  );
  Mul3 mul3_68 (
    .port_byte_in_0  (port_state_in_1_1_0    ), //i
    .port_byte_in_1  (port_state_in_1_1_1    ), //i
    .port_byte_in_2  (port_state_in_1_1_2    ), //i
    .port_byte_in_3  (port_state_in_1_1_3    ), //i
    .port_byte_in_4  (port_state_in_1_1_4    ), //i
    .port_byte_in_5  (port_state_in_1_1_5    ), //i
    .port_byte_in_6  (port_state_in_1_1_6    ), //i
    .port_byte_in_7  (port_state_in_1_1_7    ), //i
    .port_byte_out_0 (mul3_68_port_byte_out_0), //o
    .port_byte_out_1 (mul3_68_port_byte_out_1), //o
    .port_byte_out_2 (mul3_68_port_byte_out_2), //o
    .port_byte_out_3 (mul3_68_port_byte_out_3), //o
    .port_byte_out_4 (mul3_68_port_byte_out_4), //o
    .port_byte_out_5 (mul3_68_port_byte_out_5), //o
    .port_byte_out_6 (mul3_68_port_byte_out_6), //o
    .port_byte_out_7 (mul3_68_port_byte_out_7)  //o
  );
  Mul2 mul2_69 (
    .port_byte_in_0  (port_state_in_1_1_0    ), //i
    .port_byte_in_1  (port_state_in_1_1_1    ), //i
    .port_byte_in_2  (port_state_in_1_1_2    ), //i
    .port_byte_in_3  (port_state_in_1_1_3    ), //i
    .port_byte_in_4  (port_state_in_1_1_4    ), //i
    .port_byte_in_5  (port_state_in_1_1_5    ), //i
    .port_byte_in_6  (port_state_in_1_1_6    ), //i
    .port_byte_in_7  (port_state_in_1_1_7    ), //i
    .port_byte_out_0 (mul2_69_port_byte_out_0), //o
    .port_byte_out_1 (mul2_69_port_byte_out_1), //o
    .port_byte_out_2 (mul2_69_port_byte_out_2), //o
    .port_byte_out_3 (mul2_69_port_byte_out_3), //o
    .port_byte_out_4 (mul2_69_port_byte_out_4), //o
    .port_byte_out_5 (mul2_69_port_byte_out_5), //o
    .port_byte_out_6 (mul2_69_port_byte_out_6), //o
    .port_byte_out_7 (mul2_69_port_byte_out_7)  //o
  );
  Mul3 mul3_69 (
    .port_byte_in_0  (port_state_in_2_1_0    ), //i
    .port_byte_in_1  (port_state_in_2_1_1    ), //i
    .port_byte_in_2  (port_state_in_2_1_2    ), //i
    .port_byte_in_3  (port_state_in_2_1_3    ), //i
    .port_byte_in_4  (port_state_in_2_1_4    ), //i
    .port_byte_in_5  (port_state_in_2_1_5    ), //i
    .port_byte_in_6  (port_state_in_2_1_6    ), //i
    .port_byte_in_7  (port_state_in_2_1_7    ), //i
    .port_byte_out_0 (mul3_69_port_byte_out_0), //o
    .port_byte_out_1 (mul3_69_port_byte_out_1), //o
    .port_byte_out_2 (mul3_69_port_byte_out_2), //o
    .port_byte_out_3 (mul3_69_port_byte_out_3), //o
    .port_byte_out_4 (mul3_69_port_byte_out_4), //o
    .port_byte_out_5 (mul3_69_port_byte_out_5), //o
    .port_byte_out_6 (mul3_69_port_byte_out_6), //o
    .port_byte_out_7 (mul3_69_port_byte_out_7)  //o
  );
  Mul2 mul2_70 (
    .port_byte_in_0  (port_state_in_2_1_0    ), //i
    .port_byte_in_1  (port_state_in_2_1_1    ), //i
    .port_byte_in_2  (port_state_in_2_1_2    ), //i
    .port_byte_in_3  (port_state_in_2_1_3    ), //i
    .port_byte_in_4  (port_state_in_2_1_4    ), //i
    .port_byte_in_5  (port_state_in_2_1_5    ), //i
    .port_byte_in_6  (port_state_in_2_1_6    ), //i
    .port_byte_in_7  (port_state_in_2_1_7    ), //i
    .port_byte_out_0 (mul2_70_port_byte_out_0), //o
    .port_byte_out_1 (mul2_70_port_byte_out_1), //o
    .port_byte_out_2 (mul2_70_port_byte_out_2), //o
    .port_byte_out_3 (mul2_70_port_byte_out_3), //o
    .port_byte_out_4 (mul2_70_port_byte_out_4), //o
    .port_byte_out_5 (mul2_70_port_byte_out_5), //o
    .port_byte_out_6 (mul2_70_port_byte_out_6), //o
    .port_byte_out_7 (mul2_70_port_byte_out_7)  //o
  );
  Mul3 mul3_70 (
    .port_byte_in_0  (port_state_in_3_1_0    ), //i
    .port_byte_in_1  (port_state_in_3_1_1    ), //i
    .port_byte_in_2  (port_state_in_3_1_2    ), //i
    .port_byte_in_3  (port_state_in_3_1_3    ), //i
    .port_byte_in_4  (port_state_in_3_1_4    ), //i
    .port_byte_in_5  (port_state_in_3_1_5    ), //i
    .port_byte_in_6  (port_state_in_3_1_6    ), //i
    .port_byte_in_7  (port_state_in_3_1_7    ), //i
    .port_byte_out_0 (mul3_70_port_byte_out_0), //o
    .port_byte_out_1 (mul3_70_port_byte_out_1), //o
    .port_byte_out_2 (mul3_70_port_byte_out_2), //o
    .port_byte_out_3 (mul3_70_port_byte_out_3), //o
    .port_byte_out_4 (mul3_70_port_byte_out_4), //o
    .port_byte_out_5 (mul3_70_port_byte_out_5), //o
    .port_byte_out_6 (mul3_70_port_byte_out_6), //o
    .port_byte_out_7 (mul3_70_port_byte_out_7)  //o
  );
  Mul2 mul2_71 (
    .port_byte_in_0  (port_state_in_3_1_0    ), //i
    .port_byte_in_1  (port_state_in_3_1_1    ), //i
    .port_byte_in_2  (port_state_in_3_1_2    ), //i
    .port_byte_in_3  (port_state_in_3_1_3    ), //i
    .port_byte_in_4  (port_state_in_3_1_4    ), //i
    .port_byte_in_5  (port_state_in_3_1_5    ), //i
    .port_byte_in_6  (port_state_in_3_1_6    ), //i
    .port_byte_in_7  (port_state_in_3_1_7    ), //i
    .port_byte_out_0 (mul2_71_port_byte_out_0), //o
    .port_byte_out_1 (mul2_71_port_byte_out_1), //o
    .port_byte_out_2 (mul2_71_port_byte_out_2), //o
    .port_byte_out_3 (mul2_71_port_byte_out_3), //o
    .port_byte_out_4 (mul2_71_port_byte_out_4), //o
    .port_byte_out_5 (mul2_71_port_byte_out_5), //o
    .port_byte_out_6 (mul2_71_port_byte_out_6), //o
    .port_byte_out_7 (mul2_71_port_byte_out_7)  //o
  );
  Mul3 mul3_71 (
    .port_byte_in_0  (port_state_in_0_1_0    ), //i
    .port_byte_in_1  (port_state_in_0_1_1    ), //i
    .port_byte_in_2  (port_state_in_0_1_2    ), //i
    .port_byte_in_3  (port_state_in_0_1_3    ), //i
    .port_byte_in_4  (port_state_in_0_1_4    ), //i
    .port_byte_in_5  (port_state_in_0_1_5    ), //i
    .port_byte_in_6  (port_state_in_0_1_6    ), //i
    .port_byte_in_7  (port_state_in_0_1_7    ), //i
    .port_byte_out_0 (mul3_71_port_byte_out_0), //o
    .port_byte_out_1 (mul3_71_port_byte_out_1), //o
    .port_byte_out_2 (mul3_71_port_byte_out_2), //o
    .port_byte_out_3 (mul3_71_port_byte_out_3), //o
    .port_byte_out_4 (mul3_71_port_byte_out_4), //o
    .port_byte_out_5 (mul3_71_port_byte_out_5), //o
    .port_byte_out_6 (mul3_71_port_byte_out_6), //o
    .port_byte_out_7 (mul3_71_port_byte_out_7)  //o
  );
  Mul2 mul2_72 (
    .port_byte_in_0  (port_state_in_0_2_0    ), //i
    .port_byte_in_1  (port_state_in_0_2_1    ), //i
    .port_byte_in_2  (port_state_in_0_2_2    ), //i
    .port_byte_in_3  (port_state_in_0_2_3    ), //i
    .port_byte_in_4  (port_state_in_0_2_4    ), //i
    .port_byte_in_5  (port_state_in_0_2_5    ), //i
    .port_byte_in_6  (port_state_in_0_2_6    ), //i
    .port_byte_in_7  (port_state_in_0_2_7    ), //i
    .port_byte_out_0 (mul2_72_port_byte_out_0), //o
    .port_byte_out_1 (mul2_72_port_byte_out_1), //o
    .port_byte_out_2 (mul2_72_port_byte_out_2), //o
    .port_byte_out_3 (mul2_72_port_byte_out_3), //o
    .port_byte_out_4 (mul2_72_port_byte_out_4), //o
    .port_byte_out_5 (mul2_72_port_byte_out_5), //o
    .port_byte_out_6 (mul2_72_port_byte_out_6), //o
    .port_byte_out_7 (mul2_72_port_byte_out_7)  //o
  );
  Mul3 mul3_72 (
    .port_byte_in_0  (port_state_in_1_2_0    ), //i
    .port_byte_in_1  (port_state_in_1_2_1    ), //i
    .port_byte_in_2  (port_state_in_1_2_2    ), //i
    .port_byte_in_3  (port_state_in_1_2_3    ), //i
    .port_byte_in_4  (port_state_in_1_2_4    ), //i
    .port_byte_in_5  (port_state_in_1_2_5    ), //i
    .port_byte_in_6  (port_state_in_1_2_6    ), //i
    .port_byte_in_7  (port_state_in_1_2_7    ), //i
    .port_byte_out_0 (mul3_72_port_byte_out_0), //o
    .port_byte_out_1 (mul3_72_port_byte_out_1), //o
    .port_byte_out_2 (mul3_72_port_byte_out_2), //o
    .port_byte_out_3 (mul3_72_port_byte_out_3), //o
    .port_byte_out_4 (mul3_72_port_byte_out_4), //o
    .port_byte_out_5 (mul3_72_port_byte_out_5), //o
    .port_byte_out_6 (mul3_72_port_byte_out_6), //o
    .port_byte_out_7 (mul3_72_port_byte_out_7)  //o
  );
  Mul2 mul2_73 (
    .port_byte_in_0  (port_state_in_1_2_0    ), //i
    .port_byte_in_1  (port_state_in_1_2_1    ), //i
    .port_byte_in_2  (port_state_in_1_2_2    ), //i
    .port_byte_in_3  (port_state_in_1_2_3    ), //i
    .port_byte_in_4  (port_state_in_1_2_4    ), //i
    .port_byte_in_5  (port_state_in_1_2_5    ), //i
    .port_byte_in_6  (port_state_in_1_2_6    ), //i
    .port_byte_in_7  (port_state_in_1_2_7    ), //i
    .port_byte_out_0 (mul2_73_port_byte_out_0), //o
    .port_byte_out_1 (mul2_73_port_byte_out_1), //o
    .port_byte_out_2 (mul2_73_port_byte_out_2), //o
    .port_byte_out_3 (mul2_73_port_byte_out_3), //o
    .port_byte_out_4 (mul2_73_port_byte_out_4), //o
    .port_byte_out_5 (mul2_73_port_byte_out_5), //o
    .port_byte_out_6 (mul2_73_port_byte_out_6), //o
    .port_byte_out_7 (mul2_73_port_byte_out_7)  //o
  );
  Mul3 mul3_73 (
    .port_byte_in_0  (port_state_in_2_2_0    ), //i
    .port_byte_in_1  (port_state_in_2_2_1    ), //i
    .port_byte_in_2  (port_state_in_2_2_2    ), //i
    .port_byte_in_3  (port_state_in_2_2_3    ), //i
    .port_byte_in_4  (port_state_in_2_2_4    ), //i
    .port_byte_in_5  (port_state_in_2_2_5    ), //i
    .port_byte_in_6  (port_state_in_2_2_6    ), //i
    .port_byte_in_7  (port_state_in_2_2_7    ), //i
    .port_byte_out_0 (mul3_73_port_byte_out_0), //o
    .port_byte_out_1 (mul3_73_port_byte_out_1), //o
    .port_byte_out_2 (mul3_73_port_byte_out_2), //o
    .port_byte_out_3 (mul3_73_port_byte_out_3), //o
    .port_byte_out_4 (mul3_73_port_byte_out_4), //o
    .port_byte_out_5 (mul3_73_port_byte_out_5), //o
    .port_byte_out_6 (mul3_73_port_byte_out_6), //o
    .port_byte_out_7 (mul3_73_port_byte_out_7)  //o
  );
  Mul2 mul2_74 (
    .port_byte_in_0  (port_state_in_2_2_0    ), //i
    .port_byte_in_1  (port_state_in_2_2_1    ), //i
    .port_byte_in_2  (port_state_in_2_2_2    ), //i
    .port_byte_in_3  (port_state_in_2_2_3    ), //i
    .port_byte_in_4  (port_state_in_2_2_4    ), //i
    .port_byte_in_5  (port_state_in_2_2_5    ), //i
    .port_byte_in_6  (port_state_in_2_2_6    ), //i
    .port_byte_in_7  (port_state_in_2_2_7    ), //i
    .port_byte_out_0 (mul2_74_port_byte_out_0), //o
    .port_byte_out_1 (mul2_74_port_byte_out_1), //o
    .port_byte_out_2 (mul2_74_port_byte_out_2), //o
    .port_byte_out_3 (mul2_74_port_byte_out_3), //o
    .port_byte_out_4 (mul2_74_port_byte_out_4), //o
    .port_byte_out_5 (mul2_74_port_byte_out_5), //o
    .port_byte_out_6 (mul2_74_port_byte_out_6), //o
    .port_byte_out_7 (mul2_74_port_byte_out_7)  //o
  );
  Mul3 mul3_74 (
    .port_byte_in_0  (port_state_in_3_2_0    ), //i
    .port_byte_in_1  (port_state_in_3_2_1    ), //i
    .port_byte_in_2  (port_state_in_3_2_2    ), //i
    .port_byte_in_3  (port_state_in_3_2_3    ), //i
    .port_byte_in_4  (port_state_in_3_2_4    ), //i
    .port_byte_in_5  (port_state_in_3_2_5    ), //i
    .port_byte_in_6  (port_state_in_3_2_6    ), //i
    .port_byte_in_7  (port_state_in_3_2_7    ), //i
    .port_byte_out_0 (mul3_74_port_byte_out_0), //o
    .port_byte_out_1 (mul3_74_port_byte_out_1), //o
    .port_byte_out_2 (mul3_74_port_byte_out_2), //o
    .port_byte_out_3 (mul3_74_port_byte_out_3), //o
    .port_byte_out_4 (mul3_74_port_byte_out_4), //o
    .port_byte_out_5 (mul3_74_port_byte_out_5), //o
    .port_byte_out_6 (mul3_74_port_byte_out_6), //o
    .port_byte_out_7 (mul3_74_port_byte_out_7)  //o
  );
  Mul2 mul2_75 (
    .port_byte_in_0  (port_state_in_3_2_0    ), //i
    .port_byte_in_1  (port_state_in_3_2_1    ), //i
    .port_byte_in_2  (port_state_in_3_2_2    ), //i
    .port_byte_in_3  (port_state_in_3_2_3    ), //i
    .port_byte_in_4  (port_state_in_3_2_4    ), //i
    .port_byte_in_5  (port_state_in_3_2_5    ), //i
    .port_byte_in_6  (port_state_in_3_2_6    ), //i
    .port_byte_in_7  (port_state_in_3_2_7    ), //i
    .port_byte_out_0 (mul2_75_port_byte_out_0), //o
    .port_byte_out_1 (mul2_75_port_byte_out_1), //o
    .port_byte_out_2 (mul2_75_port_byte_out_2), //o
    .port_byte_out_3 (mul2_75_port_byte_out_3), //o
    .port_byte_out_4 (mul2_75_port_byte_out_4), //o
    .port_byte_out_5 (mul2_75_port_byte_out_5), //o
    .port_byte_out_6 (mul2_75_port_byte_out_6), //o
    .port_byte_out_7 (mul2_75_port_byte_out_7)  //o
  );
  Mul3 mul3_75 (
    .port_byte_in_0  (port_state_in_0_2_0    ), //i
    .port_byte_in_1  (port_state_in_0_2_1    ), //i
    .port_byte_in_2  (port_state_in_0_2_2    ), //i
    .port_byte_in_3  (port_state_in_0_2_3    ), //i
    .port_byte_in_4  (port_state_in_0_2_4    ), //i
    .port_byte_in_5  (port_state_in_0_2_5    ), //i
    .port_byte_in_6  (port_state_in_0_2_6    ), //i
    .port_byte_in_7  (port_state_in_0_2_7    ), //i
    .port_byte_out_0 (mul3_75_port_byte_out_0), //o
    .port_byte_out_1 (mul3_75_port_byte_out_1), //o
    .port_byte_out_2 (mul3_75_port_byte_out_2), //o
    .port_byte_out_3 (mul3_75_port_byte_out_3), //o
    .port_byte_out_4 (mul3_75_port_byte_out_4), //o
    .port_byte_out_5 (mul3_75_port_byte_out_5), //o
    .port_byte_out_6 (mul3_75_port_byte_out_6), //o
    .port_byte_out_7 (mul3_75_port_byte_out_7)  //o
  );
  Mul2 mul2_76 (
    .port_byte_in_0  (port_state_in_0_3_0    ), //i
    .port_byte_in_1  (port_state_in_0_3_1    ), //i
    .port_byte_in_2  (port_state_in_0_3_2    ), //i
    .port_byte_in_3  (port_state_in_0_3_3    ), //i
    .port_byte_in_4  (port_state_in_0_3_4    ), //i
    .port_byte_in_5  (port_state_in_0_3_5    ), //i
    .port_byte_in_6  (port_state_in_0_3_6    ), //i
    .port_byte_in_7  (port_state_in_0_3_7    ), //i
    .port_byte_out_0 (mul2_76_port_byte_out_0), //o
    .port_byte_out_1 (mul2_76_port_byte_out_1), //o
    .port_byte_out_2 (mul2_76_port_byte_out_2), //o
    .port_byte_out_3 (mul2_76_port_byte_out_3), //o
    .port_byte_out_4 (mul2_76_port_byte_out_4), //o
    .port_byte_out_5 (mul2_76_port_byte_out_5), //o
    .port_byte_out_6 (mul2_76_port_byte_out_6), //o
    .port_byte_out_7 (mul2_76_port_byte_out_7)  //o
  );
  Mul3 mul3_76 (
    .port_byte_in_0  (port_state_in_1_3_0    ), //i
    .port_byte_in_1  (port_state_in_1_3_1    ), //i
    .port_byte_in_2  (port_state_in_1_3_2    ), //i
    .port_byte_in_3  (port_state_in_1_3_3    ), //i
    .port_byte_in_4  (port_state_in_1_3_4    ), //i
    .port_byte_in_5  (port_state_in_1_3_5    ), //i
    .port_byte_in_6  (port_state_in_1_3_6    ), //i
    .port_byte_in_7  (port_state_in_1_3_7    ), //i
    .port_byte_out_0 (mul3_76_port_byte_out_0), //o
    .port_byte_out_1 (mul3_76_port_byte_out_1), //o
    .port_byte_out_2 (mul3_76_port_byte_out_2), //o
    .port_byte_out_3 (mul3_76_port_byte_out_3), //o
    .port_byte_out_4 (mul3_76_port_byte_out_4), //o
    .port_byte_out_5 (mul3_76_port_byte_out_5), //o
    .port_byte_out_6 (mul3_76_port_byte_out_6), //o
    .port_byte_out_7 (mul3_76_port_byte_out_7)  //o
  );
  Mul2 mul2_77 (
    .port_byte_in_0  (port_state_in_1_3_0    ), //i
    .port_byte_in_1  (port_state_in_1_3_1    ), //i
    .port_byte_in_2  (port_state_in_1_3_2    ), //i
    .port_byte_in_3  (port_state_in_1_3_3    ), //i
    .port_byte_in_4  (port_state_in_1_3_4    ), //i
    .port_byte_in_5  (port_state_in_1_3_5    ), //i
    .port_byte_in_6  (port_state_in_1_3_6    ), //i
    .port_byte_in_7  (port_state_in_1_3_7    ), //i
    .port_byte_out_0 (mul2_77_port_byte_out_0), //o
    .port_byte_out_1 (mul2_77_port_byte_out_1), //o
    .port_byte_out_2 (mul2_77_port_byte_out_2), //o
    .port_byte_out_3 (mul2_77_port_byte_out_3), //o
    .port_byte_out_4 (mul2_77_port_byte_out_4), //o
    .port_byte_out_5 (mul2_77_port_byte_out_5), //o
    .port_byte_out_6 (mul2_77_port_byte_out_6), //o
    .port_byte_out_7 (mul2_77_port_byte_out_7)  //o
  );
  Mul3 mul3_77 (
    .port_byte_in_0  (port_state_in_2_3_0    ), //i
    .port_byte_in_1  (port_state_in_2_3_1    ), //i
    .port_byte_in_2  (port_state_in_2_3_2    ), //i
    .port_byte_in_3  (port_state_in_2_3_3    ), //i
    .port_byte_in_4  (port_state_in_2_3_4    ), //i
    .port_byte_in_5  (port_state_in_2_3_5    ), //i
    .port_byte_in_6  (port_state_in_2_3_6    ), //i
    .port_byte_in_7  (port_state_in_2_3_7    ), //i
    .port_byte_out_0 (mul3_77_port_byte_out_0), //o
    .port_byte_out_1 (mul3_77_port_byte_out_1), //o
    .port_byte_out_2 (mul3_77_port_byte_out_2), //o
    .port_byte_out_3 (mul3_77_port_byte_out_3), //o
    .port_byte_out_4 (mul3_77_port_byte_out_4), //o
    .port_byte_out_5 (mul3_77_port_byte_out_5), //o
    .port_byte_out_6 (mul3_77_port_byte_out_6), //o
    .port_byte_out_7 (mul3_77_port_byte_out_7)  //o
  );
  Mul2 mul2_78 (
    .port_byte_in_0  (port_state_in_2_3_0    ), //i
    .port_byte_in_1  (port_state_in_2_3_1    ), //i
    .port_byte_in_2  (port_state_in_2_3_2    ), //i
    .port_byte_in_3  (port_state_in_2_3_3    ), //i
    .port_byte_in_4  (port_state_in_2_3_4    ), //i
    .port_byte_in_5  (port_state_in_2_3_5    ), //i
    .port_byte_in_6  (port_state_in_2_3_6    ), //i
    .port_byte_in_7  (port_state_in_2_3_7    ), //i
    .port_byte_out_0 (mul2_78_port_byte_out_0), //o
    .port_byte_out_1 (mul2_78_port_byte_out_1), //o
    .port_byte_out_2 (mul2_78_port_byte_out_2), //o
    .port_byte_out_3 (mul2_78_port_byte_out_3), //o
    .port_byte_out_4 (mul2_78_port_byte_out_4), //o
    .port_byte_out_5 (mul2_78_port_byte_out_5), //o
    .port_byte_out_6 (mul2_78_port_byte_out_6), //o
    .port_byte_out_7 (mul2_78_port_byte_out_7)  //o
  );
  Mul3 mul3_78 (
    .port_byte_in_0  (port_state_in_3_3_0    ), //i
    .port_byte_in_1  (port_state_in_3_3_1    ), //i
    .port_byte_in_2  (port_state_in_3_3_2    ), //i
    .port_byte_in_3  (port_state_in_3_3_3    ), //i
    .port_byte_in_4  (port_state_in_3_3_4    ), //i
    .port_byte_in_5  (port_state_in_3_3_5    ), //i
    .port_byte_in_6  (port_state_in_3_3_6    ), //i
    .port_byte_in_7  (port_state_in_3_3_7    ), //i
    .port_byte_out_0 (mul3_78_port_byte_out_0), //o
    .port_byte_out_1 (mul3_78_port_byte_out_1), //o
    .port_byte_out_2 (mul3_78_port_byte_out_2), //o
    .port_byte_out_3 (mul3_78_port_byte_out_3), //o
    .port_byte_out_4 (mul3_78_port_byte_out_4), //o
    .port_byte_out_5 (mul3_78_port_byte_out_5), //o
    .port_byte_out_6 (mul3_78_port_byte_out_6), //o
    .port_byte_out_7 (mul3_78_port_byte_out_7)  //o
  );
  Mul2 mul2_79 (
    .port_byte_in_0  (port_state_in_3_3_0    ), //i
    .port_byte_in_1  (port_state_in_3_3_1    ), //i
    .port_byte_in_2  (port_state_in_3_3_2    ), //i
    .port_byte_in_3  (port_state_in_3_3_3    ), //i
    .port_byte_in_4  (port_state_in_3_3_4    ), //i
    .port_byte_in_5  (port_state_in_3_3_5    ), //i
    .port_byte_in_6  (port_state_in_3_3_6    ), //i
    .port_byte_in_7  (port_state_in_3_3_7    ), //i
    .port_byte_out_0 (mul2_79_port_byte_out_0), //o
    .port_byte_out_1 (mul2_79_port_byte_out_1), //o
    .port_byte_out_2 (mul2_79_port_byte_out_2), //o
    .port_byte_out_3 (mul2_79_port_byte_out_3), //o
    .port_byte_out_4 (mul2_79_port_byte_out_4), //o
    .port_byte_out_5 (mul2_79_port_byte_out_5), //o
    .port_byte_out_6 (mul2_79_port_byte_out_6), //o
    .port_byte_out_7 (mul2_79_port_byte_out_7)  //o
  );
  Mul3 mul3_79 (
    .port_byte_in_0  (port_state_in_0_3_0    ), //i
    .port_byte_in_1  (port_state_in_0_3_1    ), //i
    .port_byte_in_2  (port_state_in_0_3_2    ), //i
    .port_byte_in_3  (port_state_in_0_3_3    ), //i
    .port_byte_in_4  (port_state_in_0_3_4    ), //i
    .port_byte_in_5  (port_state_in_0_3_5    ), //i
    .port_byte_in_6  (port_state_in_0_3_6    ), //i
    .port_byte_in_7  (port_state_in_0_3_7    ), //i
    .port_byte_out_0 (mul3_79_port_byte_out_0), //o
    .port_byte_out_1 (mul3_79_port_byte_out_1), //o
    .port_byte_out_2 (mul3_79_port_byte_out_2), //o
    .port_byte_out_3 (mul3_79_port_byte_out_3), //o
    .port_byte_out_4 (mul3_79_port_byte_out_4), //o
    .port_byte_out_5 (mul3_79_port_byte_out_5), //o
    .port_byte_out_6 (mul3_79_port_byte_out_6), //o
    .port_byte_out_7 (mul3_79_port_byte_out_7)  //o
  );
  Mul2 mul2_80 (
    .port_byte_in_0  (port_state_in_4_0_0    ), //i
    .port_byte_in_1  (port_state_in_4_0_1    ), //i
    .port_byte_in_2  (port_state_in_4_0_2    ), //i
    .port_byte_in_3  (port_state_in_4_0_3    ), //i
    .port_byte_in_4  (port_state_in_4_0_4    ), //i
    .port_byte_in_5  (port_state_in_4_0_5    ), //i
    .port_byte_in_6  (port_state_in_4_0_6    ), //i
    .port_byte_in_7  (port_state_in_4_0_7    ), //i
    .port_byte_out_0 (mul2_80_port_byte_out_0), //o
    .port_byte_out_1 (mul2_80_port_byte_out_1), //o
    .port_byte_out_2 (mul2_80_port_byte_out_2), //o
    .port_byte_out_3 (mul2_80_port_byte_out_3), //o
    .port_byte_out_4 (mul2_80_port_byte_out_4), //o
    .port_byte_out_5 (mul2_80_port_byte_out_5), //o
    .port_byte_out_6 (mul2_80_port_byte_out_6), //o
    .port_byte_out_7 (mul2_80_port_byte_out_7)  //o
  );
  Mul3 mul3_80 (
    .port_byte_in_0  (port_state_in_5_0_0    ), //i
    .port_byte_in_1  (port_state_in_5_0_1    ), //i
    .port_byte_in_2  (port_state_in_5_0_2    ), //i
    .port_byte_in_3  (port_state_in_5_0_3    ), //i
    .port_byte_in_4  (port_state_in_5_0_4    ), //i
    .port_byte_in_5  (port_state_in_5_0_5    ), //i
    .port_byte_in_6  (port_state_in_5_0_6    ), //i
    .port_byte_in_7  (port_state_in_5_0_7    ), //i
    .port_byte_out_0 (mul3_80_port_byte_out_0), //o
    .port_byte_out_1 (mul3_80_port_byte_out_1), //o
    .port_byte_out_2 (mul3_80_port_byte_out_2), //o
    .port_byte_out_3 (mul3_80_port_byte_out_3), //o
    .port_byte_out_4 (mul3_80_port_byte_out_4), //o
    .port_byte_out_5 (mul3_80_port_byte_out_5), //o
    .port_byte_out_6 (mul3_80_port_byte_out_6), //o
    .port_byte_out_7 (mul3_80_port_byte_out_7)  //o
  );
  Mul2 mul2_81 (
    .port_byte_in_0  (port_state_in_5_0_0    ), //i
    .port_byte_in_1  (port_state_in_5_0_1    ), //i
    .port_byte_in_2  (port_state_in_5_0_2    ), //i
    .port_byte_in_3  (port_state_in_5_0_3    ), //i
    .port_byte_in_4  (port_state_in_5_0_4    ), //i
    .port_byte_in_5  (port_state_in_5_0_5    ), //i
    .port_byte_in_6  (port_state_in_5_0_6    ), //i
    .port_byte_in_7  (port_state_in_5_0_7    ), //i
    .port_byte_out_0 (mul2_81_port_byte_out_0), //o
    .port_byte_out_1 (mul2_81_port_byte_out_1), //o
    .port_byte_out_2 (mul2_81_port_byte_out_2), //o
    .port_byte_out_3 (mul2_81_port_byte_out_3), //o
    .port_byte_out_4 (mul2_81_port_byte_out_4), //o
    .port_byte_out_5 (mul2_81_port_byte_out_5), //o
    .port_byte_out_6 (mul2_81_port_byte_out_6), //o
    .port_byte_out_7 (mul2_81_port_byte_out_7)  //o
  );
  Mul3 mul3_81 (
    .port_byte_in_0  (port_state_in_6_0_0    ), //i
    .port_byte_in_1  (port_state_in_6_0_1    ), //i
    .port_byte_in_2  (port_state_in_6_0_2    ), //i
    .port_byte_in_3  (port_state_in_6_0_3    ), //i
    .port_byte_in_4  (port_state_in_6_0_4    ), //i
    .port_byte_in_5  (port_state_in_6_0_5    ), //i
    .port_byte_in_6  (port_state_in_6_0_6    ), //i
    .port_byte_in_7  (port_state_in_6_0_7    ), //i
    .port_byte_out_0 (mul3_81_port_byte_out_0), //o
    .port_byte_out_1 (mul3_81_port_byte_out_1), //o
    .port_byte_out_2 (mul3_81_port_byte_out_2), //o
    .port_byte_out_3 (mul3_81_port_byte_out_3), //o
    .port_byte_out_4 (mul3_81_port_byte_out_4), //o
    .port_byte_out_5 (mul3_81_port_byte_out_5), //o
    .port_byte_out_6 (mul3_81_port_byte_out_6), //o
    .port_byte_out_7 (mul3_81_port_byte_out_7)  //o
  );
  Mul2 mul2_82 (
    .port_byte_in_0  (port_state_in_6_0_0    ), //i
    .port_byte_in_1  (port_state_in_6_0_1    ), //i
    .port_byte_in_2  (port_state_in_6_0_2    ), //i
    .port_byte_in_3  (port_state_in_6_0_3    ), //i
    .port_byte_in_4  (port_state_in_6_0_4    ), //i
    .port_byte_in_5  (port_state_in_6_0_5    ), //i
    .port_byte_in_6  (port_state_in_6_0_6    ), //i
    .port_byte_in_7  (port_state_in_6_0_7    ), //i
    .port_byte_out_0 (mul2_82_port_byte_out_0), //o
    .port_byte_out_1 (mul2_82_port_byte_out_1), //o
    .port_byte_out_2 (mul2_82_port_byte_out_2), //o
    .port_byte_out_3 (mul2_82_port_byte_out_3), //o
    .port_byte_out_4 (mul2_82_port_byte_out_4), //o
    .port_byte_out_5 (mul2_82_port_byte_out_5), //o
    .port_byte_out_6 (mul2_82_port_byte_out_6), //o
    .port_byte_out_7 (mul2_82_port_byte_out_7)  //o
  );
  Mul3 mul3_82 (
    .port_byte_in_0  (port_state_in_7_0_0    ), //i
    .port_byte_in_1  (port_state_in_7_0_1    ), //i
    .port_byte_in_2  (port_state_in_7_0_2    ), //i
    .port_byte_in_3  (port_state_in_7_0_3    ), //i
    .port_byte_in_4  (port_state_in_7_0_4    ), //i
    .port_byte_in_5  (port_state_in_7_0_5    ), //i
    .port_byte_in_6  (port_state_in_7_0_6    ), //i
    .port_byte_in_7  (port_state_in_7_0_7    ), //i
    .port_byte_out_0 (mul3_82_port_byte_out_0), //o
    .port_byte_out_1 (mul3_82_port_byte_out_1), //o
    .port_byte_out_2 (mul3_82_port_byte_out_2), //o
    .port_byte_out_3 (mul3_82_port_byte_out_3), //o
    .port_byte_out_4 (mul3_82_port_byte_out_4), //o
    .port_byte_out_5 (mul3_82_port_byte_out_5), //o
    .port_byte_out_6 (mul3_82_port_byte_out_6), //o
    .port_byte_out_7 (mul3_82_port_byte_out_7)  //o
  );
  Mul2 mul2_83 (
    .port_byte_in_0  (port_state_in_7_0_0    ), //i
    .port_byte_in_1  (port_state_in_7_0_1    ), //i
    .port_byte_in_2  (port_state_in_7_0_2    ), //i
    .port_byte_in_3  (port_state_in_7_0_3    ), //i
    .port_byte_in_4  (port_state_in_7_0_4    ), //i
    .port_byte_in_5  (port_state_in_7_0_5    ), //i
    .port_byte_in_6  (port_state_in_7_0_6    ), //i
    .port_byte_in_7  (port_state_in_7_0_7    ), //i
    .port_byte_out_0 (mul2_83_port_byte_out_0), //o
    .port_byte_out_1 (mul2_83_port_byte_out_1), //o
    .port_byte_out_2 (mul2_83_port_byte_out_2), //o
    .port_byte_out_3 (mul2_83_port_byte_out_3), //o
    .port_byte_out_4 (mul2_83_port_byte_out_4), //o
    .port_byte_out_5 (mul2_83_port_byte_out_5), //o
    .port_byte_out_6 (mul2_83_port_byte_out_6), //o
    .port_byte_out_7 (mul2_83_port_byte_out_7)  //o
  );
  Mul3 mul3_83 (
    .port_byte_in_0  (port_state_in_4_0_0    ), //i
    .port_byte_in_1  (port_state_in_4_0_1    ), //i
    .port_byte_in_2  (port_state_in_4_0_2    ), //i
    .port_byte_in_3  (port_state_in_4_0_3    ), //i
    .port_byte_in_4  (port_state_in_4_0_4    ), //i
    .port_byte_in_5  (port_state_in_4_0_5    ), //i
    .port_byte_in_6  (port_state_in_4_0_6    ), //i
    .port_byte_in_7  (port_state_in_4_0_7    ), //i
    .port_byte_out_0 (mul3_83_port_byte_out_0), //o
    .port_byte_out_1 (mul3_83_port_byte_out_1), //o
    .port_byte_out_2 (mul3_83_port_byte_out_2), //o
    .port_byte_out_3 (mul3_83_port_byte_out_3), //o
    .port_byte_out_4 (mul3_83_port_byte_out_4), //o
    .port_byte_out_5 (mul3_83_port_byte_out_5), //o
    .port_byte_out_6 (mul3_83_port_byte_out_6), //o
    .port_byte_out_7 (mul3_83_port_byte_out_7)  //o
  );
  Mul2 mul2_84 (
    .port_byte_in_0  (port_state_in_4_1_0    ), //i
    .port_byte_in_1  (port_state_in_4_1_1    ), //i
    .port_byte_in_2  (port_state_in_4_1_2    ), //i
    .port_byte_in_3  (port_state_in_4_1_3    ), //i
    .port_byte_in_4  (port_state_in_4_1_4    ), //i
    .port_byte_in_5  (port_state_in_4_1_5    ), //i
    .port_byte_in_6  (port_state_in_4_1_6    ), //i
    .port_byte_in_7  (port_state_in_4_1_7    ), //i
    .port_byte_out_0 (mul2_84_port_byte_out_0), //o
    .port_byte_out_1 (mul2_84_port_byte_out_1), //o
    .port_byte_out_2 (mul2_84_port_byte_out_2), //o
    .port_byte_out_3 (mul2_84_port_byte_out_3), //o
    .port_byte_out_4 (mul2_84_port_byte_out_4), //o
    .port_byte_out_5 (mul2_84_port_byte_out_5), //o
    .port_byte_out_6 (mul2_84_port_byte_out_6), //o
    .port_byte_out_7 (mul2_84_port_byte_out_7)  //o
  );
  Mul3 mul3_84 (
    .port_byte_in_0  (port_state_in_5_1_0    ), //i
    .port_byte_in_1  (port_state_in_5_1_1    ), //i
    .port_byte_in_2  (port_state_in_5_1_2    ), //i
    .port_byte_in_3  (port_state_in_5_1_3    ), //i
    .port_byte_in_4  (port_state_in_5_1_4    ), //i
    .port_byte_in_5  (port_state_in_5_1_5    ), //i
    .port_byte_in_6  (port_state_in_5_1_6    ), //i
    .port_byte_in_7  (port_state_in_5_1_7    ), //i
    .port_byte_out_0 (mul3_84_port_byte_out_0), //o
    .port_byte_out_1 (mul3_84_port_byte_out_1), //o
    .port_byte_out_2 (mul3_84_port_byte_out_2), //o
    .port_byte_out_3 (mul3_84_port_byte_out_3), //o
    .port_byte_out_4 (mul3_84_port_byte_out_4), //o
    .port_byte_out_5 (mul3_84_port_byte_out_5), //o
    .port_byte_out_6 (mul3_84_port_byte_out_6), //o
    .port_byte_out_7 (mul3_84_port_byte_out_7)  //o
  );
  Mul2 mul2_85 (
    .port_byte_in_0  (port_state_in_5_1_0    ), //i
    .port_byte_in_1  (port_state_in_5_1_1    ), //i
    .port_byte_in_2  (port_state_in_5_1_2    ), //i
    .port_byte_in_3  (port_state_in_5_1_3    ), //i
    .port_byte_in_4  (port_state_in_5_1_4    ), //i
    .port_byte_in_5  (port_state_in_5_1_5    ), //i
    .port_byte_in_6  (port_state_in_5_1_6    ), //i
    .port_byte_in_7  (port_state_in_5_1_7    ), //i
    .port_byte_out_0 (mul2_85_port_byte_out_0), //o
    .port_byte_out_1 (mul2_85_port_byte_out_1), //o
    .port_byte_out_2 (mul2_85_port_byte_out_2), //o
    .port_byte_out_3 (mul2_85_port_byte_out_3), //o
    .port_byte_out_4 (mul2_85_port_byte_out_4), //o
    .port_byte_out_5 (mul2_85_port_byte_out_5), //o
    .port_byte_out_6 (mul2_85_port_byte_out_6), //o
    .port_byte_out_7 (mul2_85_port_byte_out_7)  //o
  );
  Mul3 mul3_85 (
    .port_byte_in_0  (port_state_in_6_1_0    ), //i
    .port_byte_in_1  (port_state_in_6_1_1    ), //i
    .port_byte_in_2  (port_state_in_6_1_2    ), //i
    .port_byte_in_3  (port_state_in_6_1_3    ), //i
    .port_byte_in_4  (port_state_in_6_1_4    ), //i
    .port_byte_in_5  (port_state_in_6_1_5    ), //i
    .port_byte_in_6  (port_state_in_6_1_6    ), //i
    .port_byte_in_7  (port_state_in_6_1_7    ), //i
    .port_byte_out_0 (mul3_85_port_byte_out_0), //o
    .port_byte_out_1 (mul3_85_port_byte_out_1), //o
    .port_byte_out_2 (mul3_85_port_byte_out_2), //o
    .port_byte_out_3 (mul3_85_port_byte_out_3), //o
    .port_byte_out_4 (mul3_85_port_byte_out_4), //o
    .port_byte_out_5 (mul3_85_port_byte_out_5), //o
    .port_byte_out_6 (mul3_85_port_byte_out_6), //o
    .port_byte_out_7 (mul3_85_port_byte_out_7)  //o
  );
  Mul2 mul2_86 (
    .port_byte_in_0  (port_state_in_6_1_0    ), //i
    .port_byte_in_1  (port_state_in_6_1_1    ), //i
    .port_byte_in_2  (port_state_in_6_1_2    ), //i
    .port_byte_in_3  (port_state_in_6_1_3    ), //i
    .port_byte_in_4  (port_state_in_6_1_4    ), //i
    .port_byte_in_5  (port_state_in_6_1_5    ), //i
    .port_byte_in_6  (port_state_in_6_1_6    ), //i
    .port_byte_in_7  (port_state_in_6_1_7    ), //i
    .port_byte_out_0 (mul2_86_port_byte_out_0), //o
    .port_byte_out_1 (mul2_86_port_byte_out_1), //o
    .port_byte_out_2 (mul2_86_port_byte_out_2), //o
    .port_byte_out_3 (mul2_86_port_byte_out_3), //o
    .port_byte_out_4 (mul2_86_port_byte_out_4), //o
    .port_byte_out_5 (mul2_86_port_byte_out_5), //o
    .port_byte_out_6 (mul2_86_port_byte_out_6), //o
    .port_byte_out_7 (mul2_86_port_byte_out_7)  //o
  );
  Mul3 mul3_86 (
    .port_byte_in_0  (port_state_in_7_1_0    ), //i
    .port_byte_in_1  (port_state_in_7_1_1    ), //i
    .port_byte_in_2  (port_state_in_7_1_2    ), //i
    .port_byte_in_3  (port_state_in_7_1_3    ), //i
    .port_byte_in_4  (port_state_in_7_1_4    ), //i
    .port_byte_in_5  (port_state_in_7_1_5    ), //i
    .port_byte_in_6  (port_state_in_7_1_6    ), //i
    .port_byte_in_7  (port_state_in_7_1_7    ), //i
    .port_byte_out_0 (mul3_86_port_byte_out_0), //o
    .port_byte_out_1 (mul3_86_port_byte_out_1), //o
    .port_byte_out_2 (mul3_86_port_byte_out_2), //o
    .port_byte_out_3 (mul3_86_port_byte_out_3), //o
    .port_byte_out_4 (mul3_86_port_byte_out_4), //o
    .port_byte_out_5 (mul3_86_port_byte_out_5), //o
    .port_byte_out_6 (mul3_86_port_byte_out_6), //o
    .port_byte_out_7 (mul3_86_port_byte_out_7)  //o
  );
  Mul2 mul2_87 (
    .port_byte_in_0  (port_state_in_7_1_0    ), //i
    .port_byte_in_1  (port_state_in_7_1_1    ), //i
    .port_byte_in_2  (port_state_in_7_1_2    ), //i
    .port_byte_in_3  (port_state_in_7_1_3    ), //i
    .port_byte_in_4  (port_state_in_7_1_4    ), //i
    .port_byte_in_5  (port_state_in_7_1_5    ), //i
    .port_byte_in_6  (port_state_in_7_1_6    ), //i
    .port_byte_in_7  (port_state_in_7_1_7    ), //i
    .port_byte_out_0 (mul2_87_port_byte_out_0), //o
    .port_byte_out_1 (mul2_87_port_byte_out_1), //o
    .port_byte_out_2 (mul2_87_port_byte_out_2), //o
    .port_byte_out_3 (mul2_87_port_byte_out_3), //o
    .port_byte_out_4 (mul2_87_port_byte_out_4), //o
    .port_byte_out_5 (mul2_87_port_byte_out_5), //o
    .port_byte_out_6 (mul2_87_port_byte_out_6), //o
    .port_byte_out_7 (mul2_87_port_byte_out_7)  //o
  );
  Mul3 mul3_87 (
    .port_byte_in_0  (port_state_in_4_1_0    ), //i
    .port_byte_in_1  (port_state_in_4_1_1    ), //i
    .port_byte_in_2  (port_state_in_4_1_2    ), //i
    .port_byte_in_3  (port_state_in_4_1_3    ), //i
    .port_byte_in_4  (port_state_in_4_1_4    ), //i
    .port_byte_in_5  (port_state_in_4_1_5    ), //i
    .port_byte_in_6  (port_state_in_4_1_6    ), //i
    .port_byte_in_7  (port_state_in_4_1_7    ), //i
    .port_byte_out_0 (mul3_87_port_byte_out_0), //o
    .port_byte_out_1 (mul3_87_port_byte_out_1), //o
    .port_byte_out_2 (mul3_87_port_byte_out_2), //o
    .port_byte_out_3 (mul3_87_port_byte_out_3), //o
    .port_byte_out_4 (mul3_87_port_byte_out_4), //o
    .port_byte_out_5 (mul3_87_port_byte_out_5), //o
    .port_byte_out_6 (mul3_87_port_byte_out_6), //o
    .port_byte_out_7 (mul3_87_port_byte_out_7)  //o
  );
  Mul2 mul2_88 (
    .port_byte_in_0  (port_state_in_4_2_0    ), //i
    .port_byte_in_1  (port_state_in_4_2_1    ), //i
    .port_byte_in_2  (port_state_in_4_2_2    ), //i
    .port_byte_in_3  (port_state_in_4_2_3    ), //i
    .port_byte_in_4  (port_state_in_4_2_4    ), //i
    .port_byte_in_5  (port_state_in_4_2_5    ), //i
    .port_byte_in_6  (port_state_in_4_2_6    ), //i
    .port_byte_in_7  (port_state_in_4_2_7    ), //i
    .port_byte_out_0 (mul2_88_port_byte_out_0), //o
    .port_byte_out_1 (mul2_88_port_byte_out_1), //o
    .port_byte_out_2 (mul2_88_port_byte_out_2), //o
    .port_byte_out_3 (mul2_88_port_byte_out_3), //o
    .port_byte_out_4 (mul2_88_port_byte_out_4), //o
    .port_byte_out_5 (mul2_88_port_byte_out_5), //o
    .port_byte_out_6 (mul2_88_port_byte_out_6), //o
    .port_byte_out_7 (mul2_88_port_byte_out_7)  //o
  );
  Mul3 mul3_88 (
    .port_byte_in_0  (port_state_in_5_2_0    ), //i
    .port_byte_in_1  (port_state_in_5_2_1    ), //i
    .port_byte_in_2  (port_state_in_5_2_2    ), //i
    .port_byte_in_3  (port_state_in_5_2_3    ), //i
    .port_byte_in_4  (port_state_in_5_2_4    ), //i
    .port_byte_in_5  (port_state_in_5_2_5    ), //i
    .port_byte_in_6  (port_state_in_5_2_6    ), //i
    .port_byte_in_7  (port_state_in_5_2_7    ), //i
    .port_byte_out_0 (mul3_88_port_byte_out_0), //o
    .port_byte_out_1 (mul3_88_port_byte_out_1), //o
    .port_byte_out_2 (mul3_88_port_byte_out_2), //o
    .port_byte_out_3 (mul3_88_port_byte_out_3), //o
    .port_byte_out_4 (mul3_88_port_byte_out_4), //o
    .port_byte_out_5 (mul3_88_port_byte_out_5), //o
    .port_byte_out_6 (mul3_88_port_byte_out_6), //o
    .port_byte_out_7 (mul3_88_port_byte_out_7)  //o
  );
  Mul2 mul2_89 (
    .port_byte_in_0  (port_state_in_5_2_0    ), //i
    .port_byte_in_1  (port_state_in_5_2_1    ), //i
    .port_byte_in_2  (port_state_in_5_2_2    ), //i
    .port_byte_in_3  (port_state_in_5_2_3    ), //i
    .port_byte_in_4  (port_state_in_5_2_4    ), //i
    .port_byte_in_5  (port_state_in_5_2_5    ), //i
    .port_byte_in_6  (port_state_in_5_2_6    ), //i
    .port_byte_in_7  (port_state_in_5_2_7    ), //i
    .port_byte_out_0 (mul2_89_port_byte_out_0), //o
    .port_byte_out_1 (mul2_89_port_byte_out_1), //o
    .port_byte_out_2 (mul2_89_port_byte_out_2), //o
    .port_byte_out_3 (mul2_89_port_byte_out_3), //o
    .port_byte_out_4 (mul2_89_port_byte_out_4), //o
    .port_byte_out_5 (mul2_89_port_byte_out_5), //o
    .port_byte_out_6 (mul2_89_port_byte_out_6), //o
    .port_byte_out_7 (mul2_89_port_byte_out_7)  //o
  );
  Mul3 mul3_89 (
    .port_byte_in_0  (port_state_in_6_2_0    ), //i
    .port_byte_in_1  (port_state_in_6_2_1    ), //i
    .port_byte_in_2  (port_state_in_6_2_2    ), //i
    .port_byte_in_3  (port_state_in_6_2_3    ), //i
    .port_byte_in_4  (port_state_in_6_2_4    ), //i
    .port_byte_in_5  (port_state_in_6_2_5    ), //i
    .port_byte_in_6  (port_state_in_6_2_6    ), //i
    .port_byte_in_7  (port_state_in_6_2_7    ), //i
    .port_byte_out_0 (mul3_89_port_byte_out_0), //o
    .port_byte_out_1 (mul3_89_port_byte_out_1), //o
    .port_byte_out_2 (mul3_89_port_byte_out_2), //o
    .port_byte_out_3 (mul3_89_port_byte_out_3), //o
    .port_byte_out_4 (mul3_89_port_byte_out_4), //o
    .port_byte_out_5 (mul3_89_port_byte_out_5), //o
    .port_byte_out_6 (mul3_89_port_byte_out_6), //o
    .port_byte_out_7 (mul3_89_port_byte_out_7)  //o
  );
  Mul2 mul2_90 (
    .port_byte_in_0  (port_state_in_6_2_0    ), //i
    .port_byte_in_1  (port_state_in_6_2_1    ), //i
    .port_byte_in_2  (port_state_in_6_2_2    ), //i
    .port_byte_in_3  (port_state_in_6_2_3    ), //i
    .port_byte_in_4  (port_state_in_6_2_4    ), //i
    .port_byte_in_5  (port_state_in_6_2_5    ), //i
    .port_byte_in_6  (port_state_in_6_2_6    ), //i
    .port_byte_in_7  (port_state_in_6_2_7    ), //i
    .port_byte_out_0 (mul2_90_port_byte_out_0), //o
    .port_byte_out_1 (mul2_90_port_byte_out_1), //o
    .port_byte_out_2 (mul2_90_port_byte_out_2), //o
    .port_byte_out_3 (mul2_90_port_byte_out_3), //o
    .port_byte_out_4 (mul2_90_port_byte_out_4), //o
    .port_byte_out_5 (mul2_90_port_byte_out_5), //o
    .port_byte_out_6 (mul2_90_port_byte_out_6), //o
    .port_byte_out_7 (mul2_90_port_byte_out_7)  //o
  );
  Mul3 mul3_90 (
    .port_byte_in_0  (port_state_in_7_2_0    ), //i
    .port_byte_in_1  (port_state_in_7_2_1    ), //i
    .port_byte_in_2  (port_state_in_7_2_2    ), //i
    .port_byte_in_3  (port_state_in_7_2_3    ), //i
    .port_byte_in_4  (port_state_in_7_2_4    ), //i
    .port_byte_in_5  (port_state_in_7_2_5    ), //i
    .port_byte_in_6  (port_state_in_7_2_6    ), //i
    .port_byte_in_7  (port_state_in_7_2_7    ), //i
    .port_byte_out_0 (mul3_90_port_byte_out_0), //o
    .port_byte_out_1 (mul3_90_port_byte_out_1), //o
    .port_byte_out_2 (mul3_90_port_byte_out_2), //o
    .port_byte_out_3 (mul3_90_port_byte_out_3), //o
    .port_byte_out_4 (mul3_90_port_byte_out_4), //o
    .port_byte_out_5 (mul3_90_port_byte_out_5), //o
    .port_byte_out_6 (mul3_90_port_byte_out_6), //o
    .port_byte_out_7 (mul3_90_port_byte_out_7)  //o
  );
  Mul2 mul2_91 (
    .port_byte_in_0  (port_state_in_7_2_0    ), //i
    .port_byte_in_1  (port_state_in_7_2_1    ), //i
    .port_byte_in_2  (port_state_in_7_2_2    ), //i
    .port_byte_in_3  (port_state_in_7_2_3    ), //i
    .port_byte_in_4  (port_state_in_7_2_4    ), //i
    .port_byte_in_5  (port_state_in_7_2_5    ), //i
    .port_byte_in_6  (port_state_in_7_2_6    ), //i
    .port_byte_in_7  (port_state_in_7_2_7    ), //i
    .port_byte_out_0 (mul2_91_port_byte_out_0), //o
    .port_byte_out_1 (mul2_91_port_byte_out_1), //o
    .port_byte_out_2 (mul2_91_port_byte_out_2), //o
    .port_byte_out_3 (mul2_91_port_byte_out_3), //o
    .port_byte_out_4 (mul2_91_port_byte_out_4), //o
    .port_byte_out_5 (mul2_91_port_byte_out_5), //o
    .port_byte_out_6 (mul2_91_port_byte_out_6), //o
    .port_byte_out_7 (mul2_91_port_byte_out_7)  //o
  );
  Mul3 mul3_91 (
    .port_byte_in_0  (port_state_in_4_2_0    ), //i
    .port_byte_in_1  (port_state_in_4_2_1    ), //i
    .port_byte_in_2  (port_state_in_4_2_2    ), //i
    .port_byte_in_3  (port_state_in_4_2_3    ), //i
    .port_byte_in_4  (port_state_in_4_2_4    ), //i
    .port_byte_in_5  (port_state_in_4_2_5    ), //i
    .port_byte_in_6  (port_state_in_4_2_6    ), //i
    .port_byte_in_7  (port_state_in_4_2_7    ), //i
    .port_byte_out_0 (mul3_91_port_byte_out_0), //o
    .port_byte_out_1 (mul3_91_port_byte_out_1), //o
    .port_byte_out_2 (mul3_91_port_byte_out_2), //o
    .port_byte_out_3 (mul3_91_port_byte_out_3), //o
    .port_byte_out_4 (mul3_91_port_byte_out_4), //o
    .port_byte_out_5 (mul3_91_port_byte_out_5), //o
    .port_byte_out_6 (mul3_91_port_byte_out_6), //o
    .port_byte_out_7 (mul3_91_port_byte_out_7)  //o
  );
  Mul2 mul2_92 (
    .port_byte_in_0  (port_state_in_4_3_0    ), //i
    .port_byte_in_1  (port_state_in_4_3_1    ), //i
    .port_byte_in_2  (port_state_in_4_3_2    ), //i
    .port_byte_in_3  (port_state_in_4_3_3    ), //i
    .port_byte_in_4  (port_state_in_4_3_4    ), //i
    .port_byte_in_5  (port_state_in_4_3_5    ), //i
    .port_byte_in_6  (port_state_in_4_3_6    ), //i
    .port_byte_in_7  (port_state_in_4_3_7    ), //i
    .port_byte_out_0 (mul2_92_port_byte_out_0), //o
    .port_byte_out_1 (mul2_92_port_byte_out_1), //o
    .port_byte_out_2 (mul2_92_port_byte_out_2), //o
    .port_byte_out_3 (mul2_92_port_byte_out_3), //o
    .port_byte_out_4 (mul2_92_port_byte_out_4), //o
    .port_byte_out_5 (mul2_92_port_byte_out_5), //o
    .port_byte_out_6 (mul2_92_port_byte_out_6), //o
    .port_byte_out_7 (mul2_92_port_byte_out_7)  //o
  );
  Mul3 mul3_92 (
    .port_byte_in_0  (port_state_in_5_3_0    ), //i
    .port_byte_in_1  (port_state_in_5_3_1    ), //i
    .port_byte_in_2  (port_state_in_5_3_2    ), //i
    .port_byte_in_3  (port_state_in_5_3_3    ), //i
    .port_byte_in_4  (port_state_in_5_3_4    ), //i
    .port_byte_in_5  (port_state_in_5_3_5    ), //i
    .port_byte_in_6  (port_state_in_5_3_6    ), //i
    .port_byte_in_7  (port_state_in_5_3_7    ), //i
    .port_byte_out_0 (mul3_92_port_byte_out_0), //o
    .port_byte_out_1 (mul3_92_port_byte_out_1), //o
    .port_byte_out_2 (mul3_92_port_byte_out_2), //o
    .port_byte_out_3 (mul3_92_port_byte_out_3), //o
    .port_byte_out_4 (mul3_92_port_byte_out_4), //o
    .port_byte_out_5 (mul3_92_port_byte_out_5), //o
    .port_byte_out_6 (mul3_92_port_byte_out_6), //o
    .port_byte_out_7 (mul3_92_port_byte_out_7)  //o
  );
  Mul2 mul2_93 (
    .port_byte_in_0  (port_state_in_5_3_0    ), //i
    .port_byte_in_1  (port_state_in_5_3_1    ), //i
    .port_byte_in_2  (port_state_in_5_3_2    ), //i
    .port_byte_in_3  (port_state_in_5_3_3    ), //i
    .port_byte_in_4  (port_state_in_5_3_4    ), //i
    .port_byte_in_5  (port_state_in_5_3_5    ), //i
    .port_byte_in_6  (port_state_in_5_3_6    ), //i
    .port_byte_in_7  (port_state_in_5_3_7    ), //i
    .port_byte_out_0 (mul2_93_port_byte_out_0), //o
    .port_byte_out_1 (mul2_93_port_byte_out_1), //o
    .port_byte_out_2 (mul2_93_port_byte_out_2), //o
    .port_byte_out_3 (mul2_93_port_byte_out_3), //o
    .port_byte_out_4 (mul2_93_port_byte_out_4), //o
    .port_byte_out_5 (mul2_93_port_byte_out_5), //o
    .port_byte_out_6 (mul2_93_port_byte_out_6), //o
    .port_byte_out_7 (mul2_93_port_byte_out_7)  //o
  );
  Mul3 mul3_93 (
    .port_byte_in_0  (port_state_in_6_3_0    ), //i
    .port_byte_in_1  (port_state_in_6_3_1    ), //i
    .port_byte_in_2  (port_state_in_6_3_2    ), //i
    .port_byte_in_3  (port_state_in_6_3_3    ), //i
    .port_byte_in_4  (port_state_in_6_3_4    ), //i
    .port_byte_in_5  (port_state_in_6_3_5    ), //i
    .port_byte_in_6  (port_state_in_6_3_6    ), //i
    .port_byte_in_7  (port_state_in_6_3_7    ), //i
    .port_byte_out_0 (mul3_93_port_byte_out_0), //o
    .port_byte_out_1 (mul3_93_port_byte_out_1), //o
    .port_byte_out_2 (mul3_93_port_byte_out_2), //o
    .port_byte_out_3 (mul3_93_port_byte_out_3), //o
    .port_byte_out_4 (mul3_93_port_byte_out_4), //o
    .port_byte_out_5 (mul3_93_port_byte_out_5), //o
    .port_byte_out_6 (mul3_93_port_byte_out_6), //o
    .port_byte_out_7 (mul3_93_port_byte_out_7)  //o
  );
  Mul2 mul2_94 (
    .port_byte_in_0  (port_state_in_6_3_0    ), //i
    .port_byte_in_1  (port_state_in_6_3_1    ), //i
    .port_byte_in_2  (port_state_in_6_3_2    ), //i
    .port_byte_in_3  (port_state_in_6_3_3    ), //i
    .port_byte_in_4  (port_state_in_6_3_4    ), //i
    .port_byte_in_5  (port_state_in_6_3_5    ), //i
    .port_byte_in_6  (port_state_in_6_3_6    ), //i
    .port_byte_in_7  (port_state_in_6_3_7    ), //i
    .port_byte_out_0 (mul2_94_port_byte_out_0), //o
    .port_byte_out_1 (mul2_94_port_byte_out_1), //o
    .port_byte_out_2 (mul2_94_port_byte_out_2), //o
    .port_byte_out_3 (mul2_94_port_byte_out_3), //o
    .port_byte_out_4 (mul2_94_port_byte_out_4), //o
    .port_byte_out_5 (mul2_94_port_byte_out_5), //o
    .port_byte_out_6 (mul2_94_port_byte_out_6), //o
    .port_byte_out_7 (mul2_94_port_byte_out_7)  //o
  );
  Mul3 mul3_94 (
    .port_byte_in_0  (port_state_in_7_3_0    ), //i
    .port_byte_in_1  (port_state_in_7_3_1    ), //i
    .port_byte_in_2  (port_state_in_7_3_2    ), //i
    .port_byte_in_3  (port_state_in_7_3_3    ), //i
    .port_byte_in_4  (port_state_in_7_3_4    ), //i
    .port_byte_in_5  (port_state_in_7_3_5    ), //i
    .port_byte_in_6  (port_state_in_7_3_6    ), //i
    .port_byte_in_7  (port_state_in_7_3_7    ), //i
    .port_byte_out_0 (mul3_94_port_byte_out_0), //o
    .port_byte_out_1 (mul3_94_port_byte_out_1), //o
    .port_byte_out_2 (mul3_94_port_byte_out_2), //o
    .port_byte_out_3 (mul3_94_port_byte_out_3), //o
    .port_byte_out_4 (mul3_94_port_byte_out_4), //o
    .port_byte_out_5 (mul3_94_port_byte_out_5), //o
    .port_byte_out_6 (mul3_94_port_byte_out_6), //o
    .port_byte_out_7 (mul3_94_port_byte_out_7)  //o
  );
  Mul2 mul2_95 (
    .port_byte_in_0  (port_state_in_7_3_0    ), //i
    .port_byte_in_1  (port_state_in_7_3_1    ), //i
    .port_byte_in_2  (port_state_in_7_3_2    ), //i
    .port_byte_in_3  (port_state_in_7_3_3    ), //i
    .port_byte_in_4  (port_state_in_7_3_4    ), //i
    .port_byte_in_5  (port_state_in_7_3_5    ), //i
    .port_byte_in_6  (port_state_in_7_3_6    ), //i
    .port_byte_in_7  (port_state_in_7_3_7    ), //i
    .port_byte_out_0 (mul2_95_port_byte_out_0), //o
    .port_byte_out_1 (mul2_95_port_byte_out_1), //o
    .port_byte_out_2 (mul2_95_port_byte_out_2), //o
    .port_byte_out_3 (mul2_95_port_byte_out_3), //o
    .port_byte_out_4 (mul2_95_port_byte_out_4), //o
    .port_byte_out_5 (mul2_95_port_byte_out_5), //o
    .port_byte_out_6 (mul2_95_port_byte_out_6), //o
    .port_byte_out_7 (mul2_95_port_byte_out_7)  //o
  );
  Mul3 mul3_95 (
    .port_byte_in_0  (port_state_in_4_3_0    ), //i
    .port_byte_in_1  (port_state_in_4_3_1    ), //i
    .port_byte_in_2  (port_state_in_4_3_2    ), //i
    .port_byte_in_3  (port_state_in_4_3_3    ), //i
    .port_byte_in_4  (port_state_in_4_3_4    ), //i
    .port_byte_in_5  (port_state_in_4_3_5    ), //i
    .port_byte_in_6  (port_state_in_4_3_6    ), //i
    .port_byte_in_7  (port_state_in_4_3_7    ), //i
    .port_byte_out_0 (mul3_95_port_byte_out_0), //o
    .port_byte_out_1 (mul3_95_port_byte_out_1), //o
    .port_byte_out_2 (mul3_95_port_byte_out_2), //o
    .port_byte_out_3 (mul3_95_port_byte_out_3), //o
    .port_byte_out_4 (mul3_95_port_byte_out_4), //o
    .port_byte_out_5 (mul3_95_port_byte_out_5), //o
    .port_byte_out_6 (mul3_95_port_byte_out_6), //o
    .port_byte_out_7 (mul3_95_port_byte_out_7)  //o
  );
  Mul2 mul2_96 (
    .port_byte_in_0  (port_state_in_8_0_0    ), //i
    .port_byte_in_1  (port_state_in_8_0_1    ), //i
    .port_byte_in_2  (port_state_in_8_0_2    ), //i
    .port_byte_in_3  (port_state_in_8_0_3    ), //i
    .port_byte_in_4  (port_state_in_8_0_4    ), //i
    .port_byte_in_5  (port_state_in_8_0_5    ), //i
    .port_byte_in_6  (port_state_in_8_0_6    ), //i
    .port_byte_in_7  (port_state_in_8_0_7    ), //i
    .port_byte_out_0 (mul2_96_port_byte_out_0), //o
    .port_byte_out_1 (mul2_96_port_byte_out_1), //o
    .port_byte_out_2 (mul2_96_port_byte_out_2), //o
    .port_byte_out_3 (mul2_96_port_byte_out_3), //o
    .port_byte_out_4 (mul2_96_port_byte_out_4), //o
    .port_byte_out_5 (mul2_96_port_byte_out_5), //o
    .port_byte_out_6 (mul2_96_port_byte_out_6), //o
    .port_byte_out_7 (mul2_96_port_byte_out_7)  //o
  );
  Mul3 mul3_96 (
    .port_byte_in_0  (port_state_in_9_0_0    ), //i
    .port_byte_in_1  (port_state_in_9_0_1    ), //i
    .port_byte_in_2  (port_state_in_9_0_2    ), //i
    .port_byte_in_3  (port_state_in_9_0_3    ), //i
    .port_byte_in_4  (port_state_in_9_0_4    ), //i
    .port_byte_in_5  (port_state_in_9_0_5    ), //i
    .port_byte_in_6  (port_state_in_9_0_6    ), //i
    .port_byte_in_7  (port_state_in_9_0_7    ), //i
    .port_byte_out_0 (mul3_96_port_byte_out_0), //o
    .port_byte_out_1 (mul3_96_port_byte_out_1), //o
    .port_byte_out_2 (mul3_96_port_byte_out_2), //o
    .port_byte_out_3 (mul3_96_port_byte_out_3), //o
    .port_byte_out_4 (mul3_96_port_byte_out_4), //o
    .port_byte_out_5 (mul3_96_port_byte_out_5), //o
    .port_byte_out_6 (mul3_96_port_byte_out_6), //o
    .port_byte_out_7 (mul3_96_port_byte_out_7)  //o
  );
  Mul2 mul2_97 (
    .port_byte_in_0  (port_state_in_9_0_0    ), //i
    .port_byte_in_1  (port_state_in_9_0_1    ), //i
    .port_byte_in_2  (port_state_in_9_0_2    ), //i
    .port_byte_in_3  (port_state_in_9_0_3    ), //i
    .port_byte_in_4  (port_state_in_9_0_4    ), //i
    .port_byte_in_5  (port_state_in_9_0_5    ), //i
    .port_byte_in_6  (port_state_in_9_0_6    ), //i
    .port_byte_in_7  (port_state_in_9_0_7    ), //i
    .port_byte_out_0 (mul2_97_port_byte_out_0), //o
    .port_byte_out_1 (mul2_97_port_byte_out_1), //o
    .port_byte_out_2 (mul2_97_port_byte_out_2), //o
    .port_byte_out_3 (mul2_97_port_byte_out_3), //o
    .port_byte_out_4 (mul2_97_port_byte_out_4), //o
    .port_byte_out_5 (mul2_97_port_byte_out_5), //o
    .port_byte_out_6 (mul2_97_port_byte_out_6), //o
    .port_byte_out_7 (mul2_97_port_byte_out_7)  //o
  );
  Mul3 mul3_97 (
    .port_byte_in_0  (port_state_in_10_0_0   ), //i
    .port_byte_in_1  (port_state_in_10_0_1   ), //i
    .port_byte_in_2  (port_state_in_10_0_2   ), //i
    .port_byte_in_3  (port_state_in_10_0_3   ), //i
    .port_byte_in_4  (port_state_in_10_0_4   ), //i
    .port_byte_in_5  (port_state_in_10_0_5   ), //i
    .port_byte_in_6  (port_state_in_10_0_6   ), //i
    .port_byte_in_7  (port_state_in_10_0_7   ), //i
    .port_byte_out_0 (mul3_97_port_byte_out_0), //o
    .port_byte_out_1 (mul3_97_port_byte_out_1), //o
    .port_byte_out_2 (mul3_97_port_byte_out_2), //o
    .port_byte_out_3 (mul3_97_port_byte_out_3), //o
    .port_byte_out_4 (mul3_97_port_byte_out_4), //o
    .port_byte_out_5 (mul3_97_port_byte_out_5), //o
    .port_byte_out_6 (mul3_97_port_byte_out_6), //o
    .port_byte_out_7 (mul3_97_port_byte_out_7)  //o
  );
  Mul2 mul2_98 (
    .port_byte_in_0  (port_state_in_10_0_0   ), //i
    .port_byte_in_1  (port_state_in_10_0_1   ), //i
    .port_byte_in_2  (port_state_in_10_0_2   ), //i
    .port_byte_in_3  (port_state_in_10_0_3   ), //i
    .port_byte_in_4  (port_state_in_10_0_4   ), //i
    .port_byte_in_5  (port_state_in_10_0_5   ), //i
    .port_byte_in_6  (port_state_in_10_0_6   ), //i
    .port_byte_in_7  (port_state_in_10_0_7   ), //i
    .port_byte_out_0 (mul2_98_port_byte_out_0), //o
    .port_byte_out_1 (mul2_98_port_byte_out_1), //o
    .port_byte_out_2 (mul2_98_port_byte_out_2), //o
    .port_byte_out_3 (mul2_98_port_byte_out_3), //o
    .port_byte_out_4 (mul2_98_port_byte_out_4), //o
    .port_byte_out_5 (mul2_98_port_byte_out_5), //o
    .port_byte_out_6 (mul2_98_port_byte_out_6), //o
    .port_byte_out_7 (mul2_98_port_byte_out_7)  //o
  );
  Mul3 mul3_98 (
    .port_byte_in_0  (port_state_in_11_0_0   ), //i
    .port_byte_in_1  (port_state_in_11_0_1   ), //i
    .port_byte_in_2  (port_state_in_11_0_2   ), //i
    .port_byte_in_3  (port_state_in_11_0_3   ), //i
    .port_byte_in_4  (port_state_in_11_0_4   ), //i
    .port_byte_in_5  (port_state_in_11_0_5   ), //i
    .port_byte_in_6  (port_state_in_11_0_6   ), //i
    .port_byte_in_7  (port_state_in_11_0_7   ), //i
    .port_byte_out_0 (mul3_98_port_byte_out_0), //o
    .port_byte_out_1 (mul3_98_port_byte_out_1), //o
    .port_byte_out_2 (mul3_98_port_byte_out_2), //o
    .port_byte_out_3 (mul3_98_port_byte_out_3), //o
    .port_byte_out_4 (mul3_98_port_byte_out_4), //o
    .port_byte_out_5 (mul3_98_port_byte_out_5), //o
    .port_byte_out_6 (mul3_98_port_byte_out_6), //o
    .port_byte_out_7 (mul3_98_port_byte_out_7)  //o
  );
  Mul2 mul2_99 (
    .port_byte_in_0  (port_state_in_11_0_0   ), //i
    .port_byte_in_1  (port_state_in_11_0_1   ), //i
    .port_byte_in_2  (port_state_in_11_0_2   ), //i
    .port_byte_in_3  (port_state_in_11_0_3   ), //i
    .port_byte_in_4  (port_state_in_11_0_4   ), //i
    .port_byte_in_5  (port_state_in_11_0_5   ), //i
    .port_byte_in_6  (port_state_in_11_0_6   ), //i
    .port_byte_in_7  (port_state_in_11_0_7   ), //i
    .port_byte_out_0 (mul2_99_port_byte_out_0), //o
    .port_byte_out_1 (mul2_99_port_byte_out_1), //o
    .port_byte_out_2 (mul2_99_port_byte_out_2), //o
    .port_byte_out_3 (mul2_99_port_byte_out_3), //o
    .port_byte_out_4 (mul2_99_port_byte_out_4), //o
    .port_byte_out_5 (mul2_99_port_byte_out_5), //o
    .port_byte_out_6 (mul2_99_port_byte_out_6), //o
    .port_byte_out_7 (mul2_99_port_byte_out_7)  //o
  );
  Mul3 mul3_99 (
    .port_byte_in_0  (port_state_in_8_0_0    ), //i
    .port_byte_in_1  (port_state_in_8_0_1    ), //i
    .port_byte_in_2  (port_state_in_8_0_2    ), //i
    .port_byte_in_3  (port_state_in_8_0_3    ), //i
    .port_byte_in_4  (port_state_in_8_0_4    ), //i
    .port_byte_in_5  (port_state_in_8_0_5    ), //i
    .port_byte_in_6  (port_state_in_8_0_6    ), //i
    .port_byte_in_7  (port_state_in_8_0_7    ), //i
    .port_byte_out_0 (mul3_99_port_byte_out_0), //o
    .port_byte_out_1 (mul3_99_port_byte_out_1), //o
    .port_byte_out_2 (mul3_99_port_byte_out_2), //o
    .port_byte_out_3 (mul3_99_port_byte_out_3), //o
    .port_byte_out_4 (mul3_99_port_byte_out_4), //o
    .port_byte_out_5 (mul3_99_port_byte_out_5), //o
    .port_byte_out_6 (mul3_99_port_byte_out_6), //o
    .port_byte_out_7 (mul3_99_port_byte_out_7)  //o
  );
  Mul2 mul2_100 (
    .port_byte_in_0  (port_state_in_8_1_0     ), //i
    .port_byte_in_1  (port_state_in_8_1_1     ), //i
    .port_byte_in_2  (port_state_in_8_1_2     ), //i
    .port_byte_in_3  (port_state_in_8_1_3     ), //i
    .port_byte_in_4  (port_state_in_8_1_4     ), //i
    .port_byte_in_5  (port_state_in_8_1_5     ), //i
    .port_byte_in_6  (port_state_in_8_1_6     ), //i
    .port_byte_in_7  (port_state_in_8_1_7     ), //i
    .port_byte_out_0 (mul2_100_port_byte_out_0), //o
    .port_byte_out_1 (mul2_100_port_byte_out_1), //o
    .port_byte_out_2 (mul2_100_port_byte_out_2), //o
    .port_byte_out_3 (mul2_100_port_byte_out_3), //o
    .port_byte_out_4 (mul2_100_port_byte_out_4), //o
    .port_byte_out_5 (mul2_100_port_byte_out_5), //o
    .port_byte_out_6 (mul2_100_port_byte_out_6), //o
    .port_byte_out_7 (mul2_100_port_byte_out_7)  //o
  );
  Mul3 mul3_100 (
    .port_byte_in_0  (port_state_in_9_1_0     ), //i
    .port_byte_in_1  (port_state_in_9_1_1     ), //i
    .port_byte_in_2  (port_state_in_9_1_2     ), //i
    .port_byte_in_3  (port_state_in_9_1_3     ), //i
    .port_byte_in_4  (port_state_in_9_1_4     ), //i
    .port_byte_in_5  (port_state_in_9_1_5     ), //i
    .port_byte_in_6  (port_state_in_9_1_6     ), //i
    .port_byte_in_7  (port_state_in_9_1_7     ), //i
    .port_byte_out_0 (mul3_100_port_byte_out_0), //o
    .port_byte_out_1 (mul3_100_port_byte_out_1), //o
    .port_byte_out_2 (mul3_100_port_byte_out_2), //o
    .port_byte_out_3 (mul3_100_port_byte_out_3), //o
    .port_byte_out_4 (mul3_100_port_byte_out_4), //o
    .port_byte_out_5 (mul3_100_port_byte_out_5), //o
    .port_byte_out_6 (mul3_100_port_byte_out_6), //o
    .port_byte_out_7 (mul3_100_port_byte_out_7)  //o
  );
  Mul2 mul2_101 (
    .port_byte_in_0  (port_state_in_9_1_0     ), //i
    .port_byte_in_1  (port_state_in_9_1_1     ), //i
    .port_byte_in_2  (port_state_in_9_1_2     ), //i
    .port_byte_in_3  (port_state_in_9_1_3     ), //i
    .port_byte_in_4  (port_state_in_9_1_4     ), //i
    .port_byte_in_5  (port_state_in_9_1_5     ), //i
    .port_byte_in_6  (port_state_in_9_1_6     ), //i
    .port_byte_in_7  (port_state_in_9_1_7     ), //i
    .port_byte_out_0 (mul2_101_port_byte_out_0), //o
    .port_byte_out_1 (mul2_101_port_byte_out_1), //o
    .port_byte_out_2 (mul2_101_port_byte_out_2), //o
    .port_byte_out_3 (mul2_101_port_byte_out_3), //o
    .port_byte_out_4 (mul2_101_port_byte_out_4), //o
    .port_byte_out_5 (mul2_101_port_byte_out_5), //o
    .port_byte_out_6 (mul2_101_port_byte_out_6), //o
    .port_byte_out_7 (mul2_101_port_byte_out_7)  //o
  );
  Mul3 mul3_101 (
    .port_byte_in_0  (port_state_in_10_1_0    ), //i
    .port_byte_in_1  (port_state_in_10_1_1    ), //i
    .port_byte_in_2  (port_state_in_10_1_2    ), //i
    .port_byte_in_3  (port_state_in_10_1_3    ), //i
    .port_byte_in_4  (port_state_in_10_1_4    ), //i
    .port_byte_in_5  (port_state_in_10_1_5    ), //i
    .port_byte_in_6  (port_state_in_10_1_6    ), //i
    .port_byte_in_7  (port_state_in_10_1_7    ), //i
    .port_byte_out_0 (mul3_101_port_byte_out_0), //o
    .port_byte_out_1 (mul3_101_port_byte_out_1), //o
    .port_byte_out_2 (mul3_101_port_byte_out_2), //o
    .port_byte_out_3 (mul3_101_port_byte_out_3), //o
    .port_byte_out_4 (mul3_101_port_byte_out_4), //o
    .port_byte_out_5 (mul3_101_port_byte_out_5), //o
    .port_byte_out_6 (mul3_101_port_byte_out_6), //o
    .port_byte_out_7 (mul3_101_port_byte_out_7)  //o
  );
  Mul2 mul2_102 (
    .port_byte_in_0  (port_state_in_10_1_0    ), //i
    .port_byte_in_1  (port_state_in_10_1_1    ), //i
    .port_byte_in_2  (port_state_in_10_1_2    ), //i
    .port_byte_in_3  (port_state_in_10_1_3    ), //i
    .port_byte_in_4  (port_state_in_10_1_4    ), //i
    .port_byte_in_5  (port_state_in_10_1_5    ), //i
    .port_byte_in_6  (port_state_in_10_1_6    ), //i
    .port_byte_in_7  (port_state_in_10_1_7    ), //i
    .port_byte_out_0 (mul2_102_port_byte_out_0), //o
    .port_byte_out_1 (mul2_102_port_byte_out_1), //o
    .port_byte_out_2 (mul2_102_port_byte_out_2), //o
    .port_byte_out_3 (mul2_102_port_byte_out_3), //o
    .port_byte_out_4 (mul2_102_port_byte_out_4), //o
    .port_byte_out_5 (mul2_102_port_byte_out_5), //o
    .port_byte_out_6 (mul2_102_port_byte_out_6), //o
    .port_byte_out_7 (mul2_102_port_byte_out_7)  //o
  );
  Mul3 mul3_102 (
    .port_byte_in_0  (port_state_in_11_1_0    ), //i
    .port_byte_in_1  (port_state_in_11_1_1    ), //i
    .port_byte_in_2  (port_state_in_11_1_2    ), //i
    .port_byte_in_3  (port_state_in_11_1_3    ), //i
    .port_byte_in_4  (port_state_in_11_1_4    ), //i
    .port_byte_in_5  (port_state_in_11_1_5    ), //i
    .port_byte_in_6  (port_state_in_11_1_6    ), //i
    .port_byte_in_7  (port_state_in_11_1_7    ), //i
    .port_byte_out_0 (mul3_102_port_byte_out_0), //o
    .port_byte_out_1 (mul3_102_port_byte_out_1), //o
    .port_byte_out_2 (mul3_102_port_byte_out_2), //o
    .port_byte_out_3 (mul3_102_port_byte_out_3), //o
    .port_byte_out_4 (mul3_102_port_byte_out_4), //o
    .port_byte_out_5 (mul3_102_port_byte_out_5), //o
    .port_byte_out_6 (mul3_102_port_byte_out_6), //o
    .port_byte_out_7 (mul3_102_port_byte_out_7)  //o
  );
  Mul2 mul2_103 (
    .port_byte_in_0  (port_state_in_11_1_0    ), //i
    .port_byte_in_1  (port_state_in_11_1_1    ), //i
    .port_byte_in_2  (port_state_in_11_1_2    ), //i
    .port_byte_in_3  (port_state_in_11_1_3    ), //i
    .port_byte_in_4  (port_state_in_11_1_4    ), //i
    .port_byte_in_5  (port_state_in_11_1_5    ), //i
    .port_byte_in_6  (port_state_in_11_1_6    ), //i
    .port_byte_in_7  (port_state_in_11_1_7    ), //i
    .port_byte_out_0 (mul2_103_port_byte_out_0), //o
    .port_byte_out_1 (mul2_103_port_byte_out_1), //o
    .port_byte_out_2 (mul2_103_port_byte_out_2), //o
    .port_byte_out_3 (mul2_103_port_byte_out_3), //o
    .port_byte_out_4 (mul2_103_port_byte_out_4), //o
    .port_byte_out_5 (mul2_103_port_byte_out_5), //o
    .port_byte_out_6 (mul2_103_port_byte_out_6), //o
    .port_byte_out_7 (mul2_103_port_byte_out_7)  //o
  );
  Mul3 mul3_103 (
    .port_byte_in_0  (port_state_in_8_1_0     ), //i
    .port_byte_in_1  (port_state_in_8_1_1     ), //i
    .port_byte_in_2  (port_state_in_8_1_2     ), //i
    .port_byte_in_3  (port_state_in_8_1_3     ), //i
    .port_byte_in_4  (port_state_in_8_1_4     ), //i
    .port_byte_in_5  (port_state_in_8_1_5     ), //i
    .port_byte_in_6  (port_state_in_8_1_6     ), //i
    .port_byte_in_7  (port_state_in_8_1_7     ), //i
    .port_byte_out_0 (mul3_103_port_byte_out_0), //o
    .port_byte_out_1 (mul3_103_port_byte_out_1), //o
    .port_byte_out_2 (mul3_103_port_byte_out_2), //o
    .port_byte_out_3 (mul3_103_port_byte_out_3), //o
    .port_byte_out_4 (mul3_103_port_byte_out_4), //o
    .port_byte_out_5 (mul3_103_port_byte_out_5), //o
    .port_byte_out_6 (mul3_103_port_byte_out_6), //o
    .port_byte_out_7 (mul3_103_port_byte_out_7)  //o
  );
  Mul2 mul2_104 (
    .port_byte_in_0  (port_state_in_8_2_0     ), //i
    .port_byte_in_1  (port_state_in_8_2_1     ), //i
    .port_byte_in_2  (port_state_in_8_2_2     ), //i
    .port_byte_in_3  (port_state_in_8_2_3     ), //i
    .port_byte_in_4  (port_state_in_8_2_4     ), //i
    .port_byte_in_5  (port_state_in_8_2_5     ), //i
    .port_byte_in_6  (port_state_in_8_2_6     ), //i
    .port_byte_in_7  (port_state_in_8_2_7     ), //i
    .port_byte_out_0 (mul2_104_port_byte_out_0), //o
    .port_byte_out_1 (mul2_104_port_byte_out_1), //o
    .port_byte_out_2 (mul2_104_port_byte_out_2), //o
    .port_byte_out_3 (mul2_104_port_byte_out_3), //o
    .port_byte_out_4 (mul2_104_port_byte_out_4), //o
    .port_byte_out_5 (mul2_104_port_byte_out_5), //o
    .port_byte_out_6 (mul2_104_port_byte_out_6), //o
    .port_byte_out_7 (mul2_104_port_byte_out_7)  //o
  );
  Mul3 mul3_104 (
    .port_byte_in_0  (port_state_in_9_2_0     ), //i
    .port_byte_in_1  (port_state_in_9_2_1     ), //i
    .port_byte_in_2  (port_state_in_9_2_2     ), //i
    .port_byte_in_3  (port_state_in_9_2_3     ), //i
    .port_byte_in_4  (port_state_in_9_2_4     ), //i
    .port_byte_in_5  (port_state_in_9_2_5     ), //i
    .port_byte_in_6  (port_state_in_9_2_6     ), //i
    .port_byte_in_7  (port_state_in_9_2_7     ), //i
    .port_byte_out_0 (mul3_104_port_byte_out_0), //o
    .port_byte_out_1 (mul3_104_port_byte_out_1), //o
    .port_byte_out_2 (mul3_104_port_byte_out_2), //o
    .port_byte_out_3 (mul3_104_port_byte_out_3), //o
    .port_byte_out_4 (mul3_104_port_byte_out_4), //o
    .port_byte_out_5 (mul3_104_port_byte_out_5), //o
    .port_byte_out_6 (mul3_104_port_byte_out_6), //o
    .port_byte_out_7 (mul3_104_port_byte_out_7)  //o
  );
  Mul2 mul2_105 (
    .port_byte_in_0  (port_state_in_9_2_0     ), //i
    .port_byte_in_1  (port_state_in_9_2_1     ), //i
    .port_byte_in_2  (port_state_in_9_2_2     ), //i
    .port_byte_in_3  (port_state_in_9_2_3     ), //i
    .port_byte_in_4  (port_state_in_9_2_4     ), //i
    .port_byte_in_5  (port_state_in_9_2_5     ), //i
    .port_byte_in_6  (port_state_in_9_2_6     ), //i
    .port_byte_in_7  (port_state_in_9_2_7     ), //i
    .port_byte_out_0 (mul2_105_port_byte_out_0), //o
    .port_byte_out_1 (mul2_105_port_byte_out_1), //o
    .port_byte_out_2 (mul2_105_port_byte_out_2), //o
    .port_byte_out_3 (mul2_105_port_byte_out_3), //o
    .port_byte_out_4 (mul2_105_port_byte_out_4), //o
    .port_byte_out_5 (mul2_105_port_byte_out_5), //o
    .port_byte_out_6 (mul2_105_port_byte_out_6), //o
    .port_byte_out_7 (mul2_105_port_byte_out_7)  //o
  );
  Mul3 mul3_105 (
    .port_byte_in_0  (port_state_in_10_2_0    ), //i
    .port_byte_in_1  (port_state_in_10_2_1    ), //i
    .port_byte_in_2  (port_state_in_10_2_2    ), //i
    .port_byte_in_3  (port_state_in_10_2_3    ), //i
    .port_byte_in_4  (port_state_in_10_2_4    ), //i
    .port_byte_in_5  (port_state_in_10_2_5    ), //i
    .port_byte_in_6  (port_state_in_10_2_6    ), //i
    .port_byte_in_7  (port_state_in_10_2_7    ), //i
    .port_byte_out_0 (mul3_105_port_byte_out_0), //o
    .port_byte_out_1 (mul3_105_port_byte_out_1), //o
    .port_byte_out_2 (mul3_105_port_byte_out_2), //o
    .port_byte_out_3 (mul3_105_port_byte_out_3), //o
    .port_byte_out_4 (mul3_105_port_byte_out_4), //o
    .port_byte_out_5 (mul3_105_port_byte_out_5), //o
    .port_byte_out_6 (mul3_105_port_byte_out_6), //o
    .port_byte_out_7 (mul3_105_port_byte_out_7)  //o
  );
  Mul2 mul2_106 (
    .port_byte_in_0  (port_state_in_10_2_0    ), //i
    .port_byte_in_1  (port_state_in_10_2_1    ), //i
    .port_byte_in_2  (port_state_in_10_2_2    ), //i
    .port_byte_in_3  (port_state_in_10_2_3    ), //i
    .port_byte_in_4  (port_state_in_10_2_4    ), //i
    .port_byte_in_5  (port_state_in_10_2_5    ), //i
    .port_byte_in_6  (port_state_in_10_2_6    ), //i
    .port_byte_in_7  (port_state_in_10_2_7    ), //i
    .port_byte_out_0 (mul2_106_port_byte_out_0), //o
    .port_byte_out_1 (mul2_106_port_byte_out_1), //o
    .port_byte_out_2 (mul2_106_port_byte_out_2), //o
    .port_byte_out_3 (mul2_106_port_byte_out_3), //o
    .port_byte_out_4 (mul2_106_port_byte_out_4), //o
    .port_byte_out_5 (mul2_106_port_byte_out_5), //o
    .port_byte_out_6 (mul2_106_port_byte_out_6), //o
    .port_byte_out_7 (mul2_106_port_byte_out_7)  //o
  );
  Mul3 mul3_106 (
    .port_byte_in_0  (port_state_in_11_2_0    ), //i
    .port_byte_in_1  (port_state_in_11_2_1    ), //i
    .port_byte_in_2  (port_state_in_11_2_2    ), //i
    .port_byte_in_3  (port_state_in_11_2_3    ), //i
    .port_byte_in_4  (port_state_in_11_2_4    ), //i
    .port_byte_in_5  (port_state_in_11_2_5    ), //i
    .port_byte_in_6  (port_state_in_11_2_6    ), //i
    .port_byte_in_7  (port_state_in_11_2_7    ), //i
    .port_byte_out_0 (mul3_106_port_byte_out_0), //o
    .port_byte_out_1 (mul3_106_port_byte_out_1), //o
    .port_byte_out_2 (mul3_106_port_byte_out_2), //o
    .port_byte_out_3 (mul3_106_port_byte_out_3), //o
    .port_byte_out_4 (mul3_106_port_byte_out_4), //o
    .port_byte_out_5 (mul3_106_port_byte_out_5), //o
    .port_byte_out_6 (mul3_106_port_byte_out_6), //o
    .port_byte_out_7 (mul3_106_port_byte_out_7)  //o
  );
  Mul2 mul2_107 (
    .port_byte_in_0  (port_state_in_11_2_0    ), //i
    .port_byte_in_1  (port_state_in_11_2_1    ), //i
    .port_byte_in_2  (port_state_in_11_2_2    ), //i
    .port_byte_in_3  (port_state_in_11_2_3    ), //i
    .port_byte_in_4  (port_state_in_11_2_4    ), //i
    .port_byte_in_5  (port_state_in_11_2_5    ), //i
    .port_byte_in_6  (port_state_in_11_2_6    ), //i
    .port_byte_in_7  (port_state_in_11_2_7    ), //i
    .port_byte_out_0 (mul2_107_port_byte_out_0), //o
    .port_byte_out_1 (mul2_107_port_byte_out_1), //o
    .port_byte_out_2 (mul2_107_port_byte_out_2), //o
    .port_byte_out_3 (mul2_107_port_byte_out_3), //o
    .port_byte_out_4 (mul2_107_port_byte_out_4), //o
    .port_byte_out_5 (mul2_107_port_byte_out_5), //o
    .port_byte_out_6 (mul2_107_port_byte_out_6), //o
    .port_byte_out_7 (mul2_107_port_byte_out_7)  //o
  );
  Mul3 mul3_107 (
    .port_byte_in_0  (port_state_in_8_2_0     ), //i
    .port_byte_in_1  (port_state_in_8_2_1     ), //i
    .port_byte_in_2  (port_state_in_8_2_2     ), //i
    .port_byte_in_3  (port_state_in_8_2_3     ), //i
    .port_byte_in_4  (port_state_in_8_2_4     ), //i
    .port_byte_in_5  (port_state_in_8_2_5     ), //i
    .port_byte_in_6  (port_state_in_8_2_6     ), //i
    .port_byte_in_7  (port_state_in_8_2_7     ), //i
    .port_byte_out_0 (mul3_107_port_byte_out_0), //o
    .port_byte_out_1 (mul3_107_port_byte_out_1), //o
    .port_byte_out_2 (mul3_107_port_byte_out_2), //o
    .port_byte_out_3 (mul3_107_port_byte_out_3), //o
    .port_byte_out_4 (mul3_107_port_byte_out_4), //o
    .port_byte_out_5 (mul3_107_port_byte_out_5), //o
    .port_byte_out_6 (mul3_107_port_byte_out_6), //o
    .port_byte_out_7 (mul3_107_port_byte_out_7)  //o
  );
  Mul2 mul2_108 (
    .port_byte_in_0  (port_state_in_8_3_0     ), //i
    .port_byte_in_1  (port_state_in_8_3_1     ), //i
    .port_byte_in_2  (port_state_in_8_3_2     ), //i
    .port_byte_in_3  (port_state_in_8_3_3     ), //i
    .port_byte_in_4  (port_state_in_8_3_4     ), //i
    .port_byte_in_5  (port_state_in_8_3_5     ), //i
    .port_byte_in_6  (port_state_in_8_3_6     ), //i
    .port_byte_in_7  (port_state_in_8_3_7     ), //i
    .port_byte_out_0 (mul2_108_port_byte_out_0), //o
    .port_byte_out_1 (mul2_108_port_byte_out_1), //o
    .port_byte_out_2 (mul2_108_port_byte_out_2), //o
    .port_byte_out_3 (mul2_108_port_byte_out_3), //o
    .port_byte_out_4 (mul2_108_port_byte_out_4), //o
    .port_byte_out_5 (mul2_108_port_byte_out_5), //o
    .port_byte_out_6 (mul2_108_port_byte_out_6), //o
    .port_byte_out_7 (mul2_108_port_byte_out_7)  //o
  );
  Mul3 mul3_108 (
    .port_byte_in_0  (port_state_in_9_3_0     ), //i
    .port_byte_in_1  (port_state_in_9_3_1     ), //i
    .port_byte_in_2  (port_state_in_9_3_2     ), //i
    .port_byte_in_3  (port_state_in_9_3_3     ), //i
    .port_byte_in_4  (port_state_in_9_3_4     ), //i
    .port_byte_in_5  (port_state_in_9_3_5     ), //i
    .port_byte_in_6  (port_state_in_9_3_6     ), //i
    .port_byte_in_7  (port_state_in_9_3_7     ), //i
    .port_byte_out_0 (mul3_108_port_byte_out_0), //o
    .port_byte_out_1 (mul3_108_port_byte_out_1), //o
    .port_byte_out_2 (mul3_108_port_byte_out_2), //o
    .port_byte_out_3 (mul3_108_port_byte_out_3), //o
    .port_byte_out_4 (mul3_108_port_byte_out_4), //o
    .port_byte_out_5 (mul3_108_port_byte_out_5), //o
    .port_byte_out_6 (mul3_108_port_byte_out_6), //o
    .port_byte_out_7 (mul3_108_port_byte_out_7)  //o
  );
  Mul2 mul2_109 (
    .port_byte_in_0  (port_state_in_9_3_0     ), //i
    .port_byte_in_1  (port_state_in_9_3_1     ), //i
    .port_byte_in_2  (port_state_in_9_3_2     ), //i
    .port_byte_in_3  (port_state_in_9_3_3     ), //i
    .port_byte_in_4  (port_state_in_9_3_4     ), //i
    .port_byte_in_5  (port_state_in_9_3_5     ), //i
    .port_byte_in_6  (port_state_in_9_3_6     ), //i
    .port_byte_in_7  (port_state_in_9_3_7     ), //i
    .port_byte_out_0 (mul2_109_port_byte_out_0), //o
    .port_byte_out_1 (mul2_109_port_byte_out_1), //o
    .port_byte_out_2 (mul2_109_port_byte_out_2), //o
    .port_byte_out_3 (mul2_109_port_byte_out_3), //o
    .port_byte_out_4 (mul2_109_port_byte_out_4), //o
    .port_byte_out_5 (mul2_109_port_byte_out_5), //o
    .port_byte_out_6 (mul2_109_port_byte_out_6), //o
    .port_byte_out_7 (mul2_109_port_byte_out_7)  //o
  );
  Mul3 mul3_109 (
    .port_byte_in_0  (port_state_in_10_3_0    ), //i
    .port_byte_in_1  (port_state_in_10_3_1    ), //i
    .port_byte_in_2  (port_state_in_10_3_2    ), //i
    .port_byte_in_3  (port_state_in_10_3_3    ), //i
    .port_byte_in_4  (port_state_in_10_3_4    ), //i
    .port_byte_in_5  (port_state_in_10_3_5    ), //i
    .port_byte_in_6  (port_state_in_10_3_6    ), //i
    .port_byte_in_7  (port_state_in_10_3_7    ), //i
    .port_byte_out_0 (mul3_109_port_byte_out_0), //o
    .port_byte_out_1 (mul3_109_port_byte_out_1), //o
    .port_byte_out_2 (mul3_109_port_byte_out_2), //o
    .port_byte_out_3 (mul3_109_port_byte_out_3), //o
    .port_byte_out_4 (mul3_109_port_byte_out_4), //o
    .port_byte_out_5 (mul3_109_port_byte_out_5), //o
    .port_byte_out_6 (mul3_109_port_byte_out_6), //o
    .port_byte_out_7 (mul3_109_port_byte_out_7)  //o
  );
  Mul2 mul2_110 (
    .port_byte_in_0  (port_state_in_10_3_0    ), //i
    .port_byte_in_1  (port_state_in_10_3_1    ), //i
    .port_byte_in_2  (port_state_in_10_3_2    ), //i
    .port_byte_in_3  (port_state_in_10_3_3    ), //i
    .port_byte_in_4  (port_state_in_10_3_4    ), //i
    .port_byte_in_5  (port_state_in_10_3_5    ), //i
    .port_byte_in_6  (port_state_in_10_3_6    ), //i
    .port_byte_in_7  (port_state_in_10_3_7    ), //i
    .port_byte_out_0 (mul2_110_port_byte_out_0), //o
    .port_byte_out_1 (mul2_110_port_byte_out_1), //o
    .port_byte_out_2 (mul2_110_port_byte_out_2), //o
    .port_byte_out_3 (mul2_110_port_byte_out_3), //o
    .port_byte_out_4 (mul2_110_port_byte_out_4), //o
    .port_byte_out_5 (mul2_110_port_byte_out_5), //o
    .port_byte_out_6 (mul2_110_port_byte_out_6), //o
    .port_byte_out_7 (mul2_110_port_byte_out_7)  //o
  );
  Mul3 mul3_110 (
    .port_byte_in_0  (port_state_in_11_3_0    ), //i
    .port_byte_in_1  (port_state_in_11_3_1    ), //i
    .port_byte_in_2  (port_state_in_11_3_2    ), //i
    .port_byte_in_3  (port_state_in_11_3_3    ), //i
    .port_byte_in_4  (port_state_in_11_3_4    ), //i
    .port_byte_in_5  (port_state_in_11_3_5    ), //i
    .port_byte_in_6  (port_state_in_11_3_6    ), //i
    .port_byte_in_7  (port_state_in_11_3_7    ), //i
    .port_byte_out_0 (mul3_110_port_byte_out_0), //o
    .port_byte_out_1 (mul3_110_port_byte_out_1), //o
    .port_byte_out_2 (mul3_110_port_byte_out_2), //o
    .port_byte_out_3 (mul3_110_port_byte_out_3), //o
    .port_byte_out_4 (mul3_110_port_byte_out_4), //o
    .port_byte_out_5 (mul3_110_port_byte_out_5), //o
    .port_byte_out_6 (mul3_110_port_byte_out_6), //o
    .port_byte_out_7 (mul3_110_port_byte_out_7)  //o
  );
  Mul2 mul2_111 (
    .port_byte_in_0  (port_state_in_11_3_0    ), //i
    .port_byte_in_1  (port_state_in_11_3_1    ), //i
    .port_byte_in_2  (port_state_in_11_3_2    ), //i
    .port_byte_in_3  (port_state_in_11_3_3    ), //i
    .port_byte_in_4  (port_state_in_11_3_4    ), //i
    .port_byte_in_5  (port_state_in_11_3_5    ), //i
    .port_byte_in_6  (port_state_in_11_3_6    ), //i
    .port_byte_in_7  (port_state_in_11_3_7    ), //i
    .port_byte_out_0 (mul2_111_port_byte_out_0), //o
    .port_byte_out_1 (mul2_111_port_byte_out_1), //o
    .port_byte_out_2 (mul2_111_port_byte_out_2), //o
    .port_byte_out_3 (mul2_111_port_byte_out_3), //o
    .port_byte_out_4 (mul2_111_port_byte_out_4), //o
    .port_byte_out_5 (mul2_111_port_byte_out_5), //o
    .port_byte_out_6 (mul2_111_port_byte_out_6), //o
    .port_byte_out_7 (mul2_111_port_byte_out_7)  //o
  );
  Mul3 mul3_111 (
    .port_byte_in_0  (port_state_in_8_3_0     ), //i
    .port_byte_in_1  (port_state_in_8_3_1     ), //i
    .port_byte_in_2  (port_state_in_8_3_2     ), //i
    .port_byte_in_3  (port_state_in_8_3_3     ), //i
    .port_byte_in_4  (port_state_in_8_3_4     ), //i
    .port_byte_in_5  (port_state_in_8_3_5     ), //i
    .port_byte_in_6  (port_state_in_8_3_6     ), //i
    .port_byte_in_7  (port_state_in_8_3_7     ), //i
    .port_byte_out_0 (mul3_111_port_byte_out_0), //o
    .port_byte_out_1 (mul3_111_port_byte_out_1), //o
    .port_byte_out_2 (mul3_111_port_byte_out_2), //o
    .port_byte_out_3 (mul3_111_port_byte_out_3), //o
    .port_byte_out_4 (mul3_111_port_byte_out_4), //o
    .port_byte_out_5 (mul3_111_port_byte_out_5), //o
    .port_byte_out_6 (mul3_111_port_byte_out_6), //o
    .port_byte_out_7 (mul3_111_port_byte_out_7)  //o
  );
  Mul2 mul2_112 (
    .port_byte_in_0  (port_state_in_12_0_0    ), //i
    .port_byte_in_1  (port_state_in_12_0_1    ), //i
    .port_byte_in_2  (port_state_in_12_0_2    ), //i
    .port_byte_in_3  (port_state_in_12_0_3    ), //i
    .port_byte_in_4  (port_state_in_12_0_4    ), //i
    .port_byte_in_5  (port_state_in_12_0_5    ), //i
    .port_byte_in_6  (port_state_in_12_0_6    ), //i
    .port_byte_in_7  (port_state_in_12_0_7    ), //i
    .port_byte_out_0 (mul2_112_port_byte_out_0), //o
    .port_byte_out_1 (mul2_112_port_byte_out_1), //o
    .port_byte_out_2 (mul2_112_port_byte_out_2), //o
    .port_byte_out_3 (mul2_112_port_byte_out_3), //o
    .port_byte_out_4 (mul2_112_port_byte_out_4), //o
    .port_byte_out_5 (mul2_112_port_byte_out_5), //o
    .port_byte_out_6 (mul2_112_port_byte_out_6), //o
    .port_byte_out_7 (mul2_112_port_byte_out_7)  //o
  );
  Mul3 mul3_112 (
    .port_byte_in_0  (port_state_in_13_0_0    ), //i
    .port_byte_in_1  (port_state_in_13_0_1    ), //i
    .port_byte_in_2  (port_state_in_13_0_2    ), //i
    .port_byte_in_3  (port_state_in_13_0_3    ), //i
    .port_byte_in_4  (port_state_in_13_0_4    ), //i
    .port_byte_in_5  (port_state_in_13_0_5    ), //i
    .port_byte_in_6  (port_state_in_13_0_6    ), //i
    .port_byte_in_7  (port_state_in_13_0_7    ), //i
    .port_byte_out_0 (mul3_112_port_byte_out_0), //o
    .port_byte_out_1 (mul3_112_port_byte_out_1), //o
    .port_byte_out_2 (mul3_112_port_byte_out_2), //o
    .port_byte_out_3 (mul3_112_port_byte_out_3), //o
    .port_byte_out_4 (mul3_112_port_byte_out_4), //o
    .port_byte_out_5 (mul3_112_port_byte_out_5), //o
    .port_byte_out_6 (mul3_112_port_byte_out_6), //o
    .port_byte_out_7 (mul3_112_port_byte_out_7)  //o
  );
  Mul2 mul2_113 (
    .port_byte_in_0  (port_state_in_13_0_0    ), //i
    .port_byte_in_1  (port_state_in_13_0_1    ), //i
    .port_byte_in_2  (port_state_in_13_0_2    ), //i
    .port_byte_in_3  (port_state_in_13_0_3    ), //i
    .port_byte_in_4  (port_state_in_13_0_4    ), //i
    .port_byte_in_5  (port_state_in_13_0_5    ), //i
    .port_byte_in_6  (port_state_in_13_0_6    ), //i
    .port_byte_in_7  (port_state_in_13_0_7    ), //i
    .port_byte_out_0 (mul2_113_port_byte_out_0), //o
    .port_byte_out_1 (mul2_113_port_byte_out_1), //o
    .port_byte_out_2 (mul2_113_port_byte_out_2), //o
    .port_byte_out_3 (mul2_113_port_byte_out_3), //o
    .port_byte_out_4 (mul2_113_port_byte_out_4), //o
    .port_byte_out_5 (mul2_113_port_byte_out_5), //o
    .port_byte_out_6 (mul2_113_port_byte_out_6), //o
    .port_byte_out_7 (mul2_113_port_byte_out_7)  //o
  );
  Mul3 mul3_113 (
    .port_byte_in_0  (port_state_in_14_0_0    ), //i
    .port_byte_in_1  (port_state_in_14_0_1    ), //i
    .port_byte_in_2  (port_state_in_14_0_2    ), //i
    .port_byte_in_3  (port_state_in_14_0_3    ), //i
    .port_byte_in_4  (port_state_in_14_0_4    ), //i
    .port_byte_in_5  (port_state_in_14_0_5    ), //i
    .port_byte_in_6  (port_state_in_14_0_6    ), //i
    .port_byte_in_7  (port_state_in_14_0_7    ), //i
    .port_byte_out_0 (mul3_113_port_byte_out_0), //o
    .port_byte_out_1 (mul3_113_port_byte_out_1), //o
    .port_byte_out_2 (mul3_113_port_byte_out_2), //o
    .port_byte_out_3 (mul3_113_port_byte_out_3), //o
    .port_byte_out_4 (mul3_113_port_byte_out_4), //o
    .port_byte_out_5 (mul3_113_port_byte_out_5), //o
    .port_byte_out_6 (mul3_113_port_byte_out_6), //o
    .port_byte_out_7 (mul3_113_port_byte_out_7)  //o
  );
  Mul2 mul2_114 (
    .port_byte_in_0  (port_state_in_14_0_0    ), //i
    .port_byte_in_1  (port_state_in_14_0_1    ), //i
    .port_byte_in_2  (port_state_in_14_0_2    ), //i
    .port_byte_in_3  (port_state_in_14_0_3    ), //i
    .port_byte_in_4  (port_state_in_14_0_4    ), //i
    .port_byte_in_5  (port_state_in_14_0_5    ), //i
    .port_byte_in_6  (port_state_in_14_0_6    ), //i
    .port_byte_in_7  (port_state_in_14_0_7    ), //i
    .port_byte_out_0 (mul2_114_port_byte_out_0), //o
    .port_byte_out_1 (mul2_114_port_byte_out_1), //o
    .port_byte_out_2 (mul2_114_port_byte_out_2), //o
    .port_byte_out_3 (mul2_114_port_byte_out_3), //o
    .port_byte_out_4 (mul2_114_port_byte_out_4), //o
    .port_byte_out_5 (mul2_114_port_byte_out_5), //o
    .port_byte_out_6 (mul2_114_port_byte_out_6), //o
    .port_byte_out_7 (mul2_114_port_byte_out_7)  //o
  );
  Mul3 mul3_114 (
    .port_byte_in_0  (port_state_in_15_0_0    ), //i
    .port_byte_in_1  (port_state_in_15_0_1    ), //i
    .port_byte_in_2  (port_state_in_15_0_2    ), //i
    .port_byte_in_3  (port_state_in_15_0_3    ), //i
    .port_byte_in_4  (port_state_in_15_0_4    ), //i
    .port_byte_in_5  (port_state_in_15_0_5    ), //i
    .port_byte_in_6  (port_state_in_15_0_6    ), //i
    .port_byte_in_7  (port_state_in_15_0_7    ), //i
    .port_byte_out_0 (mul3_114_port_byte_out_0), //o
    .port_byte_out_1 (mul3_114_port_byte_out_1), //o
    .port_byte_out_2 (mul3_114_port_byte_out_2), //o
    .port_byte_out_3 (mul3_114_port_byte_out_3), //o
    .port_byte_out_4 (mul3_114_port_byte_out_4), //o
    .port_byte_out_5 (mul3_114_port_byte_out_5), //o
    .port_byte_out_6 (mul3_114_port_byte_out_6), //o
    .port_byte_out_7 (mul3_114_port_byte_out_7)  //o
  );
  Mul2 mul2_115 (
    .port_byte_in_0  (port_state_in_15_0_0    ), //i
    .port_byte_in_1  (port_state_in_15_0_1    ), //i
    .port_byte_in_2  (port_state_in_15_0_2    ), //i
    .port_byte_in_3  (port_state_in_15_0_3    ), //i
    .port_byte_in_4  (port_state_in_15_0_4    ), //i
    .port_byte_in_5  (port_state_in_15_0_5    ), //i
    .port_byte_in_6  (port_state_in_15_0_6    ), //i
    .port_byte_in_7  (port_state_in_15_0_7    ), //i
    .port_byte_out_0 (mul2_115_port_byte_out_0), //o
    .port_byte_out_1 (mul2_115_port_byte_out_1), //o
    .port_byte_out_2 (mul2_115_port_byte_out_2), //o
    .port_byte_out_3 (mul2_115_port_byte_out_3), //o
    .port_byte_out_4 (mul2_115_port_byte_out_4), //o
    .port_byte_out_5 (mul2_115_port_byte_out_5), //o
    .port_byte_out_6 (mul2_115_port_byte_out_6), //o
    .port_byte_out_7 (mul2_115_port_byte_out_7)  //o
  );
  Mul3 mul3_115 (
    .port_byte_in_0  (port_state_in_12_0_0    ), //i
    .port_byte_in_1  (port_state_in_12_0_1    ), //i
    .port_byte_in_2  (port_state_in_12_0_2    ), //i
    .port_byte_in_3  (port_state_in_12_0_3    ), //i
    .port_byte_in_4  (port_state_in_12_0_4    ), //i
    .port_byte_in_5  (port_state_in_12_0_5    ), //i
    .port_byte_in_6  (port_state_in_12_0_6    ), //i
    .port_byte_in_7  (port_state_in_12_0_7    ), //i
    .port_byte_out_0 (mul3_115_port_byte_out_0), //o
    .port_byte_out_1 (mul3_115_port_byte_out_1), //o
    .port_byte_out_2 (mul3_115_port_byte_out_2), //o
    .port_byte_out_3 (mul3_115_port_byte_out_3), //o
    .port_byte_out_4 (mul3_115_port_byte_out_4), //o
    .port_byte_out_5 (mul3_115_port_byte_out_5), //o
    .port_byte_out_6 (mul3_115_port_byte_out_6), //o
    .port_byte_out_7 (mul3_115_port_byte_out_7)  //o
  );
  Mul2 mul2_116 (
    .port_byte_in_0  (port_state_in_12_1_0    ), //i
    .port_byte_in_1  (port_state_in_12_1_1    ), //i
    .port_byte_in_2  (port_state_in_12_1_2    ), //i
    .port_byte_in_3  (port_state_in_12_1_3    ), //i
    .port_byte_in_4  (port_state_in_12_1_4    ), //i
    .port_byte_in_5  (port_state_in_12_1_5    ), //i
    .port_byte_in_6  (port_state_in_12_1_6    ), //i
    .port_byte_in_7  (port_state_in_12_1_7    ), //i
    .port_byte_out_0 (mul2_116_port_byte_out_0), //o
    .port_byte_out_1 (mul2_116_port_byte_out_1), //o
    .port_byte_out_2 (mul2_116_port_byte_out_2), //o
    .port_byte_out_3 (mul2_116_port_byte_out_3), //o
    .port_byte_out_4 (mul2_116_port_byte_out_4), //o
    .port_byte_out_5 (mul2_116_port_byte_out_5), //o
    .port_byte_out_6 (mul2_116_port_byte_out_6), //o
    .port_byte_out_7 (mul2_116_port_byte_out_7)  //o
  );
  Mul3 mul3_116 (
    .port_byte_in_0  (port_state_in_13_1_0    ), //i
    .port_byte_in_1  (port_state_in_13_1_1    ), //i
    .port_byte_in_2  (port_state_in_13_1_2    ), //i
    .port_byte_in_3  (port_state_in_13_1_3    ), //i
    .port_byte_in_4  (port_state_in_13_1_4    ), //i
    .port_byte_in_5  (port_state_in_13_1_5    ), //i
    .port_byte_in_6  (port_state_in_13_1_6    ), //i
    .port_byte_in_7  (port_state_in_13_1_7    ), //i
    .port_byte_out_0 (mul3_116_port_byte_out_0), //o
    .port_byte_out_1 (mul3_116_port_byte_out_1), //o
    .port_byte_out_2 (mul3_116_port_byte_out_2), //o
    .port_byte_out_3 (mul3_116_port_byte_out_3), //o
    .port_byte_out_4 (mul3_116_port_byte_out_4), //o
    .port_byte_out_5 (mul3_116_port_byte_out_5), //o
    .port_byte_out_6 (mul3_116_port_byte_out_6), //o
    .port_byte_out_7 (mul3_116_port_byte_out_7)  //o
  );
  Mul2 mul2_117 (
    .port_byte_in_0  (port_state_in_13_1_0    ), //i
    .port_byte_in_1  (port_state_in_13_1_1    ), //i
    .port_byte_in_2  (port_state_in_13_1_2    ), //i
    .port_byte_in_3  (port_state_in_13_1_3    ), //i
    .port_byte_in_4  (port_state_in_13_1_4    ), //i
    .port_byte_in_5  (port_state_in_13_1_5    ), //i
    .port_byte_in_6  (port_state_in_13_1_6    ), //i
    .port_byte_in_7  (port_state_in_13_1_7    ), //i
    .port_byte_out_0 (mul2_117_port_byte_out_0), //o
    .port_byte_out_1 (mul2_117_port_byte_out_1), //o
    .port_byte_out_2 (mul2_117_port_byte_out_2), //o
    .port_byte_out_3 (mul2_117_port_byte_out_3), //o
    .port_byte_out_4 (mul2_117_port_byte_out_4), //o
    .port_byte_out_5 (mul2_117_port_byte_out_5), //o
    .port_byte_out_6 (mul2_117_port_byte_out_6), //o
    .port_byte_out_7 (mul2_117_port_byte_out_7)  //o
  );
  Mul3 mul3_117 (
    .port_byte_in_0  (port_state_in_14_1_0    ), //i
    .port_byte_in_1  (port_state_in_14_1_1    ), //i
    .port_byte_in_2  (port_state_in_14_1_2    ), //i
    .port_byte_in_3  (port_state_in_14_1_3    ), //i
    .port_byte_in_4  (port_state_in_14_1_4    ), //i
    .port_byte_in_5  (port_state_in_14_1_5    ), //i
    .port_byte_in_6  (port_state_in_14_1_6    ), //i
    .port_byte_in_7  (port_state_in_14_1_7    ), //i
    .port_byte_out_0 (mul3_117_port_byte_out_0), //o
    .port_byte_out_1 (mul3_117_port_byte_out_1), //o
    .port_byte_out_2 (mul3_117_port_byte_out_2), //o
    .port_byte_out_3 (mul3_117_port_byte_out_3), //o
    .port_byte_out_4 (mul3_117_port_byte_out_4), //o
    .port_byte_out_5 (mul3_117_port_byte_out_5), //o
    .port_byte_out_6 (mul3_117_port_byte_out_6), //o
    .port_byte_out_7 (mul3_117_port_byte_out_7)  //o
  );
  Mul2 mul2_118 (
    .port_byte_in_0  (port_state_in_14_1_0    ), //i
    .port_byte_in_1  (port_state_in_14_1_1    ), //i
    .port_byte_in_2  (port_state_in_14_1_2    ), //i
    .port_byte_in_3  (port_state_in_14_1_3    ), //i
    .port_byte_in_4  (port_state_in_14_1_4    ), //i
    .port_byte_in_5  (port_state_in_14_1_5    ), //i
    .port_byte_in_6  (port_state_in_14_1_6    ), //i
    .port_byte_in_7  (port_state_in_14_1_7    ), //i
    .port_byte_out_0 (mul2_118_port_byte_out_0), //o
    .port_byte_out_1 (mul2_118_port_byte_out_1), //o
    .port_byte_out_2 (mul2_118_port_byte_out_2), //o
    .port_byte_out_3 (mul2_118_port_byte_out_3), //o
    .port_byte_out_4 (mul2_118_port_byte_out_4), //o
    .port_byte_out_5 (mul2_118_port_byte_out_5), //o
    .port_byte_out_6 (mul2_118_port_byte_out_6), //o
    .port_byte_out_7 (mul2_118_port_byte_out_7)  //o
  );
  Mul3 mul3_118 (
    .port_byte_in_0  (port_state_in_15_1_0    ), //i
    .port_byte_in_1  (port_state_in_15_1_1    ), //i
    .port_byte_in_2  (port_state_in_15_1_2    ), //i
    .port_byte_in_3  (port_state_in_15_1_3    ), //i
    .port_byte_in_4  (port_state_in_15_1_4    ), //i
    .port_byte_in_5  (port_state_in_15_1_5    ), //i
    .port_byte_in_6  (port_state_in_15_1_6    ), //i
    .port_byte_in_7  (port_state_in_15_1_7    ), //i
    .port_byte_out_0 (mul3_118_port_byte_out_0), //o
    .port_byte_out_1 (mul3_118_port_byte_out_1), //o
    .port_byte_out_2 (mul3_118_port_byte_out_2), //o
    .port_byte_out_3 (mul3_118_port_byte_out_3), //o
    .port_byte_out_4 (mul3_118_port_byte_out_4), //o
    .port_byte_out_5 (mul3_118_port_byte_out_5), //o
    .port_byte_out_6 (mul3_118_port_byte_out_6), //o
    .port_byte_out_7 (mul3_118_port_byte_out_7)  //o
  );
  Mul2 mul2_119 (
    .port_byte_in_0  (port_state_in_15_1_0    ), //i
    .port_byte_in_1  (port_state_in_15_1_1    ), //i
    .port_byte_in_2  (port_state_in_15_1_2    ), //i
    .port_byte_in_3  (port_state_in_15_1_3    ), //i
    .port_byte_in_4  (port_state_in_15_1_4    ), //i
    .port_byte_in_5  (port_state_in_15_1_5    ), //i
    .port_byte_in_6  (port_state_in_15_1_6    ), //i
    .port_byte_in_7  (port_state_in_15_1_7    ), //i
    .port_byte_out_0 (mul2_119_port_byte_out_0), //o
    .port_byte_out_1 (mul2_119_port_byte_out_1), //o
    .port_byte_out_2 (mul2_119_port_byte_out_2), //o
    .port_byte_out_3 (mul2_119_port_byte_out_3), //o
    .port_byte_out_4 (mul2_119_port_byte_out_4), //o
    .port_byte_out_5 (mul2_119_port_byte_out_5), //o
    .port_byte_out_6 (mul2_119_port_byte_out_6), //o
    .port_byte_out_7 (mul2_119_port_byte_out_7)  //o
  );
  Mul3 mul3_119 (
    .port_byte_in_0  (port_state_in_12_1_0    ), //i
    .port_byte_in_1  (port_state_in_12_1_1    ), //i
    .port_byte_in_2  (port_state_in_12_1_2    ), //i
    .port_byte_in_3  (port_state_in_12_1_3    ), //i
    .port_byte_in_4  (port_state_in_12_1_4    ), //i
    .port_byte_in_5  (port_state_in_12_1_5    ), //i
    .port_byte_in_6  (port_state_in_12_1_6    ), //i
    .port_byte_in_7  (port_state_in_12_1_7    ), //i
    .port_byte_out_0 (mul3_119_port_byte_out_0), //o
    .port_byte_out_1 (mul3_119_port_byte_out_1), //o
    .port_byte_out_2 (mul3_119_port_byte_out_2), //o
    .port_byte_out_3 (mul3_119_port_byte_out_3), //o
    .port_byte_out_4 (mul3_119_port_byte_out_4), //o
    .port_byte_out_5 (mul3_119_port_byte_out_5), //o
    .port_byte_out_6 (mul3_119_port_byte_out_6), //o
    .port_byte_out_7 (mul3_119_port_byte_out_7)  //o
  );
  Mul2 mul2_120 (
    .port_byte_in_0  (port_state_in_12_2_0    ), //i
    .port_byte_in_1  (port_state_in_12_2_1    ), //i
    .port_byte_in_2  (port_state_in_12_2_2    ), //i
    .port_byte_in_3  (port_state_in_12_2_3    ), //i
    .port_byte_in_4  (port_state_in_12_2_4    ), //i
    .port_byte_in_5  (port_state_in_12_2_5    ), //i
    .port_byte_in_6  (port_state_in_12_2_6    ), //i
    .port_byte_in_7  (port_state_in_12_2_7    ), //i
    .port_byte_out_0 (mul2_120_port_byte_out_0), //o
    .port_byte_out_1 (mul2_120_port_byte_out_1), //o
    .port_byte_out_2 (mul2_120_port_byte_out_2), //o
    .port_byte_out_3 (mul2_120_port_byte_out_3), //o
    .port_byte_out_4 (mul2_120_port_byte_out_4), //o
    .port_byte_out_5 (mul2_120_port_byte_out_5), //o
    .port_byte_out_6 (mul2_120_port_byte_out_6), //o
    .port_byte_out_7 (mul2_120_port_byte_out_7)  //o
  );
  Mul3 mul3_120 (
    .port_byte_in_0  (port_state_in_13_2_0    ), //i
    .port_byte_in_1  (port_state_in_13_2_1    ), //i
    .port_byte_in_2  (port_state_in_13_2_2    ), //i
    .port_byte_in_3  (port_state_in_13_2_3    ), //i
    .port_byte_in_4  (port_state_in_13_2_4    ), //i
    .port_byte_in_5  (port_state_in_13_2_5    ), //i
    .port_byte_in_6  (port_state_in_13_2_6    ), //i
    .port_byte_in_7  (port_state_in_13_2_7    ), //i
    .port_byte_out_0 (mul3_120_port_byte_out_0), //o
    .port_byte_out_1 (mul3_120_port_byte_out_1), //o
    .port_byte_out_2 (mul3_120_port_byte_out_2), //o
    .port_byte_out_3 (mul3_120_port_byte_out_3), //o
    .port_byte_out_4 (mul3_120_port_byte_out_4), //o
    .port_byte_out_5 (mul3_120_port_byte_out_5), //o
    .port_byte_out_6 (mul3_120_port_byte_out_6), //o
    .port_byte_out_7 (mul3_120_port_byte_out_7)  //o
  );
  Mul2 mul2_121 (
    .port_byte_in_0  (port_state_in_13_2_0    ), //i
    .port_byte_in_1  (port_state_in_13_2_1    ), //i
    .port_byte_in_2  (port_state_in_13_2_2    ), //i
    .port_byte_in_3  (port_state_in_13_2_3    ), //i
    .port_byte_in_4  (port_state_in_13_2_4    ), //i
    .port_byte_in_5  (port_state_in_13_2_5    ), //i
    .port_byte_in_6  (port_state_in_13_2_6    ), //i
    .port_byte_in_7  (port_state_in_13_2_7    ), //i
    .port_byte_out_0 (mul2_121_port_byte_out_0), //o
    .port_byte_out_1 (mul2_121_port_byte_out_1), //o
    .port_byte_out_2 (mul2_121_port_byte_out_2), //o
    .port_byte_out_3 (mul2_121_port_byte_out_3), //o
    .port_byte_out_4 (mul2_121_port_byte_out_4), //o
    .port_byte_out_5 (mul2_121_port_byte_out_5), //o
    .port_byte_out_6 (mul2_121_port_byte_out_6), //o
    .port_byte_out_7 (mul2_121_port_byte_out_7)  //o
  );
  Mul3 mul3_121 (
    .port_byte_in_0  (port_state_in_14_2_0    ), //i
    .port_byte_in_1  (port_state_in_14_2_1    ), //i
    .port_byte_in_2  (port_state_in_14_2_2    ), //i
    .port_byte_in_3  (port_state_in_14_2_3    ), //i
    .port_byte_in_4  (port_state_in_14_2_4    ), //i
    .port_byte_in_5  (port_state_in_14_2_5    ), //i
    .port_byte_in_6  (port_state_in_14_2_6    ), //i
    .port_byte_in_7  (port_state_in_14_2_7    ), //i
    .port_byte_out_0 (mul3_121_port_byte_out_0), //o
    .port_byte_out_1 (mul3_121_port_byte_out_1), //o
    .port_byte_out_2 (mul3_121_port_byte_out_2), //o
    .port_byte_out_3 (mul3_121_port_byte_out_3), //o
    .port_byte_out_4 (mul3_121_port_byte_out_4), //o
    .port_byte_out_5 (mul3_121_port_byte_out_5), //o
    .port_byte_out_6 (mul3_121_port_byte_out_6), //o
    .port_byte_out_7 (mul3_121_port_byte_out_7)  //o
  );
  Mul2 mul2_122 (
    .port_byte_in_0  (port_state_in_14_2_0    ), //i
    .port_byte_in_1  (port_state_in_14_2_1    ), //i
    .port_byte_in_2  (port_state_in_14_2_2    ), //i
    .port_byte_in_3  (port_state_in_14_2_3    ), //i
    .port_byte_in_4  (port_state_in_14_2_4    ), //i
    .port_byte_in_5  (port_state_in_14_2_5    ), //i
    .port_byte_in_6  (port_state_in_14_2_6    ), //i
    .port_byte_in_7  (port_state_in_14_2_7    ), //i
    .port_byte_out_0 (mul2_122_port_byte_out_0), //o
    .port_byte_out_1 (mul2_122_port_byte_out_1), //o
    .port_byte_out_2 (mul2_122_port_byte_out_2), //o
    .port_byte_out_3 (mul2_122_port_byte_out_3), //o
    .port_byte_out_4 (mul2_122_port_byte_out_4), //o
    .port_byte_out_5 (mul2_122_port_byte_out_5), //o
    .port_byte_out_6 (mul2_122_port_byte_out_6), //o
    .port_byte_out_7 (mul2_122_port_byte_out_7)  //o
  );
  Mul3 mul3_122 (
    .port_byte_in_0  (port_state_in_15_2_0    ), //i
    .port_byte_in_1  (port_state_in_15_2_1    ), //i
    .port_byte_in_2  (port_state_in_15_2_2    ), //i
    .port_byte_in_3  (port_state_in_15_2_3    ), //i
    .port_byte_in_4  (port_state_in_15_2_4    ), //i
    .port_byte_in_5  (port_state_in_15_2_5    ), //i
    .port_byte_in_6  (port_state_in_15_2_6    ), //i
    .port_byte_in_7  (port_state_in_15_2_7    ), //i
    .port_byte_out_0 (mul3_122_port_byte_out_0), //o
    .port_byte_out_1 (mul3_122_port_byte_out_1), //o
    .port_byte_out_2 (mul3_122_port_byte_out_2), //o
    .port_byte_out_3 (mul3_122_port_byte_out_3), //o
    .port_byte_out_4 (mul3_122_port_byte_out_4), //o
    .port_byte_out_5 (mul3_122_port_byte_out_5), //o
    .port_byte_out_6 (mul3_122_port_byte_out_6), //o
    .port_byte_out_7 (mul3_122_port_byte_out_7)  //o
  );
  Mul2 mul2_123 (
    .port_byte_in_0  (port_state_in_15_2_0    ), //i
    .port_byte_in_1  (port_state_in_15_2_1    ), //i
    .port_byte_in_2  (port_state_in_15_2_2    ), //i
    .port_byte_in_3  (port_state_in_15_2_3    ), //i
    .port_byte_in_4  (port_state_in_15_2_4    ), //i
    .port_byte_in_5  (port_state_in_15_2_5    ), //i
    .port_byte_in_6  (port_state_in_15_2_6    ), //i
    .port_byte_in_7  (port_state_in_15_2_7    ), //i
    .port_byte_out_0 (mul2_123_port_byte_out_0), //o
    .port_byte_out_1 (mul2_123_port_byte_out_1), //o
    .port_byte_out_2 (mul2_123_port_byte_out_2), //o
    .port_byte_out_3 (mul2_123_port_byte_out_3), //o
    .port_byte_out_4 (mul2_123_port_byte_out_4), //o
    .port_byte_out_5 (mul2_123_port_byte_out_5), //o
    .port_byte_out_6 (mul2_123_port_byte_out_6), //o
    .port_byte_out_7 (mul2_123_port_byte_out_7)  //o
  );
  Mul3 mul3_123 (
    .port_byte_in_0  (port_state_in_12_2_0    ), //i
    .port_byte_in_1  (port_state_in_12_2_1    ), //i
    .port_byte_in_2  (port_state_in_12_2_2    ), //i
    .port_byte_in_3  (port_state_in_12_2_3    ), //i
    .port_byte_in_4  (port_state_in_12_2_4    ), //i
    .port_byte_in_5  (port_state_in_12_2_5    ), //i
    .port_byte_in_6  (port_state_in_12_2_6    ), //i
    .port_byte_in_7  (port_state_in_12_2_7    ), //i
    .port_byte_out_0 (mul3_123_port_byte_out_0), //o
    .port_byte_out_1 (mul3_123_port_byte_out_1), //o
    .port_byte_out_2 (mul3_123_port_byte_out_2), //o
    .port_byte_out_3 (mul3_123_port_byte_out_3), //o
    .port_byte_out_4 (mul3_123_port_byte_out_4), //o
    .port_byte_out_5 (mul3_123_port_byte_out_5), //o
    .port_byte_out_6 (mul3_123_port_byte_out_6), //o
    .port_byte_out_7 (mul3_123_port_byte_out_7)  //o
  );
  Mul2 mul2_124 (
    .port_byte_in_0  (port_state_in_12_3_0    ), //i
    .port_byte_in_1  (port_state_in_12_3_1    ), //i
    .port_byte_in_2  (port_state_in_12_3_2    ), //i
    .port_byte_in_3  (port_state_in_12_3_3    ), //i
    .port_byte_in_4  (port_state_in_12_3_4    ), //i
    .port_byte_in_5  (port_state_in_12_3_5    ), //i
    .port_byte_in_6  (port_state_in_12_3_6    ), //i
    .port_byte_in_7  (port_state_in_12_3_7    ), //i
    .port_byte_out_0 (mul2_124_port_byte_out_0), //o
    .port_byte_out_1 (mul2_124_port_byte_out_1), //o
    .port_byte_out_2 (mul2_124_port_byte_out_2), //o
    .port_byte_out_3 (mul2_124_port_byte_out_3), //o
    .port_byte_out_4 (mul2_124_port_byte_out_4), //o
    .port_byte_out_5 (mul2_124_port_byte_out_5), //o
    .port_byte_out_6 (mul2_124_port_byte_out_6), //o
    .port_byte_out_7 (mul2_124_port_byte_out_7)  //o
  );
  Mul3 mul3_124 (
    .port_byte_in_0  (port_state_in_13_3_0    ), //i
    .port_byte_in_1  (port_state_in_13_3_1    ), //i
    .port_byte_in_2  (port_state_in_13_3_2    ), //i
    .port_byte_in_3  (port_state_in_13_3_3    ), //i
    .port_byte_in_4  (port_state_in_13_3_4    ), //i
    .port_byte_in_5  (port_state_in_13_3_5    ), //i
    .port_byte_in_6  (port_state_in_13_3_6    ), //i
    .port_byte_in_7  (port_state_in_13_3_7    ), //i
    .port_byte_out_0 (mul3_124_port_byte_out_0), //o
    .port_byte_out_1 (mul3_124_port_byte_out_1), //o
    .port_byte_out_2 (mul3_124_port_byte_out_2), //o
    .port_byte_out_3 (mul3_124_port_byte_out_3), //o
    .port_byte_out_4 (mul3_124_port_byte_out_4), //o
    .port_byte_out_5 (mul3_124_port_byte_out_5), //o
    .port_byte_out_6 (mul3_124_port_byte_out_6), //o
    .port_byte_out_7 (mul3_124_port_byte_out_7)  //o
  );
  Mul2 mul2_125 (
    .port_byte_in_0  (port_state_in_13_3_0    ), //i
    .port_byte_in_1  (port_state_in_13_3_1    ), //i
    .port_byte_in_2  (port_state_in_13_3_2    ), //i
    .port_byte_in_3  (port_state_in_13_3_3    ), //i
    .port_byte_in_4  (port_state_in_13_3_4    ), //i
    .port_byte_in_5  (port_state_in_13_3_5    ), //i
    .port_byte_in_6  (port_state_in_13_3_6    ), //i
    .port_byte_in_7  (port_state_in_13_3_7    ), //i
    .port_byte_out_0 (mul2_125_port_byte_out_0), //o
    .port_byte_out_1 (mul2_125_port_byte_out_1), //o
    .port_byte_out_2 (mul2_125_port_byte_out_2), //o
    .port_byte_out_3 (mul2_125_port_byte_out_3), //o
    .port_byte_out_4 (mul2_125_port_byte_out_4), //o
    .port_byte_out_5 (mul2_125_port_byte_out_5), //o
    .port_byte_out_6 (mul2_125_port_byte_out_6), //o
    .port_byte_out_7 (mul2_125_port_byte_out_7)  //o
  );
  Mul3 mul3_125 (
    .port_byte_in_0  (port_state_in_14_3_0    ), //i
    .port_byte_in_1  (port_state_in_14_3_1    ), //i
    .port_byte_in_2  (port_state_in_14_3_2    ), //i
    .port_byte_in_3  (port_state_in_14_3_3    ), //i
    .port_byte_in_4  (port_state_in_14_3_4    ), //i
    .port_byte_in_5  (port_state_in_14_3_5    ), //i
    .port_byte_in_6  (port_state_in_14_3_6    ), //i
    .port_byte_in_7  (port_state_in_14_3_7    ), //i
    .port_byte_out_0 (mul3_125_port_byte_out_0), //o
    .port_byte_out_1 (mul3_125_port_byte_out_1), //o
    .port_byte_out_2 (mul3_125_port_byte_out_2), //o
    .port_byte_out_3 (mul3_125_port_byte_out_3), //o
    .port_byte_out_4 (mul3_125_port_byte_out_4), //o
    .port_byte_out_5 (mul3_125_port_byte_out_5), //o
    .port_byte_out_6 (mul3_125_port_byte_out_6), //o
    .port_byte_out_7 (mul3_125_port_byte_out_7)  //o
  );
  Mul2 mul2_126 (
    .port_byte_in_0  (port_state_in_14_3_0    ), //i
    .port_byte_in_1  (port_state_in_14_3_1    ), //i
    .port_byte_in_2  (port_state_in_14_3_2    ), //i
    .port_byte_in_3  (port_state_in_14_3_3    ), //i
    .port_byte_in_4  (port_state_in_14_3_4    ), //i
    .port_byte_in_5  (port_state_in_14_3_5    ), //i
    .port_byte_in_6  (port_state_in_14_3_6    ), //i
    .port_byte_in_7  (port_state_in_14_3_7    ), //i
    .port_byte_out_0 (mul2_126_port_byte_out_0), //o
    .port_byte_out_1 (mul2_126_port_byte_out_1), //o
    .port_byte_out_2 (mul2_126_port_byte_out_2), //o
    .port_byte_out_3 (mul2_126_port_byte_out_3), //o
    .port_byte_out_4 (mul2_126_port_byte_out_4), //o
    .port_byte_out_5 (mul2_126_port_byte_out_5), //o
    .port_byte_out_6 (mul2_126_port_byte_out_6), //o
    .port_byte_out_7 (mul2_126_port_byte_out_7)  //o
  );
  Mul3 mul3_126 (
    .port_byte_in_0  (port_state_in_15_3_0    ), //i
    .port_byte_in_1  (port_state_in_15_3_1    ), //i
    .port_byte_in_2  (port_state_in_15_3_2    ), //i
    .port_byte_in_3  (port_state_in_15_3_3    ), //i
    .port_byte_in_4  (port_state_in_15_3_4    ), //i
    .port_byte_in_5  (port_state_in_15_3_5    ), //i
    .port_byte_in_6  (port_state_in_15_3_6    ), //i
    .port_byte_in_7  (port_state_in_15_3_7    ), //i
    .port_byte_out_0 (mul3_126_port_byte_out_0), //o
    .port_byte_out_1 (mul3_126_port_byte_out_1), //o
    .port_byte_out_2 (mul3_126_port_byte_out_2), //o
    .port_byte_out_3 (mul3_126_port_byte_out_3), //o
    .port_byte_out_4 (mul3_126_port_byte_out_4), //o
    .port_byte_out_5 (mul3_126_port_byte_out_5), //o
    .port_byte_out_6 (mul3_126_port_byte_out_6), //o
    .port_byte_out_7 (mul3_126_port_byte_out_7)  //o
  );
  Mul2 mul2_127 (
    .port_byte_in_0  (port_state_in_15_3_0    ), //i
    .port_byte_in_1  (port_state_in_15_3_1    ), //i
    .port_byte_in_2  (port_state_in_15_3_2    ), //i
    .port_byte_in_3  (port_state_in_15_3_3    ), //i
    .port_byte_in_4  (port_state_in_15_3_4    ), //i
    .port_byte_in_5  (port_state_in_15_3_5    ), //i
    .port_byte_in_6  (port_state_in_15_3_6    ), //i
    .port_byte_in_7  (port_state_in_15_3_7    ), //i
    .port_byte_out_0 (mul2_127_port_byte_out_0), //o
    .port_byte_out_1 (mul2_127_port_byte_out_1), //o
    .port_byte_out_2 (mul2_127_port_byte_out_2), //o
    .port_byte_out_3 (mul2_127_port_byte_out_3), //o
    .port_byte_out_4 (mul2_127_port_byte_out_4), //o
    .port_byte_out_5 (mul2_127_port_byte_out_5), //o
    .port_byte_out_6 (mul2_127_port_byte_out_6), //o
    .port_byte_out_7 (mul2_127_port_byte_out_7)  //o
  );
  Mul3 mul3_127 (
    .port_byte_in_0  (port_state_in_12_3_0    ), //i
    .port_byte_in_1  (port_state_in_12_3_1    ), //i
    .port_byte_in_2  (port_state_in_12_3_2    ), //i
    .port_byte_in_3  (port_state_in_12_3_3    ), //i
    .port_byte_in_4  (port_state_in_12_3_4    ), //i
    .port_byte_in_5  (port_state_in_12_3_5    ), //i
    .port_byte_in_6  (port_state_in_12_3_6    ), //i
    .port_byte_in_7  (port_state_in_12_3_7    ), //i
    .port_byte_out_0 (mul3_127_port_byte_out_0), //o
    .port_byte_out_1 (mul3_127_port_byte_out_1), //o
    .port_byte_out_2 (mul3_127_port_byte_out_2), //o
    .port_byte_out_3 (mul3_127_port_byte_out_3), //o
    .port_byte_out_4 (mul3_127_port_byte_out_4), //o
    .port_byte_out_5 (mul3_127_port_byte_out_5), //o
    .port_byte_out_6 (mul3_127_port_byte_out_6), //o
    .port_byte_out_7 (mul3_127_port_byte_out_7)  //o
  );
  assign state_out_0_0_0 = (((mul2_64_port_byte_out_0 ^ mul3_64_port_byte_out_0) ^ port_state_in_2_0_0) ^ port_state_in_3_0_0);
  assign state_out_1_0_0 = (((mul2_65_port_byte_out_0 ^ mul3_65_port_byte_out_0) ^ port_state_in_0_0_0) ^ port_state_in_3_0_0);
  assign state_out_2_0_0 = (((mul2_66_port_byte_out_0 ^ mul3_66_port_byte_out_0) ^ port_state_in_0_0_0) ^ port_state_in_1_0_0);
  assign state_out_3_0_0 = (((mul2_67_port_byte_out_0 ^ mul3_67_port_byte_out_0) ^ port_state_in_1_0_0) ^ port_state_in_2_0_0);
  assign state_out_0_0_1 = (((mul2_64_port_byte_out_1 ^ mul3_64_port_byte_out_1) ^ port_state_in_2_0_1) ^ port_state_in_3_0_1);
  assign state_out_1_0_1 = (((mul2_65_port_byte_out_1 ^ mul3_65_port_byte_out_1) ^ port_state_in_0_0_1) ^ port_state_in_3_0_1);
  assign state_out_2_0_1 = (((mul2_66_port_byte_out_1 ^ mul3_66_port_byte_out_1) ^ port_state_in_0_0_1) ^ port_state_in_1_0_1);
  assign state_out_3_0_1 = (((mul2_67_port_byte_out_1 ^ mul3_67_port_byte_out_1) ^ port_state_in_1_0_1) ^ port_state_in_2_0_1);
  assign state_out_0_0_2 = (((mul2_64_port_byte_out_2 ^ mul3_64_port_byte_out_2) ^ port_state_in_2_0_2) ^ port_state_in_3_0_2);
  assign state_out_1_0_2 = (((mul2_65_port_byte_out_2 ^ mul3_65_port_byte_out_2) ^ port_state_in_0_0_2) ^ port_state_in_3_0_2);
  assign state_out_2_0_2 = (((mul2_66_port_byte_out_2 ^ mul3_66_port_byte_out_2) ^ port_state_in_0_0_2) ^ port_state_in_1_0_2);
  assign state_out_3_0_2 = (((mul2_67_port_byte_out_2 ^ mul3_67_port_byte_out_2) ^ port_state_in_1_0_2) ^ port_state_in_2_0_2);
  assign state_out_0_0_3 = (((mul2_64_port_byte_out_3 ^ mul3_64_port_byte_out_3) ^ port_state_in_2_0_3) ^ port_state_in_3_0_3);
  assign state_out_1_0_3 = (((mul2_65_port_byte_out_3 ^ mul3_65_port_byte_out_3) ^ port_state_in_0_0_3) ^ port_state_in_3_0_3);
  assign state_out_2_0_3 = (((mul2_66_port_byte_out_3 ^ mul3_66_port_byte_out_3) ^ port_state_in_0_0_3) ^ port_state_in_1_0_3);
  assign state_out_3_0_3 = (((mul2_67_port_byte_out_3 ^ mul3_67_port_byte_out_3) ^ port_state_in_1_0_3) ^ port_state_in_2_0_3);
  assign state_out_0_0_4 = (((mul2_64_port_byte_out_4 ^ mul3_64_port_byte_out_4) ^ port_state_in_2_0_4) ^ port_state_in_3_0_4);
  assign state_out_1_0_4 = (((mul2_65_port_byte_out_4 ^ mul3_65_port_byte_out_4) ^ port_state_in_0_0_4) ^ port_state_in_3_0_4);
  assign state_out_2_0_4 = (((mul2_66_port_byte_out_4 ^ mul3_66_port_byte_out_4) ^ port_state_in_0_0_4) ^ port_state_in_1_0_4);
  assign state_out_3_0_4 = (((mul2_67_port_byte_out_4 ^ mul3_67_port_byte_out_4) ^ port_state_in_1_0_4) ^ port_state_in_2_0_4);
  assign state_out_0_0_5 = (((mul2_64_port_byte_out_5 ^ mul3_64_port_byte_out_5) ^ port_state_in_2_0_5) ^ port_state_in_3_0_5);
  assign state_out_1_0_5 = (((mul2_65_port_byte_out_5 ^ mul3_65_port_byte_out_5) ^ port_state_in_0_0_5) ^ port_state_in_3_0_5);
  assign state_out_2_0_5 = (((mul2_66_port_byte_out_5 ^ mul3_66_port_byte_out_5) ^ port_state_in_0_0_5) ^ port_state_in_1_0_5);
  assign state_out_3_0_5 = (((mul2_67_port_byte_out_5 ^ mul3_67_port_byte_out_5) ^ port_state_in_1_0_5) ^ port_state_in_2_0_5);
  assign state_out_0_0_6 = (((mul2_64_port_byte_out_6 ^ mul3_64_port_byte_out_6) ^ port_state_in_2_0_6) ^ port_state_in_3_0_6);
  assign state_out_1_0_6 = (((mul2_65_port_byte_out_6 ^ mul3_65_port_byte_out_6) ^ port_state_in_0_0_6) ^ port_state_in_3_0_6);
  assign state_out_2_0_6 = (((mul2_66_port_byte_out_6 ^ mul3_66_port_byte_out_6) ^ port_state_in_0_0_6) ^ port_state_in_1_0_6);
  assign state_out_3_0_6 = (((mul2_67_port_byte_out_6 ^ mul3_67_port_byte_out_6) ^ port_state_in_1_0_6) ^ port_state_in_2_0_6);
  assign state_out_0_0_7 = (((mul2_64_port_byte_out_7 ^ mul3_64_port_byte_out_7) ^ port_state_in_2_0_7) ^ port_state_in_3_0_7);
  assign state_out_1_0_7 = (((mul2_65_port_byte_out_7 ^ mul3_65_port_byte_out_7) ^ port_state_in_0_0_7) ^ port_state_in_3_0_7);
  assign state_out_2_0_7 = (((mul2_66_port_byte_out_7 ^ mul3_66_port_byte_out_7) ^ port_state_in_0_0_7) ^ port_state_in_1_0_7);
  assign state_out_3_0_7 = (((mul2_67_port_byte_out_7 ^ mul3_67_port_byte_out_7) ^ port_state_in_1_0_7) ^ port_state_in_2_0_7);
  assign state_out_0_1_0 = (((mul2_68_port_byte_out_0 ^ mul3_68_port_byte_out_0) ^ port_state_in_2_1_0) ^ port_state_in_3_1_0);
  assign state_out_1_1_0 = (((mul2_69_port_byte_out_0 ^ mul3_69_port_byte_out_0) ^ port_state_in_0_1_0) ^ port_state_in_3_1_0);
  assign state_out_2_1_0 = (((mul2_70_port_byte_out_0 ^ mul3_70_port_byte_out_0) ^ port_state_in_0_1_0) ^ port_state_in_1_1_0);
  assign state_out_3_1_0 = (((mul2_71_port_byte_out_0 ^ mul3_71_port_byte_out_0) ^ port_state_in_1_1_0) ^ port_state_in_2_1_0);
  assign state_out_0_1_1 = (((mul2_68_port_byte_out_1 ^ mul3_68_port_byte_out_1) ^ port_state_in_2_1_1) ^ port_state_in_3_1_1);
  assign state_out_1_1_1 = (((mul2_69_port_byte_out_1 ^ mul3_69_port_byte_out_1) ^ port_state_in_0_1_1) ^ port_state_in_3_1_1);
  assign state_out_2_1_1 = (((mul2_70_port_byte_out_1 ^ mul3_70_port_byte_out_1) ^ port_state_in_0_1_1) ^ port_state_in_1_1_1);
  assign state_out_3_1_1 = (((mul2_71_port_byte_out_1 ^ mul3_71_port_byte_out_1) ^ port_state_in_1_1_1) ^ port_state_in_2_1_1);
  assign state_out_0_1_2 = (((mul2_68_port_byte_out_2 ^ mul3_68_port_byte_out_2) ^ port_state_in_2_1_2) ^ port_state_in_3_1_2);
  assign state_out_1_1_2 = (((mul2_69_port_byte_out_2 ^ mul3_69_port_byte_out_2) ^ port_state_in_0_1_2) ^ port_state_in_3_1_2);
  assign state_out_2_1_2 = (((mul2_70_port_byte_out_2 ^ mul3_70_port_byte_out_2) ^ port_state_in_0_1_2) ^ port_state_in_1_1_2);
  assign state_out_3_1_2 = (((mul2_71_port_byte_out_2 ^ mul3_71_port_byte_out_2) ^ port_state_in_1_1_2) ^ port_state_in_2_1_2);
  assign state_out_0_1_3 = (((mul2_68_port_byte_out_3 ^ mul3_68_port_byte_out_3) ^ port_state_in_2_1_3) ^ port_state_in_3_1_3);
  assign state_out_1_1_3 = (((mul2_69_port_byte_out_3 ^ mul3_69_port_byte_out_3) ^ port_state_in_0_1_3) ^ port_state_in_3_1_3);
  assign state_out_2_1_3 = (((mul2_70_port_byte_out_3 ^ mul3_70_port_byte_out_3) ^ port_state_in_0_1_3) ^ port_state_in_1_1_3);
  assign state_out_3_1_3 = (((mul2_71_port_byte_out_3 ^ mul3_71_port_byte_out_3) ^ port_state_in_1_1_3) ^ port_state_in_2_1_3);
  assign state_out_0_1_4 = (((mul2_68_port_byte_out_4 ^ mul3_68_port_byte_out_4) ^ port_state_in_2_1_4) ^ port_state_in_3_1_4);
  assign state_out_1_1_4 = (((mul2_69_port_byte_out_4 ^ mul3_69_port_byte_out_4) ^ port_state_in_0_1_4) ^ port_state_in_3_1_4);
  assign state_out_2_1_4 = (((mul2_70_port_byte_out_4 ^ mul3_70_port_byte_out_4) ^ port_state_in_0_1_4) ^ port_state_in_1_1_4);
  assign state_out_3_1_4 = (((mul2_71_port_byte_out_4 ^ mul3_71_port_byte_out_4) ^ port_state_in_1_1_4) ^ port_state_in_2_1_4);
  assign state_out_0_1_5 = (((mul2_68_port_byte_out_5 ^ mul3_68_port_byte_out_5) ^ port_state_in_2_1_5) ^ port_state_in_3_1_5);
  assign state_out_1_1_5 = (((mul2_69_port_byte_out_5 ^ mul3_69_port_byte_out_5) ^ port_state_in_0_1_5) ^ port_state_in_3_1_5);
  assign state_out_2_1_5 = (((mul2_70_port_byte_out_5 ^ mul3_70_port_byte_out_5) ^ port_state_in_0_1_5) ^ port_state_in_1_1_5);
  assign state_out_3_1_5 = (((mul2_71_port_byte_out_5 ^ mul3_71_port_byte_out_5) ^ port_state_in_1_1_5) ^ port_state_in_2_1_5);
  assign state_out_0_1_6 = (((mul2_68_port_byte_out_6 ^ mul3_68_port_byte_out_6) ^ port_state_in_2_1_6) ^ port_state_in_3_1_6);
  assign state_out_1_1_6 = (((mul2_69_port_byte_out_6 ^ mul3_69_port_byte_out_6) ^ port_state_in_0_1_6) ^ port_state_in_3_1_6);
  assign state_out_2_1_6 = (((mul2_70_port_byte_out_6 ^ mul3_70_port_byte_out_6) ^ port_state_in_0_1_6) ^ port_state_in_1_1_6);
  assign state_out_3_1_6 = (((mul2_71_port_byte_out_6 ^ mul3_71_port_byte_out_6) ^ port_state_in_1_1_6) ^ port_state_in_2_1_6);
  assign state_out_0_1_7 = (((mul2_68_port_byte_out_7 ^ mul3_68_port_byte_out_7) ^ port_state_in_2_1_7) ^ port_state_in_3_1_7);
  assign state_out_1_1_7 = (((mul2_69_port_byte_out_7 ^ mul3_69_port_byte_out_7) ^ port_state_in_0_1_7) ^ port_state_in_3_1_7);
  assign state_out_2_1_7 = (((mul2_70_port_byte_out_7 ^ mul3_70_port_byte_out_7) ^ port_state_in_0_1_7) ^ port_state_in_1_1_7);
  assign state_out_3_1_7 = (((mul2_71_port_byte_out_7 ^ mul3_71_port_byte_out_7) ^ port_state_in_1_1_7) ^ port_state_in_2_1_7);
  assign state_out_0_2_0 = (((mul2_72_port_byte_out_0 ^ mul3_72_port_byte_out_0) ^ port_state_in_2_2_0) ^ port_state_in_3_2_0);
  assign state_out_1_2_0 = (((mul2_73_port_byte_out_0 ^ mul3_73_port_byte_out_0) ^ port_state_in_0_2_0) ^ port_state_in_3_2_0);
  assign state_out_2_2_0 = (((mul2_74_port_byte_out_0 ^ mul3_74_port_byte_out_0) ^ port_state_in_0_2_0) ^ port_state_in_1_2_0);
  assign state_out_3_2_0 = (((mul2_75_port_byte_out_0 ^ mul3_75_port_byte_out_0) ^ port_state_in_1_2_0) ^ port_state_in_2_2_0);
  assign state_out_0_2_1 = (((mul2_72_port_byte_out_1 ^ mul3_72_port_byte_out_1) ^ port_state_in_2_2_1) ^ port_state_in_3_2_1);
  assign state_out_1_2_1 = (((mul2_73_port_byte_out_1 ^ mul3_73_port_byte_out_1) ^ port_state_in_0_2_1) ^ port_state_in_3_2_1);
  assign state_out_2_2_1 = (((mul2_74_port_byte_out_1 ^ mul3_74_port_byte_out_1) ^ port_state_in_0_2_1) ^ port_state_in_1_2_1);
  assign state_out_3_2_1 = (((mul2_75_port_byte_out_1 ^ mul3_75_port_byte_out_1) ^ port_state_in_1_2_1) ^ port_state_in_2_2_1);
  assign state_out_0_2_2 = (((mul2_72_port_byte_out_2 ^ mul3_72_port_byte_out_2) ^ port_state_in_2_2_2) ^ port_state_in_3_2_2);
  assign state_out_1_2_2 = (((mul2_73_port_byte_out_2 ^ mul3_73_port_byte_out_2) ^ port_state_in_0_2_2) ^ port_state_in_3_2_2);
  assign state_out_2_2_2 = (((mul2_74_port_byte_out_2 ^ mul3_74_port_byte_out_2) ^ port_state_in_0_2_2) ^ port_state_in_1_2_2);
  assign state_out_3_2_2 = (((mul2_75_port_byte_out_2 ^ mul3_75_port_byte_out_2) ^ port_state_in_1_2_2) ^ port_state_in_2_2_2);
  assign state_out_0_2_3 = (((mul2_72_port_byte_out_3 ^ mul3_72_port_byte_out_3) ^ port_state_in_2_2_3) ^ port_state_in_3_2_3);
  assign state_out_1_2_3 = (((mul2_73_port_byte_out_3 ^ mul3_73_port_byte_out_3) ^ port_state_in_0_2_3) ^ port_state_in_3_2_3);
  assign state_out_2_2_3 = (((mul2_74_port_byte_out_3 ^ mul3_74_port_byte_out_3) ^ port_state_in_0_2_3) ^ port_state_in_1_2_3);
  assign state_out_3_2_3 = (((mul2_75_port_byte_out_3 ^ mul3_75_port_byte_out_3) ^ port_state_in_1_2_3) ^ port_state_in_2_2_3);
  assign state_out_0_2_4 = (((mul2_72_port_byte_out_4 ^ mul3_72_port_byte_out_4) ^ port_state_in_2_2_4) ^ port_state_in_3_2_4);
  assign state_out_1_2_4 = (((mul2_73_port_byte_out_4 ^ mul3_73_port_byte_out_4) ^ port_state_in_0_2_4) ^ port_state_in_3_2_4);
  assign state_out_2_2_4 = (((mul2_74_port_byte_out_4 ^ mul3_74_port_byte_out_4) ^ port_state_in_0_2_4) ^ port_state_in_1_2_4);
  assign state_out_3_2_4 = (((mul2_75_port_byte_out_4 ^ mul3_75_port_byte_out_4) ^ port_state_in_1_2_4) ^ port_state_in_2_2_4);
  assign state_out_0_2_5 = (((mul2_72_port_byte_out_5 ^ mul3_72_port_byte_out_5) ^ port_state_in_2_2_5) ^ port_state_in_3_2_5);
  assign state_out_1_2_5 = (((mul2_73_port_byte_out_5 ^ mul3_73_port_byte_out_5) ^ port_state_in_0_2_5) ^ port_state_in_3_2_5);
  assign state_out_2_2_5 = (((mul2_74_port_byte_out_5 ^ mul3_74_port_byte_out_5) ^ port_state_in_0_2_5) ^ port_state_in_1_2_5);
  assign state_out_3_2_5 = (((mul2_75_port_byte_out_5 ^ mul3_75_port_byte_out_5) ^ port_state_in_1_2_5) ^ port_state_in_2_2_5);
  assign state_out_0_2_6 = (((mul2_72_port_byte_out_6 ^ mul3_72_port_byte_out_6) ^ port_state_in_2_2_6) ^ port_state_in_3_2_6);
  assign state_out_1_2_6 = (((mul2_73_port_byte_out_6 ^ mul3_73_port_byte_out_6) ^ port_state_in_0_2_6) ^ port_state_in_3_2_6);
  assign state_out_2_2_6 = (((mul2_74_port_byte_out_6 ^ mul3_74_port_byte_out_6) ^ port_state_in_0_2_6) ^ port_state_in_1_2_6);
  assign state_out_3_2_6 = (((mul2_75_port_byte_out_6 ^ mul3_75_port_byte_out_6) ^ port_state_in_1_2_6) ^ port_state_in_2_2_6);
  assign state_out_0_2_7 = (((mul2_72_port_byte_out_7 ^ mul3_72_port_byte_out_7) ^ port_state_in_2_2_7) ^ port_state_in_3_2_7);
  assign state_out_1_2_7 = (((mul2_73_port_byte_out_7 ^ mul3_73_port_byte_out_7) ^ port_state_in_0_2_7) ^ port_state_in_3_2_7);
  assign state_out_2_2_7 = (((mul2_74_port_byte_out_7 ^ mul3_74_port_byte_out_7) ^ port_state_in_0_2_7) ^ port_state_in_1_2_7);
  assign state_out_3_2_7 = (((mul2_75_port_byte_out_7 ^ mul3_75_port_byte_out_7) ^ port_state_in_1_2_7) ^ port_state_in_2_2_7);
  assign state_out_0_3_0 = (((mul2_76_port_byte_out_0 ^ mul3_76_port_byte_out_0) ^ port_state_in_2_3_0) ^ port_state_in_3_3_0);
  assign state_out_1_3_0 = (((mul2_77_port_byte_out_0 ^ mul3_77_port_byte_out_0) ^ port_state_in_0_3_0) ^ port_state_in_3_3_0);
  assign state_out_2_3_0 = (((mul2_78_port_byte_out_0 ^ mul3_78_port_byte_out_0) ^ port_state_in_0_3_0) ^ port_state_in_1_3_0);
  assign state_out_3_3_0 = (((mul2_79_port_byte_out_0 ^ mul3_79_port_byte_out_0) ^ port_state_in_1_3_0) ^ port_state_in_2_3_0);
  assign state_out_0_3_1 = (((mul2_76_port_byte_out_1 ^ mul3_76_port_byte_out_1) ^ port_state_in_2_3_1) ^ port_state_in_3_3_1);
  assign state_out_1_3_1 = (((mul2_77_port_byte_out_1 ^ mul3_77_port_byte_out_1) ^ port_state_in_0_3_1) ^ port_state_in_3_3_1);
  assign state_out_2_3_1 = (((mul2_78_port_byte_out_1 ^ mul3_78_port_byte_out_1) ^ port_state_in_0_3_1) ^ port_state_in_1_3_1);
  assign state_out_3_3_1 = (((mul2_79_port_byte_out_1 ^ mul3_79_port_byte_out_1) ^ port_state_in_1_3_1) ^ port_state_in_2_3_1);
  assign state_out_0_3_2 = (((mul2_76_port_byte_out_2 ^ mul3_76_port_byte_out_2) ^ port_state_in_2_3_2) ^ port_state_in_3_3_2);
  assign state_out_1_3_2 = (((mul2_77_port_byte_out_2 ^ mul3_77_port_byte_out_2) ^ port_state_in_0_3_2) ^ port_state_in_3_3_2);
  assign state_out_2_3_2 = (((mul2_78_port_byte_out_2 ^ mul3_78_port_byte_out_2) ^ port_state_in_0_3_2) ^ port_state_in_1_3_2);
  assign state_out_3_3_2 = (((mul2_79_port_byte_out_2 ^ mul3_79_port_byte_out_2) ^ port_state_in_1_3_2) ^ port_state_in_2_3_2);
  assign state_out_0_3_3 = (((mul2_76_port_byte_out_3 ^ mul3_76_port_byte_out_3) ^ port_state_in_2_3_3) ^ port_state_in_3_3_3);
  assign state_out_1_3_3 = (((mul2_77_port_byte_out_3 ^ mul3_77_port_byte_out_3) ^ port_state_in_0_3_3) ^ port_state_in_3_3_3);
  assign state_out_2_3_3 = (((mul2_78_port_byte_out_3 ^ mul3_78_port_byte_out_3) ^ port_state_in_0_3_3) ^ port_state_in_1_3_3);
  assign state_out_3_3_3 = (((mul2_79_port_byte_out_3 ^ mul3_79_port_byte_out_3) ^ port_state_in_1_3_3) ^ port_state_in_2_3_3);
  assign state_out_0_3_4 = (((mul2_76_port_byte_out_4 ^ mul3_76_port_byte_out_4) ^ port_state_in_2_3_4) ^ port_state_in_3_3_4);
  assign state_out_1_3_4 = (((mul2_77_port_byte_out_4 ^ mul3_77_port_byte_out_4) ^ port_state_in_0_3_4) ^ port_state_in_3_3_4);
  assign state_out_2_3_4 = (((mul2_78_port_byte_out_4 ^ mul3_78_port_byte_out_4) ^ port_state_in_0_3_4) ^ port_state_in_1_3_4);
  assign state_out_3_3_4 = (((mul2_79_port_byte_out_4 ^ mul3_79_port_byte_out_4) ^ port_state_in_1_3_4) ^ port_state_in_2_3_4);
  assign state_out_0_3_5 = (((mul2_76_port_byte_out_5 ^ mul3_76_port_byte_out_5) ^ port_state_in_2_3_5) ^ port_state_in_3_3_5);
  assign state_out_1_3_5 = (((mul2_77_port_byte_out_5 ^ mul3_77_port_byte_out_5) ^ port_state_in_0_3_5) ^ port_state_in_3_3_5);
  assign state_out_2_3_5 = (((mul2_78_port_byte_out_5 ^ mul3_78_port_byte_out_5) ^ port_state_in_0_3_5) ^ port_state_in_1_3_5);
  assign state_out_3_3_5 = (((mul2_79_port_byte_out_5 ^ mul3_79_port_byte_out_5) ^ port_state_in_1_3_5) ^ port_state_in_2_3_5);
  assign state_out_0_3_6 = (((mul2_76_port_byte_out_6 ^ mul3_76_port_byte_out_6) ^ port_state_in_2_3_6) ^ port_state_in_3_3_6);
  assign state_out_1_3_6 = (((mul2_77_port_byte_out_6 ^ mul3_77_port_byte_out_6) ^ port_state_in_0_3_6) ^ port_state_in_3_3_6);
  assign state_out_2_3_6 = (((mul2_78_port_byte_out_6 ^ mul3_78_port_byte_out_6) ^ port_state_in_0_3_6) ^ port_state_in_1_3_6);
  assign state_out_3_3_6 = (((mul2_79_port_byte_out_6 ^ mul3_79_port_byte_out_6) ^ port_state_in_1_3_6) ^ port_state_in_2_3_6);
  assign state_out_0_3_7 = (((mul2_76_port_byte_out_7 ^ mul3_76_port_byte_out_7) ^ port_state_in_2_3_7) ^ port_state_in_3_3_7);
  assign state_out_1_3_7 = (((mul2_77_port_byte_out_7 ^ mul3_77_port_byte_out_7) ^ port_state_in_0_3_7) ^ port_state_in_3_3_7);
  assign state_out_2_3_7 = (((mul2_78_port_byte_out_7 ^ mul3_78_port_byte_out_7) ^ port_state_in_0_3_7) ^ port_state_in_1_3_7);
  assign state_out_3_3_7 = (((mul2_79_port_byte_out_7 ^ mul3_79_port_byte_out_7) ^ port_state_in_1_3_7) ^ port_state_in_2_3_7);
  assign state_out_4_0_0 = (((mul2_80_port_byte_out_0 ^ mul3_80_port_byte_out_0) ^ port_state_in_6_0_0) ^ port_state_in_7_0_0);
  assign state_out_5_0_0 = (((mul2_81_port_byte_out_0 ^ mul3_81_port_byte_out_0) ^ port_state_in_4_0_0) ^ port_state_in_7_0_0);
  assign state_out_6_0_0 = (((mul2_82_port_byte_out_0 ^ mul3_82_port_byte_out_0) ^ port_state_in_4_0_0) ^ port_state_in_5_0_0);
  assign state_out_7_0_0 = (((mul2_83_port_byte_out_0 ^ mul3_83_port_byte_out_0) ^ port_state_in_5_0_0) ^ port_state_in_6_0_0);
  assign state_out_4_0_1 = (((mul2_80_port_byte_out_1 ^ mul3_80_port_byte_out_1) ^ port_state_in_6_0_1) ^ port_state_in_7_0_1);
  assign state_out_5_0_1 = (((mul2_81_port_byte_out_1 ^ mul3_81_port_byte_out_1) ^ port_state_in_4_0_1) ^ port_state_in_7_0_1);
  assign state_out_6_0_1 = (((mul2_82_port_byte_out_1 ^ mul3_82_port_byte_out_1) ^ port_state_in_4_0_1) ^ port_state_in_5_0_1);
  assign state_out_7_0_1 = (((mul2_83_port_byte_out_1 ^ mul3_83_port_byte_out_1) ^ port_state_in_5_0_1) ^ port_state_in_6_0_1);
  assign state_out_4_0_2 = (((mul2_80_port_byte_out_2 ^ mul3_80_port_byte_out_2) ^ port_state_in_6_0_2) ^ port_state_in_7_0_2);
  assign state_out_5_0_2 = (((mul2_81_port_byte_out_2 ^ mul3_81_port_byte_out_2) ^ port_state_in_4_0_2) ^ port_state_in_7_0_2);
  assign state_out_6_0_2 = (((mul2_82_port_byte_out_2 ^ mul3_82_port_byte_out_2) ^ port_state_in_4_0_2) ^ port_state_in_5_0_2);
  assign state_out_7_0_2 = (((mul2_83_port_byte_out_2 ^ mul3_83_port_byte_out_2) ^ port_state_in_5_0_2) ^ port_state_in_6_0_2);
  assign state_out_4_0_3 = (((mul2_80_port_byte_out_3 ^ mul3_80_port_byte_out_3) ^ port_state_in_6_0_3) ^ port_state_in_7_0_3);
  assign state_out_5_0_3 = (((mul2_81_port_byte_out_3 ^ mul3_81_port_byte_out_3) ^ port_state_in_4_0_3) ^ port_state_in_7_0_3);
  assign state_out_6_0_3 = (((mul2_82_port_byte_out_3 ^ mul3_82_port_byte_out_3) ^ port_state_in_4_0_3) ^ port_state_in_5_0_3);
  assign state_out_7_0_3 = (((mul2_83_port_byte_out_3 ^ mul3_83_port_byte_out_3) ^ port_state_in_5_0_3) ^ port_state_in_6_0_3);
  assign state_out_4_0_4 = (((mul2_80_port_byte_out_4 ^ mul3_80_port_byte_out_4) ^ port_state_in_6_0_4) ^ port_state_in_7_0_4);
  assign state_out_5_0_4 = (((mul2_81_port_byte_out_4 ^ mul3_81_port_byte_out_4) ^ port_state_in_4_0_4) ^ port_state_in_7_0_4);
  assign state_out_6_0_4 = (((mul2_82_port_byte_out_4 ^ mul3_82_port_byte_out_4) ^ port_state_in_4_0_4) ^ port_state_in_5_0_4);
  assign state_out_7_0_4 = (((mul2_83_port_byte_out_4 ^ mul3_83_port_byte_out_4) ^ port_state_in_5_0_4) ^ port_state_in_6_0_4);
  assign state_out_4_0_5 = (((mul2_80_port_byte_out_5 ^ mul3_80_port_byte_out_5) ^ port_state_in_6_0_5) ^ port_state_in_7_0_5);
  assign state_out_5_0_5 = (((mul2_81_port_byte_out_5 ^ mul3_81_port_byte_out_5) ^ port_state_in_4_0_5) ^ port_state_in_7_0_5);
  assign state_out_6_0_5 = (((mul2_82_port_byte_out_5 ^ mul3_82_port_byte_out_5) ^ port_state_in_4_0_5) ^ port_state_in_5_0_5);
  assign state_out_7_0_5 = (((mul2_83_port_byte_out_5 ^ mul3_83_port_byte_out_5) ^ port_state_in_5_0_5) ^ port_state_in_6_0_5);
  assign state_out_4_0_6 = (((mul2_80_port_byte_out_6 ^ mul3_80_port_byte_out_6) ^ port_state_in_6_0_6) ^ port_state_in_7_0_6);
  assign state_out_5_0_6 = (((mul2_81_port_byte_out_6 ^ mul3_81_port_byte_out_6) ^ port_state_in_4_0_6) ^ port_state_in_7_0_6);
  assign state_out_6_0_6 = (((mul2_82_port_byte_out_6 ^ mul3_82_port_byte_out_6) ^ port_state_in_4_0_6) ^ port_state_in_5_0_6);
  assign state_out_7_0_6 = (((mul2_83_port_byte_out_6 ^ mul3_83_port_byte_out_6) ^ port_state_in_5_0_6) ^ port_state_in_6_0_6);
  assign state_out_4_0_7 = (((mul2_80_port_byte_out_7 ^ mul3_80_port_byte_out_7) ^ port_state_in_6_0_7) ^ port_state_in_7_0_7);
  assign state_out_5_0_7 = (((mul2_81_port_byte_out_7 ^ mul3_81_port_byte_out_7) ^ port_state_in_4_0_7) ^ port_state_in_7_0_7);
  assign state_out_6_0_7 = (((mul2_82_port_byte_out_7 ^ mul3_82_port_byte_out_7) ^ port_state_in_4_0_7) ^ port_state_in_5_0_7);
  assign state_out_7_0_7 = (((mul2_83_port_byte_out_7 ^ mul3_83_port_byte_out_7) ^ port_state_in_5_0_7) ^ port_state_in_6_0_7);
  assign state_out_4_1_0 = (((mul2_84_port_byte_out_0 ^ mul3_84_port_byte_out_0) ^ port_state_in_6_1_0) ^ port_state_in_7_1_0);
  assign state_out_5_1_0 = (((mul2_85_port_byte_out_0 ^ mul3_85_port_byte_out_0) ^ port_state_in_4_1_0) ^ port_state_in_7_1_0);
  assign state_out_6_1_0 = (((mul2_86_port_byte_out_0 ^ mul3_86_port_byte_out_0) ^ port_state_in_4_1_0) ^ port_state_in_5_1_0);
  assign state_out_7_1_0 = (((mul2_87_port_byte_out_0 ^ mul3_87_port_byte_out_0) ^ port_state_in_5_1_0) ^ port_state_in_6_1_0);
  assign state_out_4_1_1 = (((mul2_84_port_byte_out_1 ^ mul3_84_port_byte_out_1) ^ port_state_in_6_1_1) ^ port_state_in_7_1_1);
  assign state_out_5_1_1 = (((mul2_85_port_byte_out_1 ^ mul3_85_port_byte_out_1) ^ port_state_in_4_1_1) ^ port_state_in_7_1_1);
  assign state_out_6_1_1 = (((mul2_86_port_byte_out_1 ^ mul3_86_port_byte_out_1) ^ port_state_in_4_1_1) ^ port_state_in_5_1_1);
  assign state_out_7_1_1 = (((mul2_87_port_byte_out_1 ^ mul3_87_port_byte_out_1) ^ port_state_in_5_1_1) ^ port_state_in_6_1_1);
  assign state_out_4_1_2 = (((mul2_84_port_byte_out_2 ^ mul3_84_port_byte_out_2) ^ port_state_in_6_1_2) ^ port_state_in_7_1_2);
  assign state_out_5_1_2 = (((mul2_85_port_byte_out_2 ^ mul3_85_port_byte_out_2) ^ port_state_in_4_1_2) ^ port_state_in_7_1_2);
  assign state_out_6_1_2 = (((mul2_86_port_byte_out_2 ^ mul3_86_port_byte_out_2) ^ port_state_in_4_1_2) ^ port_state_in_5_1_2);
  assign state_out_7_1_2 = (((mul2_87_port_byte_out_2 ^ mul3_87_port_byte_out_2) ^ port_state_in_5_1_2) ^ port_state_in_6_1_2);
  assign state_out_4_1_3 = (((mul2_84_port_byte_out_3 ^ mul3_84_port_byte_out_3) ^ port_state_in_6_1_3) ^ port_state_in_7_1_3);
  assign state_out_5_1_3 = (((mul2_85_port_byte_out_3 ^ mul3_85_port_byte_out_3) ^ port_state_in_4_1_3) ^ port_state_in_7_1_3);
  assign state_out_6_1_3 = (((mul2_86_port_byte_out_3 ^ mul3_86_port_byte_out_3) ^ port_state_in_4_1_3) ^ port_state_in_5_1_3);
  assign state_out_7_1_3 = (((mul2_87_port_byte_out_3 ^ mul3_87_port_byte_out_3) ^ port_state_in_5_1_3) ^ port_state_in_6_1_3);
  assign state_out_4_1_4 = (((mul2_84_port_byte_out_4 ^ mul3_84_port_byte_out_4) ^ port_state_in_6_1_4) ^ port_state_in_7_1_4);
  assign state_out_5_1_4 = (((mul2_85_port_byte_out_4 ^ mul3_85_port_byte_out_4) ^ port_state_in_4_1_4) ^ port_state_in_7_1_4);
  assign state_out_6_1_4 = (((mul2_86_port_byte_out_4 ^ mul3_86_port_byte_out_4) ^ port_state_in_4_1_4) ^ port_state_in_5_1_4);
  assign state_out_7_1_4 = (((mul2_87_port_byte_out_4 ^ mul3_87_port_byte_out_4) ^ port_state_in_5_1_4) ^ port_state_in_6_1_4);
  assign state_out_4_1_5 = (((mul2_84_port_byte_out_5 ^ mul3_84_port_byte_out_5) ^ port_state_in_6_1_5) ^ port_state_in_7_1_5);
  assign state_out_5_1_5 = (((mul2_85_port_byte_out_5 ^ mul3_85_port_byte_out_5) ^ port_state_in_4_1_5) ^ port_state_in_7_1_5);
  assign state_out_6_1_5 = (((mul2_86_port_byte_out_5 ^ mul3_86_port_byte_out_5) ^ port_state_in_4_1_5) ^ port_state_in_5_1_5);
  assign state_out_7_1_5 = (((mul2_87_port_byte_out_5 ^ mul3_87_port_byte_out_5) ^ port_state_in_5_1_5) ^ port_state_in_6_1_5);
  assign state_out_4_1_6 = (((mul2_84_port_byte_out_6 ^ mul3_84_port_byte_out_6) ^ port_state_in_6_1_6) ^ port_state_in_7_1_6);
  assign state_out_5_1_6 = (((mul2_85_port_byte_out_6 ^ mul3_85_port_byte_out_6) ^ port_state_in_4_1_6) ^ port_state_in_7_1_6);
  assign state_out_6_1_6 = (((mul2_86_port_byte_out_6 ^ mul3_86_port_byte_out_6) ^ port_state_in_4_1_6) ^ port_state_in_5_1_6);
  assign state_out_7_1_6 = (((mul2_87_port_byte_out_6 ^ mul3_87_port_byte_out_6) ^ port_state_in_5_1_6) ^ port_state_in_6_1_6);
  assign state_out_4_1_7 = (((mul2_84_port_byte_out_7 ^ mul3_84_port_byte_out_7) ^ port_state_in_6_1_7) ^ port_state_in_7_1_7);
  assign state_out_5_1_7 = (((mul2_85_port_byte_out_7 ^ mul3_85_port_byte_out_7) ^ port_state_in_4_1_7) ^ port_state_in_7_1_7);
  assign state_out_6_1_7 = (((mul2_86_port_byte_out_7 ^ mul3_86_port_byte_out_7) ^ port_state_in_4_1_7) ^ port_state_in_5_1_7);
  assign state_out_7_1_7 = (((mul2_87_port_byte_out_7 ^ mul3_87_port_byte_out_7) ^ port_state_in_5_1_7) ^ port_state_in_6_1_7);
  assign state_out_4_2_0 = (((mul2_88_port_byte_out_0 ^ mul3_88_port_byte_out_0) ^ port_state_in_6_2_0) ^ port_state_in_7_2_0);
  assign state_out_5_2_0 = (((mul2_89_port_byte_out_0 ^ mul3_89_port_byte_out_0) ^ port_state_in_4_2_0) ^ port_state_in_7_2_0);
  assign state_out_6_2_0 = (((mul2_90_port_byte_out_0 ^ mul3_90_port_byte_out_0) ^ port_state_in_4_2_0) ^ port_state_in_5_2_0);
  assign state_out_7_2_0 = (((mul2_91_port_byte_out_0 ^ mul3_91_port_byte_out_0) ^ port_state_in_5_2_0) ^ port_state_in_6_2_0);
  assign state_out_4_2_1 = (((mul2_88_port_byte_out_1 ^ mul3_88_port_byte_out_1) ^ port_state_in_6_2_1) ^ port_state_in_7_2_1);
  assign state_out_5_2_1 = (((mul2_89_port_byte_out_1 ^ mul3_89_port_byte_out_1) ^ port_state_in_4_2_1) ^ port_state_in_7_2_1);
  assign state_out_6_2_1 = (((mul2_90_port_byte_out_1 ^ mul3_90_port_byte_out_1) ^ port_state_in_4_2_1) ^ port_state_in_5_2_1);
  assign state_out_7_2_1 = (((mul2_91_port_byte_out_1 ^ mul3_91_port_byte_out_1) ^ port_state_in_5_2_1) ^ port_state_in_6_2_1);
  assign state_out_4_2_2 = (((mul2_88_port_byte_out_2 ^ mul3_88_port_byte_out_2) ^ port_state_in_6_2_2) ^ port_state_in_7_2_2);
  assign state_out_5_2_2 = (((mul2_89_port_byte_out_2 ^ mul3_89_port_byte_out_2) ^ port_state_in_4_2_2) ^ port_state_in_7_2_2);
  assign state_out_6_2_2 = (((mul2_90_port_byte_out_2 ^ mul3_90_port_byte_out_2) ^ port_state_in_4_2_2) ^ port_state_in_5_2_2);
  assign state_out_7_2_2 = (((mul2_91_port_byte_out_2 ^ mul3_91_port_byte_out_2) ^ port_state_in_5_2_2) ^ port_state_in_6_2_2);
  assign state_out_4_2_3 = (((mul2_88_port_byte_out_3 ^ mul3_88_port_byte_out_3) ^ port_state_in_6_2_3) ^ port_state_in_7_2_3);
  assign state_out_5_2_3 = (((mul2_89_port_byte_out_3 ^ mul3_89_port_byte_out_3) ^ port_state_in_4_2_3) ^ port_state_in_7_2_3);
  assign state_out_6_2_3 = (((mul2_90_port_byte_out_3 ^ mul3_90_port_byte_out_3) ^ port_state_in_4_2_3) ^ port_state_in_5_2_3);
  assign state_out_7_2_3 = (((mul2_91_port_byte_out_3 ^ mul3_91_port_byte_out_3) ^ port_state_in_5_2_3) ^ port_state_in_6_2_3);
  assign state_out_4_2_4 = (((mul2_88_port_byte_out_4 ^ mul3_88_port_byte_out_4) ^ port_state_in_6_2_4) ^ port_state_in_7_2_4);
  assign state_out_5_2_4 = (((mul2_89_port_byte_out_4 ^ mul3_89_port_byte_out_4) ^ port_state_in_4_2_4) ^ port_state_in_7_2_4);
  assign state_out_6_2_4 = (((mul2_90_port_byte_out_4 ^ mul3_90_port_byte_out_4) ^ port_state_in_4_2_4) ^ port_state_in_5_2_4);
  assign state_out_7_2_4 = (((mul2_91_port_byte_out_4 ^ mul3_91_port_byte_out_4) ^ port_state_in_5_2_4) ^ port_state_in_6_2_4);
  assign state_out_4_2_5 = (((mul2_88_port_byte_out_5 ^ mul3_88_port_byte_out_5) ^ port_state_in_6_2_5) ^ port_state_in_7_2_5);
  assign state_out_5_2_5 = (((mul2_89_port_byte_out_5 ^ mul3_89_port_byte_out_5) ^ port_state_in_4_2_5) ^ port_state_in_7_2_5);
  assign state_out_6_2_5 = (((mul2_90_port_byte_out_5 ^ mul3_90_port_byte_out_5) ^ port_state_in_4_2_5) ^ port_state_in_5_2_5);
  assign state_out_7_2_5 = (((mul2_91_port_byte_out_5 ^ mul3_91_port_byte_out_5) ^ port_state_in_5_2_5) ^ port_state_in_6_2_5);
  assign state_out_4_2_6 = (((mul2_88_port_byte_out_6 ^ mul3_88_port_byte_out_6) ^ port_state_in_6_2_6) ^ port_state_in_7_2_6);
  assign state_out_5_2_6 = (((mul2_89_port_byte_out_6 ^ mul3_89_port_byte_out_6) ^ port_state_in_4_2_6) ^ port_state_in_7_2_6);
  assign state_out_6_2_6 = (((mul2_90_port_byte_out_6 ^ mul3_90_port_byte_out_6) ^ port_state_in_4_2_6) ^ port_state_in_5_2_6);
  assign state_out_7_2_6 = (((mul2_91_port_byte_out_6 ^ mul3_91_port_byte_out_6) ^ port_state_in_5_2_6) ^ port_state_in_6_2_6);
  assign state_out_4_2_7 = (((mul2_88_port_byte_out_7 ^ mul3_88_port_byte_out_7) ^ port_state_in_6_2_7) ^ port_state_in_7_2_7);
  assign state_out_5_2_7 = (((mul2_89_port_byte_out_7 ^ mul3_89_port_byte_out_7) ^ port_state_in_4_2_7) ^ port_state_in_7_2_7);
  assign state_out_6_2_7 = (((mul2_90_port_byte_out_7 ^ mul3_90_port_byte_out_7) ^ port_state_in_4_2_7) ^ port_state_in_5_2_7);
  assign state_out_7_2_7 = (((mul2_91_port_byte_out_7 ^ mul3_91_port_byte_out_7) ^ port_state_in_5_2_7) ^ port_state_in_6_2_7);
  assign state_out_4_3_0 = (((mul2_92_port_byte_out_0 ^ mul3_92_port_byte_out_0) ^ port_state_in_6_3_0) ^ port_state_in_7_3_0);
  assign state_out_5_3_0 = (((mul2_93_port_byte_out_0 ^ mul3_93_port_byte_out_0) ^ port_state_in_4_3_0) ^ port_state_in_7_3_0);
  assign state_out_6_3_0 = (((mul2_94_port_byte_out_0 ^ mul3_94_port_byte_out_0) ^ port_state_in_4_3_0) ^ port_state_in_5_3_0);
  assign state_out_7_3_0 = (((mul2_95_port_byte_out_0 ^ mul3_95_port_byte_out_0) ^ port_state_in_5_3_0) ^ port_state_in_6_3_0);
  assign state_out_4_3_1 = (((mul2_92_port_byte_out_1 ^ mul3_92_port_byte_out_1) ^ port_state_in_6_3_1) ^ port_state_in_7_3_1);
  assign state_out_5_3_1 = (((mul2_93_port_byte_out_1 ^ mul3_93_port_byte_out_1) ^ port_state_in_4_3_1) ^ port_state_in_7_3_1);
  assign state_out_6_3_1 = (((mul2_94_port_byte_out_1 ^ mul3_94_port_byte_out_1) ^ port_state_in_4_3_1) ^ port_state_in_5_3_1);
  assign state_out_7_3_1 = (((mul2_95_port_byte_out_1 ^ mul3_95_port_byte_out_1) ^ port_state_in_5_3_1) ^ port_state_in_6_3_1);
  assign state_out_4_3_2 = (((mul2_92_port_byte_out_2 ^ mul3_92_port_byte_out_2) ^ port_state_in_6_3_2) ^ port_state_in_7_3_2);
  assign state_out_5_3_2 = (((mul2_93_port_byte_out_2 ^ mul3_93_port_byte_out_2) ^ port_state_in_4_3_2) ^ port_state_in_7_3_2);
  assign state_out_6_3_2 = (((mul2_94_port_byte_out_2 ^ mul3_94_port_byte_out_2) ^ port_state_in_4_3_2) ^ port_state_in_5_3_2);
  assign state_out_7_3_2 = (((mul2_95_port_byte_out_2 ^ mul3_95_port_byte_out_2) ^ port_state_in_5_3_2) ^ port_state_in_6_3_2);
  assign state_out_4_3_3 = (((mul2_92_port_byte_out_3 ^ mul3_92_port_byte_out_3) ^ port_state_in_6_3_3) ^ port_state_in_7_3_3);
  assign state_out_5_3_3 = (((mul2_93_port_byte_out_3 ^ mul3_93_port_byte_out_3) ^ port_state_in_4_3_3) ^ port_state_in_7_3_3);
  assign state_out_6_3_3 = (((mul2_94_port_byte_out_3 ^ mul3_94_port_byte_out_3) ^ port_state_in_4_3_3) ^ port_state_in_5_3_3);
  assign state_out_7_3_3 = (((mul2_95_port_byte_out_3 ^ mul3_95_port_byte_out_3) ^ port_state_in_5_3_3) ^ port_state_in_6_3_3);
  assign state_out_4_3_4 = (((mul2_92_port_byte_out_4 ^ mul3_92_port_byte_out_4) ^ port_state_in_6_3_4) ^ port_state_in_7_3_4);
  assign state_out_5_3_4 = (((mul2_93_port_byte_out_4 ^ mul3_93_port_byte_out_4) ^ port_state_in_4_3_4) ^ port_state_in_7_3_4);
  assign state_out_6_3_4 = (((mul2_94_port_byte_out_4 ^ mul3_94_port_byte_out_4) ^ port_state_in_4_3_4) ^ port_state_in_5_3_4);
  assign state_out_7_3_4 = (((mul2_95_port_byte_out_4 ^ mul3_95_port_byte_out_4) ^ port_state_in_5_3_4) ^ port_state_in_6_3_4);
  assign state_out_4_3_5 = (((mul2_92_port_byte_out_5 ^ mul3_92_port_byte_out_5) ^ port_state_in_6_3_5) ^ port_state_in_7_3_5);
  assign state_out_5_3_5 = (((mul2_93_port_byte_out_5 ^ mul3_93_port_byte_out_5) ^ port_state_in_4_3_5) ^ port_state_in_7_3_5);
  assign state_out_6_3_5 = (((mul2_94_port_byte_out_5 ^ mul3_94_port_byte_out_5) ^ port_state_in_4_3_5) ^ port_state_in_5_3_5);
  assign state_out_7_3_5 = (((mul2_95_port_byte_out_5 ^ mul3_95_port_byte_out_5) ^ port_state_in_5_3_5) ^ port_state_in_6_3_5);
  assign state_out_4_3_6 = (((mul2_92_port_byte_out_6 ^ mul3_92_port_byte_out_6) ^ port_state_in_6_3_6) ^ port_state_in_7_3_6);
  assign state_out_5_3_6 = (((mul2_93_port_byte_out_6 ^ mul3_93_port_byte_out_6) ^ port_state_in_4_3_6) ^ port_state_in_7_3_6);
  assign state_out_6_3_6 = (((mul2_94_port_byte_out_6 ^ mul3_94_port_byte_out_6) ^ port_state_in_4_3_6) ^ port_state_in_5_3_6);
  assign state_out_7_3_6 = (((mul2_95_port_byte_out_6 ^ mul3_95_port_byte_out_6) ^ port_state_in_5_3_6) ^ port_state_in_6_3_6);
  assign state_out_4_3_7 = (((mul2_92_port_byte_out_7 ^ mul3_92_port_byte_out_7) ^ port_state_in_6_3_7) ^ port_state_in_7_3_7);
  assign state_out_5_3_7 = (((mul2_93_port_byte_out_7 ^ mul3_93_port_byte_out_7) ^ port_state_in_4_3_7) ^ port_state_in_7_3_7);
  assign state_out_6_3_7 = (((mul2_94_port_byte_out_7 ^ mul3_94_port_byte_out_7) ^ port_state_in_4_3_7) ^ port_state_in_5_3_7);
  assign state_out_7_3_7 = (((mul2_95_port_byte_out_7 ^ mul3_95_port_byte_out_7) ^ port_state_in_5_3_7) ^ port_state_in_6_3_7);
  assign state_out_8_0_0 = (((mul2_96_port_byte_out_0 ^ mul3_96_port_byte_out_0) ^ port_state_in_10_0_0) ^ port_state_in_11_0_0);
  assign state_out_9_0_0 = (((mul2_97_port_byte_out_0 ^ mul3_97_port_byte_out_0) ^ port_state_in_8_0_0) ^ port_state_in_11_0_0);
  assign state_out_10_0_0 = (((mul2_98_port_byte_out_0 ^ mul3_98_port_byte_out_0) ^ port_state_in_8_0_0) ^ port_state_in_9_0_0);
  assign state_out_11_0_0 = (((mul2_99_port_byte_out_0 ^ mul3_99_port_byte_out_0) ^ port_state_in_9_0_0) ^ port_state_in_10_0_0);
  assign state_out_8_0_1 = (((mul2_96_port_byte_out_1 ^ mul3_96_port_byte_out_1) ^ port_state_in_10_0_1) ^ port_state_in_11_0_1);
  assign state_out_9_0_1 = (((mul2_97_port_byte_out_1 ^ mul3_97_port_byte_out_1) ^ port_state_in_8_0_1) ^ port_state_in_11_0_1);
  assign state_out_10_0_1 = (((mul2_98_port_byte_out_1 ^ mul3_98_port_byte_out_1) ^ port_state_in_8_0_1) ^ port_state_in_9_0_1);
  assign state_out_11_0_1 = (((mul2_99_port_byte_out_1 ^ mul3_99_port_byte_out_1) ^ port_state_in_9_0_1) ^ port_state_in_10_0_1);
  assign state_out_8_0_2 = (((mul2_96_port_byte_out_2 ^ mul3_96_port_byte_out_2) ^ port_state_in_10_0_2) ^ port_state_in_11_0_2);
  assign state_out_9_0_2 = (((mul2_97_port_byte_out_2 ^ mul3_97_port_byte_out_2) ^ port_state_in_8_0_2) ^ port_state_in_11_0_2);
  assign state_out_10_0_2 = (((mul2_98_port_byte_out_2 ^ mul3_98_port_byte_out_2) ^ port_state_in_8_0_2) ^ port_state_in_9_0_2);
  assign state_out_11_0_2 = (((mul2_99_port_byte_out_2 ^ mul3_99_port_byte_out_2) ^ port_state_in_9_0_2) ^ port_state_in_10_0_2);
  assign state_out_8_0_3 = (((mul2_96_port_byte_out_3 ^ mul3_96_port_byte_out_3) ^ port_state_in_10_0_3) ^ port_state_in_11_0_3);
  assign state_out_9_0_3 = (((mul2_97_port_byte_out_3 ^ mul3_97_port_byte_out_3) ^ port_state_in_8_0_3) ^ port_state_in_11_0_3);
  assign state_out_10_0_3 = (((mul2_98_port_byte_out_3 ^ mul3_98_port_byte_out_3) ^ port_state_in_8_0_3) ^ port_state_in_9_0_3);
  assign state_out_11_0_3 = (((mul2_99_port_byte_out_3 ^ mul3_99_port_byte_out_3) ^ port_state_in_9_0_3) ^ port_state_in_10_0_3);
  assign state_out_8_0_4 = (((mul2_96_port_byte_out_4 ^ mul3_96_port_byte_out_4) ^ port_state_in_10_0_4) ^ port_state_in_11_0_4);
  assign state_out_9_0_4 = (((mul2_97_port_byte_out_4 ^ mul3_97_port_byte_out_4) ^ port_state_in_8_0_4) ^ port_state_in_11_0_4);
  assign state_out_10_0_4 = (((mul2_98_port_byte_out_4 ^ mul3_98_port_byte_out_4) ^ port_state_in_8_0_4) ^ port_state_in_9_0_4);
  assign state_out_11_0_4 = (((mul2_99_port_byte_out_4 ^ mul3_99_port_byte_out_4) ^ port_state_in_9_0_4) ^ port_state_in_10_0_4);
  assign state_out_8_0_5 = (((mul2_96_port_byte_out_5 ^ mul3_96_port_byte_out_5) ^ port_state_in_10_0_5) ^ port_state_in_11_0_5);
  assign state_out_9_0_5 = (((mul2_97_port_byte_out_5 ^ mul3_97_port_byte_out_5) ^ port_state_in_8_0_5) ^ port_state_in_11_0_5);
  assign state_out_10_0_5 = (((mul2_98_port_byte_out_5 ^ mul3_98_port_byte_out_5) ^ port_state_in_8_0_5) ^ port_state_in_9_0_5);
  assign state_out_11_0_5 = (((mul2_99_port_byte_out_5 ^ mul3_99_port_byte_out_5) ^ port_state_in_9_0_5) ^ port_state_in_10_0_5);
  assign state_out_8_0_6 = (((mul2_96_port_byte_out_6 ^ mul3_96_port_byte_out_6) ^ port_state_in_10_0_6) ^ port_state_in_11_0_6);
  assign state_out_9_0_6 = (((mul2_97_port_byte_out_6 ^ mul3_97_port_byte_out_6) ^ port_state_in_8_0_6) ^ port_state_in_11_0_6);
  assign state_out_10_0_6 = (((mul2_98_port_byte_out_6 ^ mul3_98_port_byte_out_6) ^ port_state_in_8_0_6) ^ port_state_in_9_0_6);
  assign state_out_11_0_6 = (((mul2_99_port_byte_out_6 ^ mul3_99_port_byte_out_6) ^ port_state_in_9_0_6) ^ port_state_in_10_0_6);
  assign state_out_8_0_7 = (((mul2_96_port_byte_out_7 ^ mul3_96_port_byte_out_7) ^ port_state_in_10_0_7) ^ port_state_in_11_0_7);
  assign state_out_9_0_7 = (((mul2_97_port_byte_out_7 ^ mul3_97_port_byte_out_7) ^ port_state_in_8_0_7) ^ port_state_in_11_0_7);
  assign state_out_10_0_7 = (((mul2_98_port_byte_out_7 ^ mul3_98_port_byte_out_7) ^ port_state_in_8_0_7) ^ port_state_in_9_0_7);
  assign state_out_11_0_7 = (((mul2_99_port_byte_out_7 ^ mul3_99_port_byte_out_7) ^ port_state_in_9_0_7) ^ port_state_in_10_0_7);
  assign state_out_8_1_0 = (((mul2_100_port_byte_out_0 ^ mul3_100_port_byte_out_0) ^ port_state_in_10_1_0) ^ port_state_in_11_1_0);
  assign state_out_9_1_0 = (((mul2_101_port_byte_out_0 ^ mul3_101_port_byte_out_0) ^ port_state_in_8_1_0) ^ port_state_in_11_1_0);
  assign state_out_10_1_0 = (((mul2_102_port_byte_out_0 ^ mul3_102_port_byte_out_0) ^ port_state_in_8_1_0) ^ port_state_in_9_1_0);
  assign state_out_11_1_0 = (((mul2_103_port_byte_out_0 ^ mul3_103_port_byte_out_0) ^ port_state_in_9_1_0) ^ port_state_in_10_1_0);
  assign state_out_8_1_1 = (((mul2_100_port_byte_out_1 ^ mul3_100_port_byte_out_1) ^ port_state_in_10_1_1) ^ port_state_in_11_1_1);
  assign state_out_9_1_1 = (((mul2_101_port_byte_out_1 ^ mul3_101_port_byte_out_1) ^ port_state_in_8_1_1) ^ port_state_in_11_1_1);
  assign state_out_10_1_1 = (((mul2_102_port_byte_out_1 ^ mul3_102_port_byte_out_1) ^ port_state_in_8_1_1) ^ port_state_in_9_1_1);
  assign state_out_11_1_1 = (((mul2_103_port_byte_out_1 ^ mul3_103_port_byte_out_1) ^ port_state_in_9_1_1) ^ port_state_in_10_1_1);
  assign state_out_8_1_2 = (((mul2_100_port_byte_out_2 ^ mul3_100_port_byte_out_2) ^ port_state_in_10_1_2) ^ port_state_in_11_1_2);
  assign state_out_9_1_2 = (((mul2_101_port_byte_out_2 ^ mul3_101_port_byte_out_2) ^ port_state_in_8_1_2) ^ port_state_in_11_1_2);
  assign state_out_10_1_2 = (((mul2_102_port_byte_out_2 ^ mul3_102_port_byte_out_2) ^ port_state_in_8_1_2) ^ port_state_in_9_1_2);
  assign state_out_11_1_2 = (((mul2_103_port_byte_out_2 ^ mul3_103_port_byte_out_2) ^ port_state_in_9_1_2) ^ port_state_in_10_1_2);
  assign state_out_8_1_3 = (((mul2_100_port_byte_out_3 ^ mul3_100_port_byte_out_3) ^ port_state_in_10_1_3) ^ port_state_in_11_1_3);
  assign state_out_9_1_3 = (((mul2_101_port_byte_out_3 ^ mul3_101_port_byte_out_3) ^ port_state_in_8_1_3) ^ port_state_in_11_1_3);
  assign state_out_10_1_3 = (((mul2_102_port_byte_out_3 ^ mul3_102_port_byte_out_3) ^ port_state_in_8_1_3) ^ port_state_in_9_1_3);
  assign state_out_11_1_3 = (((mul2_103_port_byte_out_3 ^ mul3_103_port_byte_out_3) ^ port_state_in_9_1_3) ^ port_state_in_10_1_3);
  assign state_out_8_1_4 = (((mul2_100_port_byte_out_4 ^ mul3_100_port_byte_out_4) ^ port_state_in_10_1_4) ^ port_state_in_11_1_4);
  assign state_out_9_1_4 = (((mul2_101_port_byte_out_4 ^ mul3_101_port_byte_out_4) ^ port_state_in_8_1_4) ^ port_state_in_11_1_4);
  assign state_out_10_1_4 = (((mul2_102_port_byte_out_4 ^ mul3_102_port_byte_out_4) ^ port_state_in_8_1_4) ^ port_state_in_9_1_4);
  assign state_out_11_1_4 = (((mul2_103_port_byte_out_4 ^ mul3_103_port_byte_out_4) ^ port_state_in_9_1_4) ^ port_state_in_10_1_4);
  assign state_out_8_1_5 = (((mul2_100_port_byte_out_5 ^ mul3_100_port_byte_out_5) ^ port_state_in_10_1_5) ^ port_state_in_11_1_5);
  assign state_out_9_1_5 = (((mul2_101_port_byte_out_5 ^ mul3_101_port_byte_out_5) ^ port_state_in_8_1_5) ^ port_state_in_11_1_5);
  assign state_out_10_1_5 = (((mul2_102_port_byte_out_5 ^ mul3_102_port_byte_out_5) ^ port_state_in_8_1_5) ^ port_state_in_9_1_5);
  assign state_out_11_1_5 = (((mul2_103_port_byte_out_5 ^ mul3_103_port_byte_out_5) ^ port_state_in_9_1_5) ^ port_state_in_10_1_5);
  assign state_out_8_1_6 = (((mul2_100_port_byte_out_6 ^ mul3_100_port_byte_out_6) ^ port_state_in_10_1_6) ^ port_state_in_11_1_6);
  assign state_out_9_1_6 = (((mul2_101_port_byte_out_6 ^ mul3_101_port_byte_out_6) ^ port_state_in_8_1_6) ^ port_state_in_11_1_6);
  assign state_out_10_1_6 = (((mul2_102_port_byte_out_6 ^ mul3_102_port_byte_out_6) ^ port_state_in_8_1_6) ^ port_state_in_9_1_6);
  assign state_out_11_1_6 = (((mul2_103_port_byte_out_6 ^ mul3_103_port_byte_out_6) ^ port_state_in_9_1_6) ^ port_state_in_10_1_6);
  assign state_out_8_1_7 = (((mul2_100_port_byte_out_7 ^ mul3_100_port_byte_out_7) ^ port_state_in_10_1_7) ^ port_state_in_11_1_7);
  assign state_out_9_1_7 = (((mul2_101_port_byte_out_7 ^ mul3_101_port_byte_out_7) ^ port_state_in_8_1_7) ^ port_state_in_11_1_7);
  assign state_out_10_1_7 = (((mul2_102_port_byte_out_7 ^ mul3_102_port_byte_out_7) ^ port_state_in_8_1_7) ^ port_state_in_9_1_7);
  assign state_out_11_1_7 = (((mul2_103_port_byte_out_7 ^ mul3_103_port_byte_out_7) ^ port_state_in_9_1_7) ^ port_state_in_10_1_7);
  assign state_out_8_2_0 = (((mul2_104_port_byte_out_0 ^ mul3_104_port_byte_out_0) ^ port_state_in_10_2_0) ^ port_state_in_11_2_0);
  assign state_out_9_2_0 = (((mul2_105_port_byte_out_0 ^ mul3_105_port_byte_out_0) ^ port_state_in_8_2_0) ^ port_state_in_11_2_0);
  assign state_out_10_2_0 = (((mul2_106_port_byte_out_0 ^ mul3_106_port_byte_out_0) ^ port_state_in_8_2_0) ^ port_state_in_9_2_0);
  assign state_out_11_2_0 = (((mul2_107_port_byte_out_0 ^ mul3_107_port_byte_out_0) ^ port_state_in_9_2_0) ^ port_state_in_10_2_0);
  assign state_out_8_2_1 = (((mul2_104_port_byte_out_1 ^ mul3_104_port_byte_out_1) ^ port_state_in_10_2_1) ^ port_state_in_11_2_1);
  assign state_out_9_2_1 = (((mul2_105_port_byte_out_1 ^ mul3_105_port_byte_out_1) ^ port_state_in_8_2_1) ^ port_state_in_11_2_1);
  assign state_out_10_2_1 = (((mul2_106_port_byte_out_1 ^ mul3_106_port_byte_out_1) ^ port_state_in_8_2_1) ^ port_state_in_9_2_1);
  assign state_out_11_2_1 = (((mul2_107_port_byte_out_1 ^ mul3_107_port_byte_out_1) ^ port_state_in_9_2_1) ^ port_state_in_10_2_1);
  assign state_out_8_2_2 = (((mul2_104_port_byte_out_2 ^ mul3_104_port_byte_out_2) ^ port_state_in_10_2_2) ^ port_state_in_11_2_2);
  assign state_out_9_2_2 = (((mul2_105_port_byte_out_2 ^ mul3_105_port_byte_out_2) ^ port_state_in_8_2_2) ^ port_state_in_11_2_2);
  assign state_out_10_2_2 = (((mul2_106_port_byte_out_2 ^ mul3_106_port_byte_out_2) ^ port_state_in_8_2_2) ^ port_state_in_9_2_2);
  assign state_out_11_2_2 = (((mul2_107_port_byte_out_2 ^ mul3_107_port_byte_out_2) ^ port_state_in_9_2_2) ^ port_state_in_10_2_2);
  assign state_out_8_2_3 = (((mul2_104_port_byte_out_3 ^ mul3_104_port_byte_out_3) ^ port_state_in_10_2_3) ^ port_state_in_11_2_3);
  assign state_out_9_2_3 = (((mul2_105_port_byte_out_3 ^ mul3_105_port_byte_out_3) ^ port_state_in_8_2_3) ^ port_state_in_11_2_3);
  assign state_out_10_2_3 = (((mul2_106_port_byte_out_3 ^ mul3_106_port_byte_out_3) ^ port_state_in_8_2_3) ^ port_state_in_9_2_3);
  assign state_out_11_2_3 = (((mul2_107_port_byte_out_3 ^ mul3_107_port_byte_out_3) ^ port_state_in_9_2_3) ^ port_state_in_10_2_3);
  assign state_out_8_2_4 = (((mul2_104_port_byte_out_4 ^ mul3_104_port_byte_out_4) ^ port_state_in_10_2_4) ^ port_state_in_11_2_4);
  assign state_out_9_2_4 = (((mul2_105_port_byte_out_4 ^ mul3_105_port_byte_out_4) ^ port_state_in_8_2_4) ^ port_state_in_11_2_4);
  assign state_out_10_2_4 = (((mul2_106_port_byte_out_4 ^ mul3_106_port_byte_out_4) ^ port_state_in_8_2_4) ^ port_state_in_9_2_4);
  assign state_out_11_2_4 = (((mul2_107_port_byte_out_4 ^ mul3_107_port_byte_out_4) ^ port_state_in_9_2_4) ^ port_state_in_10_2_4);
  assign state_out_8_2_5 = (((mul2_104_port_byte_out_5 ^ mul3_104_port_byte_out_5) ^ port_state_in_10_2_5) ^ port_state_in_11_2_5);
  assign state_out_9_2_5 = (((mul2_105_port_byte_out_5 ^ mul3_105_port_byte_out_5) ^ port_state_in_8_2_5) ^ port_state_in_11_2_5);
  assign state_out_10_2_5 = (((mul2_106_port_byte_out_5 ^ mul3_106_port_byte_out_5) ^ port_state_in_8_2_5) ^ port_state_in_9_2_5);
  assign state_out_11_2_5 = (((mul2_107_port_byte_out_5 ^ mul3_107_port_byte_out_5) ^ port_state_in_9_2_5) ^ port_state_in_10_2_5);
  assign state_out_8_2_6 = (((mul2_104_port_byte_out_6 ^ mul3_104_port_byte_out_6) ^ port_state_in_10_2_6) ^ port_state_in_11_2_6);
  assign state_out_9_2_6 = (((mul2_105_port_byte_out_6 ^ mul3_105_port_byte_out_6) ^ port_state_in_8_2_6) ^ port_state_in_11_2_6);
  assign state_out_10_2_6 = (((mul2_106_port_byte_out_6 ^ mul3_106_port_byte_out_6) ^ port_state_in_8_2_6) ^ port_state_in_9_2_6);
  assign state_out_11_2_6 = (((mul2_107_port_byte_out_6 ^ mul3_107_port_byte_out_6) ^ port_state_in_9_2_6) ^ port_state_in_10_2_6);
  assign state_out_8_2_7 = (((mul2_104_port_byte_out_7 ^ mul3_104_port_byte_out_7) ^ port_state_in_10_2_7) ^ port_state_in_11_2_7);
  assign state_out_9_2_7 = (((mul2_105_port_byte_out_7 ^ mul3_105_port_byte_out_7) ^ port_state_in_8_2_7) ^ port_state_in_11_2_7);
  assign state_out_10_2_7 = (((mul2_106_port_byte_out_7 ^ mul3_106_port_byte_out_7) ^ port_state_in_8_2_7) ^ port_state_in_9_2_7);
  assign state_out_11_2_7 = (((mul2_107_port_byte_out_7 ^ mul3_107_port_byte_out_7) ^ port_state_in_9_2_7) ^ port_state_in_10_2_7);
  assign state_out_8_3_0 = (((mul2_108_port_byte_out_0 ^ mul3_108_port_byte_out_0) ^ port_state_in_10_3_0) ^ port_state_in_11_3_0);
  assign state_out_9_3_0 = (((mul2_109_port_byte_out_0 ^ mul3_109_port_byte_out_0) ^ port_state_in_8_3_0) ^ port_state_in_11_3_0);
  assign state_out_10_3_0 = (((mul2_110_port_byte_out_0 ^ mul3_110_port_byte_out_0) ^ port_state_in_8_3_0) ^ port_state_in_9_3_0);
  assign state_out_11_3_0 = (((mul2_111_port_byte_out_0 ^ mul3_111_port_byte_out_0) ^ port_state_in_9_3_0) ^ port_state_in_10_3_0);
  assign state_out_8_3_1 = (((mul2_108_port_byte_out_1 ^ mul3_108_port_byte_out_1) ^ port_state_in_10_3_1) ^ port_state_in_11_3_1);
  assign state_out_9_3_1 = (((mul2_109_port_byte_out_1 ^ mul3_109_port_byte_out_1) ^ port_state_in_8_3_1) ^ port_state_in_11_3_1);
  assign state_out_10_3_1 = (((mul2_110_port_byte_out_1 ^ mul3_110_port_byte_out_1) ^ port_state_in_8_3_1) ^ port_state_in_9_3_1);
  assign state_out_11_3_1 = (((mul2_111_port_byte_out_1 ^ mul3_111_port_byte_out_1) ^ port_state_in_9_3_1) ^ port_state_in_10_3_1);
  assign state_out_8_3_2 = (((mul2_108_port_byte_out_2 ^ mul3_108_port_byte_out_2) ^ port_state_in_10_3_2) ^ port_state_in_11_3_2);
  assign state_out_9_3_2 = (((mul2_109_port_byte_out_2 ^ mul3_109_port_byte_out_2) ^ port_state_in_8_3_2) ^ port_state_in_11_3_2);
  assign state_out_10_3_2 = (((mul2_110_port_byte_out_2 ^ mul3_110_port_byte_out_2) ^ port_state_in_8_3_2) ^ port_state_in_9_3_2);
  assign state_out_11_3_2 = (((mul2_111_port_byte_out_2 ^ mul3_111_port_byte_out_2) ^ port_state_in_9_3_2) ^ port_state_in_10_3_2);
  assign state_out_8_3_3 = (((mul2_108_port_byte_out_3 ^ mul3_108_port_byte_out_3) ^ port_state_in_10_3_3) ^ port_state_in_11_3_3);
  assign state_out_9_3_3 = (((mul2_109_port_byte_out_3 ^ mul3_109_port_byte_out_3) ^ port_state_in_8_3_3) ^ port_state_in_11_3_3);
  assign state_out_10_3_3 = (((mul2_110_port_byte_out_3 ^ mul3_110_port_byte_out_3) ^ port_state_in_8_3_3) ^ port_state_in_9_3_3);
  assign state_out_11_3_3 = (((mul2_111_port_byte_out_3 ^ mul3_111_port_byte_out_3) ^ port_state_in_9_3_3) ^ port_state_in_10_3_3);
  assign state_out_8_3_4 = (((mul2_108_port_byte_out_4 ^ mul3_108_port_byte_out_4) ^ port_state_in_10_3_4) ^ port_state_in_11_3_4);
  assign state_out_9_3_4 = (((mul2_109_port_byte_out_4 ^ mul3_109_port_byte_out_4) ^ port_state_in_8_3_4) ^ port_state_in_11_3_4);
  assign state_out_10_3_4 = (((mul2_110_port_byte_out_4 ^ mul3_110_port_byte_out_4) ^ port_state_in_8_3_4) ^ port_state_in_9_3_4);
  assign state_out_11_3_4 = (((mul2_111_port_byte_out_4 ^ mul3_111_port_byte_out_4) ^ port_state_in_9_3_4) ^ port_state_in_10_3_4);
  assign state_out_8_3_5 = (((mul2_108_port_byte_out_5 ^ mul3_108_port_byte_out_5) ^ port_state_in_10_3_5) ^ port_state_in_11_3_5);
  assign state_out_9_3_5 = (((mul2_109_port_byte_out_5 ^ mul3_109_port_byte_out_5) ^ port_state_in_8_3_5) ^ port_state_in_11_3_5);
  assign state_out_10_3_5 = (((mul2_110_port_byte_out_5 ^ mul3_110_port_byte_out_5) ^ port_state_in_8_3_5) ^ port_state_in_9_3_5);
  assign state_out_11_3_5 = (((mul2_111_port_byte_out_5 ^ mul3_111_port_byte_out_5) ^ port_state_in_9_3_5) ^ port_state_in_10_3_5);
  assign state_out_8_3_6 = (((mul2_108_port_byte_out_6 ^ mul3_108_port_byte_out_6) ^ port_state_in_10_3_6) ^ port_state_in_11_3_6);
  assign state_out_9_3_6 = (((mul2_109_port_byte_out_6 ^ mul3_109_port_byte_out_6) ^ port_state_in_8_3_6) ^ port_state_in_11_3_6);
  assign state_out_10_3_6 = (((mul2_110_port_byte_out_6 ^ mul3_110_port_byte_out_6) ^ port_state_in_8_3_6) ^ port_state_in_9_3_6);
  assign state_out_11_3_6 = (((mul2_111_port_byte_out_6 ^ mul3_111_port_byte_out_6) ^ port_state_in_9_3_6) ^ port_state_in_10_3_6);
  assign state_out_8_3_7 = (((mul2_108_port_byte_out_7 ^ mul3_108_port_byte_out_7) ^ port_state_in_10_3_7) ^ port_state_in_11_3_7);
  assign state_out_9_3_7 = (((mul2_109_port_byte_out_7 ^ mul3_109_port_byte_out_7) ^ port_state_in_8_3_7) ^ port_state_in_11_3_7);
  assign state_out_10_3_7 = (((mul2_110_port_byte_out_7 ^ mul3_110_port_byte_out_7) ^ port_state_in_8_3_7) ^ port_state_in_9_3_7);
  assign state_out_11_3_7 = (((mul2_111_port_byte_out_7 ^ mul3_111_port_byte_out_7) ^ port_state_in_9_3_7) ^ port_state_in_10_3_7);
  assign state_out_12_0_0 = (((mul2_112_port_byte_out_0 ^ mul3_112_port_byte_out_0) ^ port_state_in_14_0_0) ^ port_state_in_15_0_0);
  assign state_out_13_0_0 = (((mul2_113_port_byte_out_0 ^ mul3_113_port_byte_out_0) ^ port_state_in_12_0_0) ^ port_state_in_15_0_0);
  assign state_out_14_0_0 = (((mul2_114_port_byte_out_0 ^ mul3_114_port_byte_out_0) ^ port_state_in_12_0_0) ^ port_state_in_13_0_0);
  assign state_out_15_0_0 = (((mul2_115_port_byte_out_0 ^ mul3_115_port_byte_out_0) ^ port_state_in_13_0_0) ^ port_state_in_14_0_0);
  assign state_out_12_0_1 = (((mul2_112_port_byte_out_1 ^ mul3_112_port_byte_out_1) ^ port_state_in_14_0_1) ^ port_state_in_15_0_1);
  assign state_out_13_0_1 = (((mul2_113_port_byte_out_1 ^ mul3_113_port_byte_out_1) ^ port_state_in_12_0_1) ^ port_state_in_15_0_1);
  assign state_out_14_0_1 = (((mul2_114_port_byte_out_1 ^ mul3_114_port_byte_out_1) ^ port_state_in_12_0_1) ^ port_state_in_13_0_1);
  assign state_out_15_0_1 = (((mul2_115_port_byte_out_1 ^ mul3_115_port_byte_out_1) ^ port_state_in_13_0_1) ^ port_state_in_14_0_1);
  assign state_out_12_0_2 = (((mul2_112_port_byte_out_2 ^ mul3_112_port_byte_out_2) ^ port_state_in_14_0_2) ^ port_state_in_15_0_2);
  assign state_out_13_0_2 = (((mul2_113_port_byte_out_2 ^ mul3_113_port_byte_out_2) ^ port_state_in_12_0_2) ^ port_state_in_15_0_2);
  assign state_out_14_0_2 = (((mul2_114_port_byte_out_2 ^ mul3_114_port_byte_out_2) ^ port_state_in_12_0_2) ^ port_state_in_13_0_2);
  assign state_out_15_0_2 = (((mul2_115_port_byte_out_2 ^ mul3_115_port_byte_out_2) ^ port_state_in_13_0_2) ^ port_state_in_14_0_2);
  assign state_out_12_0_3 = (((mul2_112_port_byte_out_3 ^ mul3_112_port_byte_out_3) ^ port_state_in_14_0_3) ^ port_state_in_15_0_3);
  assign state_out_13_0_3 = (((mul2_113_port_byte_out_3 ^ mul3_113_port_byte_out_3) ^ port_state_in_12_0_3) ^ port_state_in_15_0_3);
  assign state_out_14_0_3 = (((mul2_114_port_byte_out_3 ^ mul3_114_port_byte_out_3) ^ port_state_in_12_0_3) ^ port_state_in_13_0_3);
  assign state_out_15_0_3 = (((mul2_115_port_byte_out_3 ^ mul3_115_port_byte_out_3) ^ port_state_in_13_0_3) ^ port_state_in_14_0_3);
  assign state_out_12_0_4 = (((mul2_112_port_byte_out_4 ^ mul3_112_port_byte_out_4) ^ port_state_in_14_0_4) ^ port_state_in_15_0_4);
  assign state_out_13_0_4 = (((mul2_113_port_byte_out_4 ^ mul3_113_port_byte_out_4) ^ port_state_in_12_0_4) ^ port_state_in_15_0_4);
  assign state_out_14_0_4 = (((mul2_114_port_byte_out_4 ^ mul3_114_port_byte_out_4) ^ port_state_in_12_0_4) ^ port_state_in_13_0_4);
  assign state_out_15_0_4 = (((mul2_115_port_byte_out_4 ^ mul3_115_port_byte_out_4) ^ port_state_in_13_0_4) ^ port_state_in_14_0_4);
  assign state_out_12_0_5 = (((mul2_112_port_byte_out_5 ^ mul3_112_port_byte_out_5) ^ port_state_in_14_0_5) ^ port_state_in_15_0_5);
  assign state_out_13_0_5 = (((mul2_113_port_byte_out_5 ^ mul3_113_port_byte_out_5) ^ port_state_in_12_0_5) ^ port_state_in_15_0_5);
  assign state_out_14_0_5 = (((mul2_114_port_byte_out_5 ^ mul3_114_port_byte_out_5) ^ port_state_in_12_0_5) ^ port_state_in_13_0_5);
  assign state_out_15_0_5 = (((mul2_115_port_byte_out_5 ^ mul3_115_port_byte_out_5) ^ port_state_in_13_0_5) ^ port_state_in_14_0_5);
  assign state_out_12_0_6 = (((mul2_112_port_byte_out_6 ^ mul3_112_port_byte_out_6) ^ port_state_in_14_0_6) ^ port_state_in_15_0_6);
  assign state_out_13_0_6 = (((mul2_113_port_byte_out_6 ^ mul3_113_port_byte_out_6) ^ port_state_in_12_0_6) ^ port_state_in_15_0_6);
  assign state_out_14_0_6 = (((mul2_114_port_byte_out_6 ^ mul3_114_port_byte_out_6) ^ port_state_in_12_0_6) ^ port_state_in_13_0_6);
  assign state_out_15_0_6 = (((mul2_115_port_byte_out_6 ^ mul3_115_port_byte_out_6) ^ port_state_in_13_0_6) ^ port_state_in_14_0_6);
  assign state_out_12_0_7 = (((mul2_112_port_byte_out_7 ^ mul3_112_port_byte_out_7) ^ port_state_in_14_0_7) ^ port_state_in_15_0_7);
  assign state_out_13_0_7 = (((mul2_113_port_byte_out_7 ^ mul3_113_port_byte_out_7) ^ port_state_in_12_0_7) ^ port_state_in_15_0_7);
  assign state_out_14_0_7 = (((mul2_114_port_byte_out_7 ^ mul3_114_port_byte_out_7) ^ port_state_in_12_0_7) ^ port_state_in_13_0_7);
  assign state_out_15_0_7 = (((mul2_115_port_byte_out_7 ^ mul3_115_port_byte_out_7) ^ port_state_in_13_0_7) ^ port_state_in_14_0_7);
  assign state_out_12_1_0 = (((mul2_116_port_byte_out_0 ^ mul3_116_port_byte_out_0) ^ port_state_in_14_1_0) ^ port_state_in_15_1_0);
  assign state_out_13_1_0 = (((mul2_117_port_byte_out_0 ^ mul3_117_port_byte_out_0) ^ port_state_in_12_1_0) ^ port_state_in_15_1_0);
  assign state_out_14_1_0 = (((mul2_118_port_byte_out_0 ^ mul3_118_port_byte_out_0) ^ port_state_in_12_1_0) ^ port_state_in_13_1_0);
  assign state_out_15_1_0 = (((mul2_119_port_byte_out_0 ^ mul3_119_port_byte_out_0) ^ port_state_in_13_1_0) ^ port_state_in_14_1_0);
  assign state_out_12_1_1 = (((mul2_116_port_byte_out_1 ^ mul3_116_port_byte_out_1) ^ port_state_in_14_1_1) ^ port_state_in_15_1_1);
  assign state_out_13_1_1 = (((mul2_117_port_byte_out_1 ^ mul3_117_port_byte_out_1) ^ port_state_in_12_1_1) ^ port_state_in_15_1_1);
  assign state_out_14_1_1 = (((mul2_118_port_byte_out_1 ^ mul3_118_port_byte_out_1) ^ port_state_in_12_1_1) ^ port_state_in_13_1_1);
  assign state_out_15_1_1 = (((mul2_119_port_byte_out_1 ^ mul3_119_port_byte_out_1) ^ port_state_in_13_1_1) ^ port_state_in_14_1_1);
  assign state_out_12_1_2 = (((mul2_116_port_byte_out_2 ^ mul3_116_port_byte_out_2) ^ port_state_in_14_1_2) ^ port_state_in_15_1_2);
  assign state_out_13_1_2 = (((mul2_117_port_byte_out_2 ^ mul3_117_port_byte_out_2) ^ port_state_in_12_1_2) ^ port_state_in_15_1_2);
  assign state_out_14_1_2 = (((mul2_118_port_byte_out_2 ^ mul3_118_port_byte_out_2) ^ port_state_in_12_1_2) ^ port_state_in_13_1_2);
  assign state_out_15_1_2 = (((mul2_119_port_byte_out_2 ^ mul3_119_port_byte_out_2) ^ port_state_in_13_1_2) ^ port_state_in_14_1_2);
  assign state_out_12_1_3 = (((mul2_116_port_byte_out_3 ^ mul3_116_port_byte_out_3) ^ port_state_in_14_1_3) ^ port_state_in_15_1_3);
  assign state_out_13_1_3 = (((mul2_117_port_byte_out_3 ^ mul3_117_port_byte_out_3) ^ port_state_in_12_1_3) ^ port_state_in_15_1_3);
  assign state_out_14_1_3 = (((mul2_118_port_byte_out_3 ^ mul3_118_port_byte_out_3) ^ port_state_in_12_1_3) ^ port_state_in_13_1_3);
  assign state_out_15_1_3 = (((mul2_119_port_byte_out_3 ^ mul3_119_port_byte_out_3) ^ port_state_in_13_1_3) ^ port_state_in_14_1_3);
  assign state_out_12_1_4 = (((mul2_116_port_byte_out_4 ^ mul3_116_port_byte_out_4) ^ port_state_in_14_1_4) ^ port_state_in_15_1_4);
  assign state_out_13_1_4 = (((mul2_117_port_byte_out_4 ^ mul3_117_port_byte_out_4) ^ port_state_in_12_1_4) ^ port_state_in_15_1_4);
  assign state_out_14_1_4 = (((mul2_118_port_byte_out_4 ^ mul3_118_port_byte_out_4) ^ port_state_in_12_1_4) ^ port_state_in_13_1_4);
  assign state_out_15_1_4 = (((mul2_119_port_byte_out_4 ^ mul3_119_port_byte_out_4) ^ port_state_in_13_1_4) ^ port_state_in_14_1_4);
  assign state_out_12_1_5 = (((mul2_116_port_byte_out_5 ^ mul3_116_port_byte_out_5) ^ port_state_in_14_1_5) ^ port_state_in_15_1_5);
  assign state_out_13_1_5 = (((mul2_117_port_byte_out_5 ^ mul3_117_port_byte_out_5) ^ port_state_in_12_1_5) ^ port_state_in_15_1_5);
  assign state_out_14_1_5 = (((mul2_118_port_byte_out_5 ^ mul3_118_port_byte_out_5) ^ port_state_in_12_1_5) ^ port_state_in_13_1_5);
  assign state_out_15_1_5 = (((mul2_119_port_byte_out_5 ^ mul3_119_port_byte_out_5) ^ port_state_in_13_1_5) ^ port_state_in_14_1_5);
  assign state_out_12_1_6 = (((mul2_116_port_byte_out_6 ^ mul3_116_port_byte_out_6) ^ port_state_in_14_1_6) ^ port_state_in_15_1_6);
  assign state_out_13_1_6 = (((mul2_117_port_byte_out_6 ^ mul3_117_port_byte_out_6) ^ port_state_in_12_1_6) ^ port_state_in_15_1_6);
  assign state_out_14_1_6 = (((mul2_118_port_byte_out_6 ^ mul3_118_port_byte_out_6) ^ port_state_in_12_1_6) ^ port_state_in_13_1_6);
  assign state_out_15_1_6 = (((mul2_119_port_byte_out_6 ^ mul3_119_port_byte_out_6) ^ port_state_in_13_1_6) ^ port_state_in_14_1_6);
  assign state_out_12_1_7 = (((mul2_116_port_byte_out_7 ^ mul3_116_port_byte_out_7) ^ port_state_in_14_1_7) ^ port_state_in_15_1_7);
  assign state_out_13_1_7 = (((mul2_117_port_byte_out_7 ^ mul3_117_port_byte_out_7) ^ port_state_in_12_1_7) ^ port_state_in_15_1_7);
  assign state_out_14_1_7 = (((mul2_118_port_byte_out_7 ^ mul3_118_port_byte_out_7) ^ port_state_in_12_1_7) ^ port_state_in_13_1_7);
  assign state_out_15_1_7 = (((mul2_119_port_byte_out_7 ^ mul3_119_port_byte_out_7) ^ port_state_in_13_1_7) ^ port_state_in_14_1_7);
  assign state_out_12_2_0 = (((mul2_120_port_byte_out_0 ^ mul3_120_port_byte_out_0) ^ port_state_in_14_2_0) ^ port_state_in_15_2_0);
  assign state_out_13_2_0 = (((mul2_121_port_byte_out_0 ^ mul3_121_port_byte_out_0) ^ port_state_in_12_2_0) ^ port_state_in_15_2_0);
  assign state_out_14_2_0 = (((mul2_122_port_byte_out_0 ^ mul3_122_port_byte_out_0) ^ port_state_in_12_2_0) ^ port_state_in_13_2_0);
  assign state_out_15_2_0 = (((mul2_123_port_byte_out_0 ^ mul3_123_port_byte_out_0) ^ port_state_in_13_2_0) ^ port_state_in_14_2_0);
  assign state_out_12_2_1 = (((mul2_120_port_byte_out_1 ^ mul3_120_port_byte_out_1) ^ port_state_in_14_2_1) ^ port_state_in_15_2_1);
  assign state_out_13_2_1 = (((mul2_121_port_byte_out_1 ^ mul3_121_port_byte_out_1) ^ port_state_in_12_2_1) ^ port_state_in_15_2_1);
  assign state_out_14_2_1 = (((mul2_122_port_byte_out_1 ^ mul3_122_port_byte_out_1) ^ port_state_in_12_2_1) ^ port_state_in_13_2_1);
  assign state_out_15_2_1 = (((mul2_123_port_byte_out_1 ^ mul3_123_port_byte_out_1) ^ port_state_in_13_2_1) ^ port_state_in_14_2_1);
  assign state_out_12_2_2 = (((mul2_120_port_byte_out_2 ^ mul3_120_port_byte_out_2) ^ port_state_in_14_2_2) ^ port_state_in_15_2_2);
  assign state_out_13_2_2 = (((mul2_121_port_byte_out_2 ^ mul3_121_port_byte_out_2) ^ port_state_in_12_2_2) ^ port_state_in_15_2_2);
  assign state_out_14_2_2 = (((mul2_122_port_byte_out_2 ^ mul3_122_port_byte_out_2) ^ port_state_in_12_2_2) ^ port_state_in_13_2_2);
  assign state_out_15_2_2 = (((mul2_123_port_byte_out_2 ^ mul3_123_port_byte_out_2) ^ port_state_in_13_2_2) ^ port_state_in_14_2_2);
  assign state_out_12_2_3 = (((mul2_120_port_byte_out_3 ^ mul3_120_port_byte_out_3) ^ port_state_in_14_2_3) ^ port_state_in_15_2_3);
  assign state_out_13_2_3 = (((mul2_121_port_byte_out_3 ^ mul3_121_port_byte_out_3) ^ port_state_in_12_2_3) ^ port_state_in_15_2_3);
  assign state_out_14_2_3 = (((mul2_122_port_byte_out_3 ^ mul3_122_port_byte_out_3) ^ port_state_in_12_2_3) ^ port_state_in_13_2_3);
  assign state_out_15_2_3 = (((mul2_123_port_byte_out_3 ^ mul3_123_port_byte_out_3) ^ port_state_in_13_2_3) ^ port_state_in_14_2_3);
  assign state_out_12_2_4 = (((mul2_120_port_byte_out_4 ^ mul3_120_port_byte_out_4) ^ port_state_in_14_2_4) ^ port_state_in_15_2_4);
  assign state_out_13_2_4 = (((mul2_121_port_byte_out_4 ^ mul3_121_port_byte_out_4) ^ port_state_in_12_2_4) ^ port_state_in_15_2_4);
  assign state_out_14_2_4 = (((mul2_122_port_byte_out_4 ^ mul3_122_port_byte_out_4) ^ port_state_in_12_2_4) ^ port_state_in_13_2_4);
  assign state_out_15_2_4 = (((mul2_123_port_byte_out_4 ^ mul3_123_port_byte_out_4) ^ port_state_in_13_2_4) ^ port_state_in_14_2_4);
  assign state_out_12_2_5 = (((mul2_120_port_byte_out_5 ^ mul3_120_port_byte_out_5) ^ port_state_in_14_2_5) ^ port_state_in_15_2_5);
  assign state_out_13_2_5 = (((mul2_121_port_byte_out_5 ^ mul3_121_port_byte_out_5) ^ port_state_in_12_2_5) ^ port_state_in_15_2_5);
  assign state_out_14_2_5 = (((mul2_122_port_byte_out_5 ^ mul3_122_port_byte_out_5) ^ port_state_in_12_2_5) ^ port_state_in_13_2_5);
  assign state_out_15_2_5 = (((mul2_123_port_byte_out_5 ^ mul3_123_port_byte_out_5) ^ port_state_in_13_2_5) ^ port_state_in_14_2_5);
  assign state_out_12_2_6 = (((mul2_120_port_byte_out_6 ^ mul3_120_port_byte_out_6) ^ port_state_in_14_2_6) ^ port_state_in_15_2_6);
  assign state_out_13_2_6 = (((mul2_121_port_byte_out_6 ^ mul3_121_port_byte_out_6) ^ port_state_in_12_2_6) ^ port_state_in_15_2_6);
  assign state_out_14_2_6 = (((mul2_122_port_byte_out_6 ^ mul3_122_port_byte_out_6) ^ port_state_in_12_2_6) ^ port_state_in_13_2_6);
  assign state_out_15_2_6 = (((mul2_123_port_byte_out_6 ^ mul3_123_port_byte_out_6) ^ port_state_in_13_2_6) ^ port_state_in_14_2_6);
  assign state_out_12_2_7 = (((mul2_120_port_byte_out_7 ^ mul3_120_port_byte_out_7) ^ port_state_in_14_2_7) ^ port_state_in_15_2_7);
  assign state_out_13_2_7 = (((mul2_121_port_byte_out_7 ^ mul3_121_port_byte_out_7) ^ port_state_in_12_2_7) ^ port_state_in_15_2_7);
  assign state_out_14_2_7 = (((mul2_122_port_byte_out_7 ^ mul3_122_port_byte_out_7) ^ port_state_in_12_2_7) ^ port_state_in_13_2_7);
  assign state_out_15_2_7 = (((mul2_123_port_byte_out_7 ^ mul3_123_port_byte_out_7) ^ port_state_in_13_2_7) ^ port_state_in_14_2_7);
  assign state_out_12_3_0 = (((mul2_124_port_byte_out_0 ^ mul3_124_port_byte_out_0) ^ port_state_in_14_3_0) ^ port_state_in_15_3_0);
  assign state_out_13_3_0 = (((mul2_125_port_byte_out_0 ^ mul3_125_port_byte_out_0) ^ port_state_in_12_3_0) ^ port_state_in_15_3_0);
  assign state_out_14_3_0 = (((mul2_126_port_byte_out_0 ^ mul3_126_port_byte_out_0) ^ port_state_in_12_3_0) ^ port_state_in_13_3_0);
  assign state_out_15_3_0 = (((mul2_127_port_byte_out_0 ^ mul3_127_port_byte_out_0) ^ port_state_in_13_3_0) ^ port_state_in_14_3_0);
  assign state_out_12_3_1 = (((mul2_124_port_byte_out_1 ^ mul3_124_port_byte_out_1) ^ port_state_in_14_3_1) ^ port_state_in_15_3_1);
  assign state_out_13_3_1 = (((mul2_125_port_byte_out_1 ^ mul3_125_port_byte_out_1) ^ port_state_in_12_3_1) ^ port_state_in_15_3_1);
  assign state_out_14_3_1 = (((mul2_126_port_byte_out_1 ^ mul3_126_port_byte_out_1) ^ port_state_in_12_3_1) ^ port_state_in_13_3_1);
  assign state_out_15_3_1 = (((mul2_127_port_byte_out_1 ^ mul3_127_port_byte_out_1) ^ port_state_in_13_3_1) ^ port_state_in_14_3_1);
  assign state_out_12_3_2 = (((mul2_124_port_byte_out_2 ^ mul3_124_port_byte_out_2) ^ port_state_in_14_3_2) ^ port_state_in_15_3_2);
  assign state_out_13_3_2 = (((mul2_125_port_byte_out_2 ^ mul3_125_port_byte_out_2) ^ port_state_in_12_3_2) ^ port_state_in_15_3_2);
  assign state_out_14_3_2 = (((mul2_126_port_byte_out_2 ^ mul3_126_port_byte_out_2) ^ port_state_in_12_3_2) ^ port_state_in_13_3_2);
  assign state_out_15_3_2 = (((mul2_127_port_byte_out_2 ^ mul3_127_port_byte_out_2) ^ port_state_in_13_3_2) ^ port_state_in_14_3_2);
  assign state_out_12_3_3 = (((mul2_124_port_byte_out_3 ^ mul3_124_port_byte_out_3) ^ port_state_in_14_3_3) ^ port_state_in_15_3_3);
  assign state_out_13_3_3 = (((mul2_125_port_byte_out_3 ^ mul3_125_port_byte_out_3) ^ port_state_in_12_3_3) ^ port_state_in_15_3_3);
  assign state_out_14_3_3 = (((mul2_126_port_byte_out_3 ^ mul3_126_port_byte_out_3) ^ port_state_in_12_3_3) ^ port_state_in_13_3_3);
  assign state_out_15_3_3 = (((mul2_127_port_byte_out_3 ^ mul3_127_port_byte_out_3) ^ port_state_in_13_3_3) ^ port_state_in_14_3_3);
  assign state_out_12_3_4 = (((mul2_124_port_byte_out_4 ^ mul3_124_port_byte_out_4) ^ port_state_in_14_3_4) ^ port_state_in_15_3_4);
  assign state_out_13_3_4 = (((mul2_125_port_byte_out_4 ^ mul3_125_port_byte_out_4) ^ port_state_in_12_3_4) ^ port_state_in_15_3_4);
  assign state_out_14_3_4 = (((mul2_126_port_byte_out_4 ^ mul3_126_port_byte_out_4) ^ port_state_in_12_3_4) ^ port_state_in_13_3_4);
  assign state_out_15_3_4 = (((mul2_127_port_byte_out_4 ^ mul3_127_port_byte_out_4) ^ port_state_in_13_3_4) ^ port_state_in_14_3_4);
  assign state_out_12_3_5 = (((mul2_124_port_byte_out_5 ^ mul3_124_port_byte_out_5) ^ port_state_in_14_3_5) ^ port_state_in_15_3_5);
  assign state_out_13_3_5 = (((mul2_125_port_byte_out_5 ^ mul3_125_port_byte_out_5) ^ port_state_in_12_3_5) ^ port_state_in_15_3_5);
  assign state_out_14_3_5 = (((mul2_126_port_byte_out_5 ^ mul3_126_port_byte_out_5) ^ port_state_in_12_3_5) ^ port_state_in_13_3_5);
  assign state_out_15_3_5 = (((mul2_127_port_byte_out_5 ^ mul3_127_port_byte_out_5) ^ port_state_in_13_3_5) ^ port_state_in_14_3_5);
  assign state_out_12_3_6 = (((mul2_124_port_byte_out_6 ^ mul3_124_port_byte_out_6) ^ port_state_in_14_3_6) ^ port_state_in_15_3_6);
  assign state_out_13_3_6 = (((mul2_125_port_byte_out_6 ^ mul3_125_port_byte_out_6) ^ port_state_in_12_3_6) ^ port_state_in_15_3_6);
  assign state_out_14_3_6 = (((mul2_126_port_byte_out_6 ^ mul3_126_port_byte_out_6) ^ port_state_in_12_3_6) ^ port_state_in_13_3_6);
  assign state_out_15_3_6 = (((mul2_127_port_byte_out_6 ^ mul3_127_port_byte_out_6) ^ port_state_in_13_3_6) ^ port_state_in_14_3_6);
  assign state_out_12_3_7 = (((mul2_124_port_byte_out_7 ^ mul3_124_port_byte_out_7) ^ port_state_in_14_3_7) ^ port_state_in_15_3_7);
  assign state_out_13_3_7 = (((mul2_125_port_byte_out_7 ^ mul3_125_port_byte_out_7) ^ port_state_in_12_3_7) ^ port_state_in_15_3_7);
  assign state_out_14_3_7 = (((mul2_126_port_byte_out_7 ^ mul3_126_port_byte_out_7) ^ port_state_in_12_3_7) ^ port_state_in_13_3_7);
  assign state_out_15_3_7 = (((mul2_127_port_byte_out_7 ^ mul3_127_port_byte_out_7) ^ port_state_in_13_3_7) ^ port_state_in_14_3_7);
  assign port_state_out_0_0_0 = state_out_0_0_0;
  assign port_state_out_0_0_1 = state_out_0_0_1;
  assign port_state_out_0_0_2 = state_out_0_0_2;
  assign port_state_out_0_0_3 = state_out_0_0_3;
  assign port_state_out_0_0_4 = state_out_0_0_4;
  assign port_state_out_0_0_5 = state_out_0_0_5;
  assign port_state_out_0_0_6 = state_out_0_0_6;
  assign port_state_out_0_0_7 = state_out_0_0_7;
  assign port_state_out_0_1_0 = state_out_0_1_0;
  assign port_state_out_0_1_1 = state_out_0_1_1;
  assign port_state_out_0_1_2 = state_out_0_1_2;
  assign port_state_out_0_1_3 = state_out_0_1_3;
  assign port_state_out_0_1_4 = state_out_0_1_4;
  assign port_state_out_0_1_5 = state_out_0_1_5;
  assign port_state_out_0_1_6 = state_out_0_1_6;
  assign port_state_out_0_1_7 = state_out_0_1_7;
  assign port_state_out_0_2_0 = state_out_0_2_0;
  assign port_state_out_0_2_1 = state_out_0_2_1;
  assign port_state_out_0_2_2 = state_out_0_2_2;
  assign port_state_out_0_2_3 = state_out_0_2_3;
  assign port_state_out_0_2_4 = state_out_0_2_4;
  assign port_state_out_0_2_5 = state_out_0_2_5;
  assign port_state_out_0_2_6 = state_out_0_2_6;
  assign port_state_out_0_2_7 = state_out_0_2_7;
  assign port_state_out_0_3_0 = state_out_0_3_0;
  assign port_state_out_0_3_1 = state_out_0_3_1;
  assign port_state_out_0_3_2 = state_out_0_3_2;
  assign port_state_out_0_3_3 = state_out_0_3_3;
  assign port_state_out_0_3_4 = state_out_0_3_4;
  assign port_state_out_0_3_5 = state_out_0_3_5;
  assign port_state_out_0_3_6 = state_out_0_3_6;
  assign port_state_out_0_3_7 = state_out_0_3_7;
  assign port_state_out_1_0_0 = state_out_1_0_0;
  assign port_state_out_1_0_1 = state_out_1_0_1;
  assign port_state_out_1_0_2 = state_out_1_0_2;
  assign port_state_out_1_0_3 = state_out_1_0_3;
  assign port_state_out_1_0_4 = state_out_1_0_4;
  assign port_state_out_1_0_5 = state_out_1_0_5;
  assign port_state_out_1_0_6 = state_out_1_0_6;
  assign port_state_out_1_0_7 = state_out_1_0_7;
  assign port_state_out_1_1_0 = state_out_1_1_0;
  assign port_state_out_1_1_1 = state_out_1_1_1;
  assign port_state_out_1_1_2 = state_out_1_1_2;
  assign port_state_out_1_1_3 = state_out_1_1_3;
  assign port_state_out_1_1_4 = state_out_1_1_4;
  assign port_state_out_1_1_5 = state_out_1_1_5;
  assign port_state_out_1_1_6 = state_out_1_1_6;
  assign port_state_out_1_1_7 = state_out_1_1_7;
  assign port_state_out_1_2_0 = state_out_1_2_0;
  assign port_state_out_1_2_1 = state_out_1_2_1;
  assign port_state_out_1_2_2 = state_out_1_2_2;
  assign port_state_out_1_2_3 = state_out_1_2_3;
  assign port_state_out_1_2_4 = state_out_1_2_4;
  assign port_state_out_1_2_5 = state_out_1_2_5;
  assign port_state_out_1_2_6 = state_out_1_2_6;
  assign port_state_out_1_2_7 = state_out_1_2_7;
  assign port_state_out_1_3_0 = state_out_1_3_0;
  assign port_state_out_1_3_1 = state_out_1_3_1;
  assign port_state_out_1_3_2 = state_out_1_3_2;
  assign port_state_out_1_3_3 = state_out_1_3_3;
  assign port_state_out_1_3_4 = state_out_1_3_4;
  assign port_state_out_1_3_5 = state_out_1_3_5;
  assign port_state_out_1_3_6 = state_out_1_3_6;
  assign port_state_out_1_3_7 = state_out_1_3_7;
  assign port_state_out_2_0_0 = state_out_2_0_0;
  assign port_state_out_2_0_1 = state_out_2_0_1;
  assign port_state_out_2_0_2 = state_out_2_0_2;
  assign port_state_out_2_0_3 = state_out_2_0_3;
  assign port_state_out_2_0_4 = state_out_2_0_4;
  assign port_state_out_2_0_5 = state_out_2_0_5;
  assign port_state_out_2_0_6 = state_out_2_0_6;
  assign port_state_out_2_0_7 = state_out_2_0_7;
  assign port_state_out_2_1_0 = state_out_2_1_0;
  assign port_state_out_2_1_1 = state_out_2_1_1;
  assign port_state_out_2_1_2 = state_out_2_1_2;
  assign port_state_out_2_1_3 = state_out_2_1_3;
  assign port_state_out_2_1_4 = state_out_2_1_4;
  assign port_state_out_2_1_5 = state_out_2_1_5;
  assign port_state_out_2_1_6 = state_out_2_1_6;
  assign port_state_out_2_1_7 = state_out_2_1_7;
  assign port_state_out_2_2_0 = state_out_2_2_0;
  assign port_state_out_2_2_1 = state_out_2_2_1;
  assign port_state_out_2_2_2 = state_out_2_2_2;
  assign port_state_out_2_2_3 = state_out_2_2_3;
  assign port_state_out_2_2_4 = state_out_2_2_4;
  assign port_state_out_2_2_5 = state_out_2_2_5;
  assign port_state_out_2_2_6 = state_out_2_2_6;
  assign port_state_out_2_2_7 = state_out_2_2_7;
  assign port_state_out_2_3_0 = state_out_2_3_0;
  assign port_state_out_2_3_1 = state_out_2_3_1;
  assign port_state_out_2_3_2 = state_out_2_3_2;
  assign port_state_out_2_3_3 = state_out_2_3_3;
  assign port_state_out_2_3_4 = state_out_2_3_4;
  assign port_state_out_2_3_5 = state_out_2_3_5;
  assign port_state_out_2_3_6 = state_out_2_3_6;
  assign port_state_out_2_3_7 = state_out_2_3_7;
  assign port_state_out_3_0_0 = state_out_3_0_0;
  assign port_state_out_3_0_1 = state_out_3_0_1;
  assign port_state_out_3_0_2 = state_out_3_0_2;
  assign port_state_out_3_0_3 = state_out_3_0_3;
  assign port_state_out_3_0_4 = state_out_3_0_4;
  assign port_state_out_3_0_5 = state_out_3_0_5;
  assign port_state_out_3_0_6 = state_out_3_0_6;
  assign port_state_out_3_0_7 = state_out_3_0_7;
  assign port_state_out_3_1_0 = state_out_3_1_0;
  assign port_state_out_3_1_1 = state_out_3_1_1;
  assign port_state_out_3_1_2 = state_out_3_1_2;
  assign port_state_out_3_1_3 = state_out_3_1_3;
  assign port_state_out_3_1_4 = state_out_3_1_4;
  assign port_state_out_3_1_5 = state_out_3_1_5;
  assign port_state_out_3_1_6 = state_out_3_1_6;
  assign port_state_out_3_1_7 = state_out_3_1_7;
  assign port_state_out_3_2_0 = state_out_3_2_0;
  assign port_state_out_3_2_1 = state_out_3_2_1;
  assign port_state_out_3_2_2 = state_out_3_2_2;
  assign port_state_out_3_2_3 = state_out_3_2_3;
  assign port_state_out_3_2_4 = state_out_3_2_4;
  assign port_state_out_3_2_5 = state_out_3_2_5;
  assign port_state_out_3_2_6 = state_out_3_2_6;
  assign port_state_out_3_2_7 = state_out_3_2_7;
  assign port_state_out_3_3_0 = state_out_3_3_0;
  assign port_state_out_3_3_1 = state_out_3_3_1;
  assign port_state_out_3_3_2 = state_out_3_3_2;
  assign port_state_out_3_3_3 = state_out_3_3_3;
  assign port_state_out_3_3_4 = state_out_3_3_4;
  assign port_state_out_3_3_5 = state_out_3_3_5;
  assign port_state_out_3_3_6 = state_out_3_3_6;
  assign port_state_out_3_3_7 = state_out_3_3_7;
  assign port_state_out_4_0_0 = state_out_4_0_0;
  assign port_state_out_4_0_1 = state_out_4_0_1;
  assign port_state_out_4_0_2 = state_out_4_0_2;
  assign port_state_out_4_0_3 = state_out_4_0_3;
  assign port_state_out_4_0_4 = state_out_4_0_4;
  assign port_state_out_4_0_5 = state_out_4_0_5;
  assign port_state_out_4_0_6 = state_out_4_0_6;
  assign port_state_out_4_0_7 = state_out_4_0_7;
  assign port_state_out_4_1_0 = state_out_4_1_0;
  assign port_state_out_4_1_1 = state_out_4_1_1;
  assign port_state_out_4_1_2 = state_out_4_1_2;
  assign port_state_out_4_1_3 = state_out_4_1_3;
  assign port_state_out_4_1_4 = state_out_4_1_4;
  assign port_state_out_4_1_5 = state_out_4_1_5;
  assign port_state_out_4_1_6 = state_out_4_1_6;
  assign port_state_out_4_1_7 = state_out_4_1_7;
  assign port_state_out_4_2_0 = state_out_4_2_0;
  assign port_state_out_4_2_1 = state_out_4_2_1;
  assign port_state_out_4_2_2 = state_out_4_2_2;
  assign port_state_out_4_2_3 = state_out_4_2_3;
  assign port_state_out_4_2_4 = state_out_4_2_4;
  assign port_state_out_4_2_5 = state_out_4_2_5;
  assign port_state_out_4_2_6 = state_out_4_2_6;
  assign port_state_out_4_2_7 = state_out_4_2_7;
  assign port_state_out_4_3_0 = state_out_4_3_0;
  assign port_state_out_4_3_1 = state_out_4_3_1;
  assign port_state_out_4_3_2 = state_out_4_3_2;
  assign port_state_out_4_3_3 = state_out_4_3_3;
  assign port_state_out_4_3_4 = state_out_4_3_4;
  assign port_state_out_4_3_5 = state_out_4_3_5;
  assign port_state_out_4_3_6 = state_out_4_3_6;
  assign port_state_out_4_3_7 = state_out_4_3_7;
  assign port_state_out_5_0_0 = state_out_5_0_0;
  assign port_state_out_5_0_1 = state_out_5_0_1;
  assign port_state_out_5_0_2 = state_out_5_0_2;
  assign port_state_out_5_0_3 = state_out_5_0_3;
  assign port_state_out_5_0_4 = state_out_5_0_4;
  assign port_state_out_5_0_5 = state_out_5_0_5;
  assign port_state_out_5_0_6 = state_out_5_0_6;
  assign port_state_out_5_0_7 = state_out_5_0_7;
  assign port_state_out_5_1_0 = state_out_5_1_0;
  assign port_state_out_5_1_1 = state_out_5_1_1;
  assign port_state_out_5_1_2 = state_out_5_1_2;
  assign port_state_out_5_1_3 = state_out_5_1_3;
  assign port_state_out_5_1_4 = state_out_5_1_4;
  assign port_state_out_5_1_5 = state_out_5_1_5;
  assign port_state_out_5_1_6 = state_out_5_1_6;
  assign port_state_out_5_1_7 = state_out_5_1_7;
  assign port_state_out_5_2_0 = state_out_5_2_0;
  assign port_state_out_5_2_1 = state_out_5_2_1;
  assign port_state_out_5_2_2 = state_out_5_2_2;
  assign port_state_out_5_2_3 = state_out_5_2_3;
  assign port_state_out_5_2_4 = state_out_5_2_4;
  assign port_state_out_5_2_5 = state_out_5_2_5;
  assign port_state_out_5_2_6 = state_out_5_2_6;
  assign port_state_out_5_2_7 = state_out_5_2_7;
  assign port_state_out_5_3_0 = state_out_5_3_0;
  assign port_state_out_5_3_1 = state_out_5_3_1;
  assign port_state_out_5_3_2 = state_out_5_3_2;
  assign port_state_out_5_3_3 = state_out_5_3_3;
  assign port_state_out_5_3_4 = state_out_5_3_4;
  assign port_state_out_5_3_5 = state_out_5_3_5;
  assign port_state_out_5_3_6 = state_out_5_3_6;
  assign port_state_out_5_3_7 = state_out_5_3_7;
  assign port_state_out_6_0_0 = state_out_6_0_0;
  assign port_state_out_6_0_1 = state_out_6_0_1;
  assign port_state_out_6_0_2 = state_out_6_0_2;
  assign port_state_out_6_0_3 = state_out_6_0_3;
  assign port_state_out_6_0_4 = state_out_6_0_4;
  assign port_state_out_6_0_5 = state_out_6_0_5;
  assign port_state_out_6_0_6 = state_out_6_0_6;
  assign port_state_out_6_0_7 = state_out_6_0_7;
  assign port_state_out_6_1_0 = state_out_6_1_0;
  assign port_state_out_6_1_1 = state_out_6_1_1;
  assign port_state_out_6_1_2 = state_out_6_1_2;
  assign port_state_out_6_1_3 = state_out_6_1_3;
  assign port_state_out_6_1_4 = state_out_6_1_4;
  assign port_state_out_6_1_5 = state_out_6_1_5;
  assign port_state_out_6_1_6 = state_out_6_1_6;
  assign port_state_out_6_1_7 = state_out_6_1_7;
  assign port_state_out_6_2_0 = state_out_6_2_0;
  assign port_state_out_6_2_1 = state_out_6_2_1;
  assign port_state_out_6_2_2 = state_out_6_2_2;
  assign port_state_out_6_2_3 = state_out_6_2_3;
  assign port_state_out_6_2_4 = state_out_6_2_4;
  assign port_state_out_6_2_5 = state_out_6_2_5;
  assign port_state_out_6_2_6 = state_out_6_2_6;
  assign port_state_out_6_2_7 = state_out_6_2_7;
  assign port_state_out_6_3_0 = state_out_6_3_0;
  assign port_state_out_6_3_1 = state_out_6_3_1;
  assign port_state_out_6_3_2 = state_out_6_3_2;
  assign port_state_out_6_3_3 = state_out_6_3_3;
  assign port_state_out_6_3_4 = state_out_6_3_4;
  assign port_state_out_6_3_5 = state_out_6_3_5;
  assign port_state_out_6_3_6 = state_out_6_3_6;
  assign port_state_out_6_3_7 = state_out_6_3_7;
  assign port_state_out_7_0_0 = state_out_7_0_0;
  assign port_state_out_7_0_1 = state_out_7_0_1;
  assign port_state_out_7_0_2 = state_out_7_0_2;
  assign port_state_out_7_0_3 = state_out_7_0_3;
  assign port_state_out_7_0_4 = state_out_7_0_4;
  assign port_state_out_7_0_5 = state_out_7_0_5;
  assign port_state_out_7_0_6 = state_out_7_0_6;
  assign port_state_out_7_0_7 = state_out_7_0_7;
  assign port_state_out_7_1_0 = state_out_7_1_0;
  assign port_state_out_7_1_1 = state_out_7_1_1;
  assign port_state_out_7_1_2 = state_out_7_1_2;
  assign port_state_out_7_1_3 = state_out_7_1_3;
  assign port_state_out_7_1_4 = state_out_7_1_4;
  assign port_state_out_7_1_5 = state_out_7_1_5;
  assign port_state_out_7_1_6 = state_out_7_1_6;
  assign port_state_out_7_1_7 = state_out_7_1_7;
  assign port_state_out_7_2_0 = state_out_7_2_0;
  assign port_state_out_7_2_1 = state_out_7_2_1;
  assign port_state_out_7_2_2 = state_out_7_2_2;
  assign port_state_out_7_2_3 = state_out_7_2_3;
  assign port_state_out_7_2_4 = state_out_7_2_4;
  assign port_state_out_7_2_5 = state_out_7_2_5;
  assign port_state_out_7_2_6 = state_out_7_2_6;
  assign port_state_out_7_2_7 = state_out_7_2_7;
  assign port_state_out_7_3_0 = state_out_7_3_0;
  assign port_state_out_7_3_1 = state_out_7_3_1;
  assign port_state_out_7_3_2 = state_out_7_3_2;
  assign port_state_out_7_3_3 = state_out_7_3_3;
  assign port_state_out_7_3_4 = state_out_7_3_4;
  assign port_state_out_7_3_5 = state_out_7_3_5;
  assign port_state_out_7_3_6 = state_out_7_3_6;
  assign port_state_out_7_3_7 = state_out_7_3_7;
  assign port_state_out_8_0_0 = state_out_8_0_0;
  assign port_state_out_8_0_1 = state_out_8_0_1;
  assign port_state_out_8_0_2 = state_out_8_0_2;
  assign port_state_out_8_0_3 = state_out_8_0_3;
  assign port_state_out_8_0_4 = state_out_8_0_4;
  assign port_state_out_8_0_5 = state_out_8_0_5;
  assign port_state_out_8_0_6 = state_out_8_0_6;
  assign port_state_out_8_0_7 = state_out_8_0_7;
  assign port_state_out_8_1_0 = state_out_8_1_0;
  assign port_state_out_8_1_1 = state_out_8_1_1;
  assign port_state_out_8_1_2 = state_out_8_1_2;
  assign port_state_out_8_1_3 = state_out_8_1_3;
  assign port_state_out_8_1_4 = state_out_8_1_4;
  assign port_state_out_8_1_5 = state_out_8_1_5;
  assign port_state_out_8_1_6 = state_out_8_1_6;
  assign port_state_out_8_1_7 = state_out_8_1_7;
  assign port_state_out_8_2_0 = state_out_8_2_0;
  assign port_state_out_8_2_1 = state_out_8_2_1;
  assign port_state_out_8_2_2 = state_out_8_2_2;
  assign port_state_out_8_2_3 = state_out_8_2_3;
  assign port_state_out_8_2_4 = state_out_8_2_4;
  assign port_state_out_8_2_5 = state_out_8_2_5;
  assign port_state_out_8_2_6 = state_out_8_2_6;
  assign port_state_out_8_2_7 = state_out_8_2_7;
  assign port_state_out_8_3_0 = state_out_8_3_0;
  assign port_state_out_8_3_1 = state_out_8_3_1;
  assign port_state_out_8_3_2 = state_out_8_3_2;
  assign port_state_out_8_3_3 = state_out_8_3_3;
  assign port_state_out_8_3_4 = state_out_8_3_4;
  assign port_state_out_8_3_5 = state_out_8_3_5;
  assign port_state_out_8_3_6 = state_out_8_3_6;
  assign port_state_out_8_3_7 = state_out_8_3_7;
  assign port_state_out_9_0_0 = state_out_9_0_0;
  assign port_state_out_9_0_1 = state_out_9_0_1;
  assign port_state_out_9_0_2 = state_out_9_0_2;
  assign port_state_out_9_0_3 = state_out_9_0_3;
  assign port_state_out_9_0_4 = state_out_9_0_4;
  assign port_state_out_9_0_5 = state_out_9_0_5;
  assign port_state_out_9_0_6 = state_out_9_0_6;
  assign port_state_out_9_0_7 = state_out_9_0_7;
  assign port_state_out_9_1_0 = state_out_9_1_0;
  assign port_state_out_9_1_1 = state_out_9_1_1;
  assign port_state_out_9_1_2 = state_out_9_1_2;
  assign port_state_out_9_1_3 = state_out_9_1_3;
  assign port_state_out_9_1_4 = state_out_9_1_4;
  assign port_state_out_9_1_5 = state_out_9_1_5;
  assign port_state_out_9_1_6 = state_out_9_1_6;
  assign port_state_out_9_1_7 = state_out_9_1_7;
  assign port_state_out_9_2_0 = state_out_9_2_0;
  assign port_state_out_9_2_1 = state_out_9_2_1;
  assign port_state_out_9_2_2 = state_out_9_2_2;
  assign port_state_out_9_2_3 = state_out_9_2_3;
  assign port_state_out_9_2_4 = state_out_9_2_4;
  assign port_state_out_9_2_5 = state_out_9_2_5;
  assign port_state_out_9_2_6 = state_out_9_2_6;
  assign port_state_out_9_2_7 = state_out_9_2_7;
  assign port_state_out_9_3_0 = state_out_9_3_0;
  assign port_state_out_9_3_1 = state_out_9_3_1;
  assign port_state_out_9_3_2 = state_out_9_3_2;
  assign port_state_out_9_3_3 = state_out_9_3_3;
  assign port_state_out_9_3_4 = state_out_9_3_4;
  assign port_state_out_9_3_5 = state_out_9_3_5;
  assign port_state_out_9_3_6 = state_out_9_3_6;
  assign port_state_out_9_3_7 = state_out_9_3_7;
  assign port_state_out_10_0_0 = state_out_10_0_0;
  assign port_state_out_10_0_1 = state_out_10_0_1;
  assign port_state_out_10_0_2 = state_out_10_0_2;
  assign port_state_out_10_0_3 = state_out_10_0_3;
  assign port_state_out_10_0_4 = state_out_10_0_4;
  assign port_state_out_10_0_5 = state_out_10_0_5;
  assign port_state_out_10_0_6 = state_out_10_0_6;
  assign port_state_out_10_0_7 = state_out_10_0_7;
  assign port_state_out_10_1_0 = state_out_10_1_0;
  assign port_state_out_10_1_1 = state_out_10_1_1;
  assign port_state_out_10_1_2 = state_out_10_1_2;
  assign port_state_out_10_1_3 = state_out_10_1_3;
  assign port_state_out_10_1_4 = state_out_10_1_4;
  assign port_state_out_10_1_5 = state_out_10_1_5;
  assign port_state_out_10_1_6 = state_out_10_1_6;
  assign port_state_out_10_1_7 = state_out_10_1_7;
  assign port_state_out_10_2_0 = state_out_10_2_0;
  assign port_state_out_10_2_1 = state_out_10_2_1;
  assign port_state_out_10_2_2 = state_out_10_2_2;
  assign port_state_out_10_2_3 = state_out_10_2_3;
  assign port_state_out_10_2_4 = state_out_10_2_4;
  assign port_state_out_10_2_5 = state_out_10_2_5;
  assign port_state_out_10_2_6 = state_out_10_2_6;
  assign port_state_out_10_2_7 = state_out_10_2_7;
  assign port_state_out_10_3_0 = state_out_10_3_0;
  assign port_state_out_10_3_1 = state_out_10_3_1;
  assign port_state_out_10_3_2 = state_out_10_3_2;
  assign port_state_out_10_3_3 = state_out_10_3_3;
  assign port_state_out_10_3_4 = state_out_10_3_4;
  assign port_state_out_10_3_5 = state_out_10_3_5;
  assign port_state_out_10_3_6 = state_out_10_3_6;
  assign port_state_out_10_3_7 = state_out_10_3_7;
  assign port_state_out_11_0_0 = state_out_11_0_0;
  assign port_state_out_11_0_1 = state_out_11_0_1;
  assign port_state_out_11_0_2 = state_out_11_0_2;
  assign port_state_out_11_0_3 = state_out_11_0_3;
  assign port_state_out_11_0_4 = state_out_11_0_4;
  assign port_state_out_11_0_5 = state_out_11_0_5;
  assign port_state_out_11_0_6 = state_out_11_0_6;
  assign port_state_out_11_0_7 = state_out_11_0_7;
  assign port_state_out_11_1_0 = state_out_11_1_0;
  assign port_state_out_11_1_1 = state_out_11_1_1;
  assign port_state_out_11_1_2 = state_out_11_1_2;
  assign port_state_out_11_1_3 = state_out_11_1_3;
  assign port_state_out_11_1_4 = state_out_11_1_4;
  assign port_state_out_11_1_5 = state_out_11_1_5;
  assign port_state_out_11_1_6 = state_out_11_1_6;
  assign port_state_out_11_1_7 = state_out_11_1_7;
  assign port_state_out_11_2_0 = state_out_11_2_0;
  assign port_state_out_11_2_1 = state_out_11_2_1;
  assign port_state_out_11_2_2 = state_out_11_2_2;
  assign port_state_out_11_2_3 = state_out_11_2_3;
  assign port_state_out_11_2_4 = state_out_11_2_4;
  assign port_state_out_11_2_5 = state_out_11_2_5;
  assign port_state_out_11_2_6 = state_out_11_2_6;
  assign port_state_out_11_2_7 = state_out_11_2_7;
  assign port_state_out_11_3_0 = state_out_11_3_0;
  assign port_state_out_11_3_1 = state_out_11_3_1;
  assign port_state_out_11_3_2 = state_out_11_3_2;
  assign port_state_out_11_3_3 = state_out_11_3_3;
  assign port_state_out_11_3_4 = state_out_11_3_4;
  assign port_state_out_11_3_5 = state_out_11_3_5;
  assign port_state_out_11_3_6 = state_out_11_3_6;
  assign port_state_out_11_3_7 = state_out_11_3_7;
  assign port_state_out_12_0_0 = state_out_12_0_0;
  assign port_state_out_12_0_1 = state_out_12_0_1;
  assign port_state_out_12_0_2 = state_out_12_0_2;
  assign port_state_out_12_0_3 = state_out_12_0_3;
  assign port_state_out_12_0_4 = state_out_12_0_4;
  assign port_state_out_12_0_5 = state_out_12_0_5;
  assign port_state_out_12_0_6 = state_out_12_0_6;
  assign port_state_out_12_0_7 = state_out_12_0_7;
  assign port_state_out_12_1_0 = state_out_12_1_0;
  assign port_state_out_12_1_1 = state_out_12_1_1;
  assign port_state_out_12_1_2 = state_out_12_1_2;
  assign port_state_out_12_1_3 = state_out_12_1_3;
  assign port_state_out_12_1_4 = state_out_12_1_4;
  assign port_state_out_12_1_5 = state_out_12_1_5;
  assign port_state_out_12_1_6 = state_out_12_1_6;
  assign port_state_out_12_1_7 = state_out_12_1_7;
  assign port_state_out_12_2_0 = state_out_12_2_0;
  assign port_state_out_12_2_1 = state_out_12_2_1;
  assign port_state_out_12_2_2 = state_out_12_2_2;
  assign port_state_out_12_2_3 = state_out_12_2_3;
  assign port_state_out_12_2_4 = state_out_12_2_4;
  assign port_state_out_12_2_5 = state_out_12_2_5;
  assign port_state_out_12_2_6 = state_out_12_2_6;
  assign port_state_out_12_2_7 = state_out_12_2_7;
  assign port_state_out_12_3_0 = state_out_12_3_0;
  assign port_state_out_12_3_1 = state_out_12_3_1;
  assign port_state_out_12_3_2 = state_out_12_3_2;
  assign port_state_out_12_3_3 = state_out_12_3_3;
  assign port_state_out_12_3_4 = state_out_12_3_4;
  assign port_state_out_12_3_5 = state_out_12_3_5;
  assign port_state_out_12_3_6 = state_out_12_3_6;
  assign port_state_out_12_3_7 = state_out_12_3_7;
  assign port_state_out_13_0_0 = state_out_13_0_0;
  assign port_state_out_13_0_1 = state_out_13_0_1;
  assign port_state_out_13_0_2 = state_out_13_0_2;
  assign port_state_out_13_0_3 = state_out_13_0_3;
  assign port_state_out_13_0_4 = state_out_13_0_4;
  assign port_state_out_13_0_5 = state_out_13_0_5;
  assign port_state_out_13_0_6 = state_out_13_0_6;
  assign port_state_out_13_0_7 = state_out_13_0_7;
  assign port_state_out_13_1_0 = state_out_13_1_0;
  assign port_state_out_13_1_1 = state_out_13_1_1;
  assign port_state_out_13_1_2 = state_out_13_1_2;
  assign port_state_out_13_1_3 = state_out_13_1_3;
  assign port_state_out_13_1_4 = state_out_13_1_4;
  assign port_state_out_13_1_5 = state_out_13_1_5;
  assign port_state_out_13_1_6 = state_out_13_1_6;
  assign port_state_out_13_1_7 = state_out_13_1_7;
  assign port_state_out_13_2_0 = state_out_13_2_0;
  assign port_state_out_13_2_1 = state_out_13_2_1;
  assign port_state_out_13_2_2 = state_out_13_2_2;
  assign port_state_out_13_2_3 = state_out_13_2_3;
  assign port_state_out_13_2_4 = state_out_13_2_4;
  assign port_state_out_13_2_5 = state_out_13_2_5;
  assign port_state_out_13_2_6 = state_out_13_2_6;
  assign port_state_out_13_2_7 = state_out_13_2_7;
  assign port_state_out_13_3_0 = state_out_13_3_0;
  assign port_state_out_13_3_1 = state_out_13_3_1;
  assign port_state_out_13_3_2 = state_out_13_3_2;
  assign port_state_out_13_3_3 = state_out_13_3_3;
  assign port_state_out_13_3_4 = state_out_13_3_4;
  assign port_state_out_13_3_5 = state_out_13_3_5;
  assign port_state_out_13_3_6 = state_out_13_3_6;
  assign port_state_out_13_3_7 = state_out_13_3_7;
  assign port_state_out_14_0_0 = state_out_14_0_0;
  assign port_state_out_14_0_1 = state_out_14_0_1;
  assign port_state_out_14_0_2 = state_out_14_0_2;
  assign port_state_out_14_0_3 = state_out_14_0_3;
  assign port_state_out_14_0_4 = state_out_14_0_4;
  assign port_state_out_14_0_5 = state_out_14_0_5;
  assign port_state_out_14_0_6 = state_out_14_0_6;
  assign port_state_out_14_0_7 = state_out_14_0_7;
  assign port_state_out_14_1_0 = state_out_14_1_0;
  assign port_state_out_14_1_1 = state_out_14_1_1;
  assign port_state_out_14_1_2 = state_out_14_1_2;
  assign port_state_out_14_1_3 = state_out_14_1_3;
  assign port_state_out_14_1_4 = state_out_14_1_4;
  assign port_state_out_14_1_5 = state_out_14_1_5;
  assign port_state_out_14_1_6 = state_out_14_1_6;
  assign port_state_out_14_1_7 = state_out_14_1_7;
  assign port_state_out_14_2_0 = state_out_14_2_0;
  assign port_state_out_14_2_1 = state_out_14_2_1;
  assign port_state_out_14_2_2 = state_out_14_2_2;
  assign port_state_out_14_2_3 = state_out_14_2_3;
  assign port_state_out_14_2_4 = state_out_14_2_4;
  assign port_state_out_14_2_5 = state_out_14_2_5;
  assign port_state_out_14_2_6 = state_out_14_2_6;
  assign port_state_out_14_2_7 = state_out_14_2_7;
  assign port_state_out_14_3_0 = state_out_14_3_0;
  assign port_state_out_14_3_1 = state_out_14_3_1;
  assign port_state_out_14_3_2 = state_out_14_3_2;
  assign port_state_out_14_3_3 = state_out_14_3_3;
  assign port_state_out_14_3_4 = state_out_14_3_4;
  assign port_state_out_14_3_5 = state_out_14_3_5;
  assign port_state_out_14_3_6 = state_out_14_3_6;
  assign port_state_out_14_3_7 = state_out_14_3_7;
  assign port_state_out_15_0_0 = state_out_15_0_0;
  assign port_state_out_15_0_1 = state_out_15_0_1;
  assign port_state_out_15_0_2 = state_out_15_0_2;
  assign port_state_out_15_0_3 = state_out_15_0_3;
  assign port_state_out_15_0_4 = state_out_15_0_4;
  assign port_state_out_15_0_5 = state_out_15_0_5;
  assign port_state_out_15_0_6 = state_out_15_0_6;
  assign port_state_out_15_0_7 = state_out_15_0_7;
  assign port_state_out_15_1_0 = state_out_15_1_0;
  assign port_state_out_15_1_1 = state_out_15_1_1;
  assign port_state_out_15_1_2 = state_out_15_1_2;
  assign port_state_out_15_1_3 = state_out_15_1_3;
  assign port_state_out_15_1_4 = state_out_15_1_4;
  assign port_state_out_15_1_5 = state_out_15_1_5;
  assign port_state_out_15_1_6 = state_out_15_1_6;
  assign port_state_out_15_1_7 = state_out_15_1_7;
  assign port_state_out_15_2_0 = state_out_15_2_0;
  assign port_state_out_15_2_1 = state_out_15_2_1;
  assign port_state_out_15_2_2 = state_out_15_2_2;
  assign port_state_out_15_2_3 = state_out_15_2_3;
  assign port_state_out_15_2_4 = state_out_15_2_4;
  assign port_state_out_15_2_5 = state_out_15_2_5;
  assign port_state_out_15_2_6 = state_out_15_2_6;
  assign port_state_out_15_2_7 = state_out_15_2_7;
  assign port_state_out_15_3_0 = state_out_15_3_0;
  assign port_state_out_15_3_1 = state_out_15_3_1;
  assign port_state_out_15_3_2 = state_out_15_3_2;
  assign port_state_out_15_3_3 = state_out_15_3_3;
  assign port_state_out_15_3_4 = state_out_15_3_4;
  assign port_state_out_15_3_5 = state_out_15_3_5;
  assign port_state_out_15_3_6 = state_out_15_3_6;
  assign port_state_out_15_3_7 = state_out_15_3_7;

endmodule

module AES_ShiftRows (
  input      [0:0]    port_state_in_0_0_0,
  input      [0:0]    port_state_in_0_0_1,
  input      [0:0]    port_state_in_0_0_2,
  input      [0:0]    port_state_in_0_0_3,
  input      [0:0]    port_state_in_0_0_4,
  input      [0:0]    port_state_in_0_0_5,
  input      [0:0]    port_state_in_0_0_6,
  input      [0:0]    port_state_in_0_0_7,
  input      [0:0]    port_state_in_0_1_0,
  input      [0:0]    port_state_in_0_1_1,
  input      [0:0]    port_state_in_0_1_2,
  input      [0:0]    port_state_in_0_1_3,
  input      [0:0]    port_state_in_0_1_4,
  input      [0:0]    port_state_in_0_1_5,
  input      [0:0]    port_state_in_0_1_6,
  input      [0:0]    port_state_in_0_1_7,
  input      [0:0]    port_state_in_0_2_0,
  input      [0:0]    port_state_in_0_2_1,
  input      [0:0]    port_state_in_0_2_2,
  input      [0:0]    port_state_in_0_2_3,
  input      [0:0]    port_state_in_0_2_4,
  input      [0:0]    port_state_in_0_2_5,
  input      [0:0]    port_state_in_0_2_6,
  input      [0:0]    port_state_in_0_2_7,
  input      [0:0]    port_state_in_0_3_0,
  input      [0:0]    port_state_in_0_3_1,
  input      [0:0]    port_state_in_0_3_2,
  input      [0:0]    port_state_in_0_3_3,
  input      [0:0]    port_state_in_0_3_4,
  input      [0:0]    port_state_in_0_3_5,
  input      [0:0]    port_state_in_0_3_6,
  input      [0:0]    port_state_in_0_3_7,
  input      [0:0]    port_state_in_1_0_0,
  input      [0:0]    port_state_in_1_0_1,
  input      [0:0]    port_state_in_1_0_2,
  input      [0:0]    port_state_in_1_0_3,
  input      [0:0]    port_state_in_1_0_4,
  input      [0:0]    port_state_in_1_0_5,
  input      [0:0]    port_state_in_1_0_6,
  input      [0:0]    port_state_in_1_0_7,
  input      [0:0]    port_state_in_1_1_0,
  input      [0:0]    port_state_in_1_1_1,
  input      [0:0]    port_state_in_1_1_2,
  input      [0:0]    port_state_in_1_1_3,
  input      [0:0]    port_state_in_1_1_4,
  input      [0:0]    port_state_in_1_1_5,
  input      [0:0]    port_state_in_1_1_6,
  input      [0:0]    port_state_in_1_1_7,
  input      [0:0]    port_state_in_1_2_0,
  input      [0:0]    port_state_in_1_2_1,
  input      [0:0]    port_state_in_1_2_2,
  input      [0:0]    port_state_in_1_2_3,
  input      [0:0]    port_state_in_1_2_4,
  input      [0:0]    port_state_in_1_2_5,
  input      [0:0]    port_state_in_1_2_6,
  input      [0:0]    port_state_in_1_2_7,
  input      [0:0]    port_state_in_1_3_0,
  input      [0:0]    port_state_in_1_3_1,
  input      [0:0]    port_state_in_1_3_2,
  input      [0:0]    port_state_in_1_3_3,
  input      [0:0]    port_state_in_1_3_4,
  input      [0:0]    port_state_in_1_3_5,
  input      [0:0]    port_state_in_1_3_6,
  input      [0:0]    port_state_in_1_3_7,
  input      [0:0]    port_state_in_2_0_0,
  input      [0:0]    port_state_in_2_0_1,
  input      [0:0]    port_state_in_2_0_2,
  input      [0:0]    port_state_in_2_0_3,
  input      [0:0]    port_state_in_2_0_4,
  input      [0:0]    port_state_in_2_0_5,
  input      [0:0]    port_state_in_2_0_6,
  input      [0:0]    port_state_in_2_0_7,
  input      [0:0]    port_state_in_2_1_0,
  input      [0:0]    port_state_in_2_1_1,
  input      [0:0]    port_state_in_2_1_2,
  input      [0:0]    port_state_in_2_1_3,
  input      [0:0]    port_state_in_2_1_4,
  input      [0:0]    port_state_in_2_1_5,
  input      [0:0]    port_state_in_2_1_6,
  input      [0:0]    port_state_in_2_1_7,
  input      [0:0]    port_state_in_2_2_0,
  input      [0:0]    port_state_in_2_2_1,
  input      [0:0]    port_state_in_2_2_2,
  input      [0:0]    port_state_in_2_2_3,
  input      [0:0]    port_state_in_2_2_4,
  input      [0:0]    port_state_in_2_2_5,
  input      [0:0]    port_state_in_2_2_6,
  input      [0:0]    port_state_in_2_2_7,
  input      [0:0]    port_state_in_2_3_0,
  input      [0:0]    port_state_in_2_3_1,
  input      [0:0]    port_state_in_2_3_2,
  input      [0:0]    port_state_in_2_3_3,
  input      [0:0]    port_state_in_2_3_4,
  input      [0:0]    port_state_in_2_3_5,
  input      [0:0]    port_state_in_2_3_6,
  input      [0:0]    port_state_in_2_3_7,
  input      [0:0]    port_state_in_3_0_0,
  input      [0:0]    port_state_in_3_0_1,
  input      [0:0]    port_state_in_3_0_2,
  input      [0:0]    port_state_in_3_0_3,
  input      [0:0]    port_state_in_3_0_4,
  input      [0:0]    port_state_in_3_0_5,
  input      [0:0]    port_state_in_3_0_6,
  input      [0:0]    port_state_in_3_0_7,
  input      [0:0]    port_state_in_3_1_0,
  input      [0:0]    port_state_in_3_1_1,
  input      [0:0]    port_state_in_3_1_2,
  input      [0:0]    port_state_in_3_1_3,
  input      [0:0]    port_state_in_3_1_4,
  input      [0:0]    port_state_in_3_1_5,
  input      [0:0]    port_state_in_3_1_6,
  input      [0:0]    port_state_in_3_1_7,
  input      [0:0]    port_state_in_3_2_0,
  input      [0:0]    port_state_in_3_2_1,
  input      [0:0]    port_state_in_3_2_2,
  input      [0:0]    port_state_in_3_2_3,
  input      [0:0]    port_state_in_3_2_4,
  input      [0:0]    port_state_in_3_2_5,
  input      [0:0]    port_state_in_3_2_6,
  input      [0:0]    port_state_in_3_2_7,
  input      [0:0]    port_state_in_3_3_0,
  input      [0:0]    port_state_in_3_3_1,
  input      [0:0]    port_state_in_3_3_2,
  input      [0:0]    port_state_in_3_3_3,
  input      [0:0]    port_state_in_3_3_4,
  input      [0:0]    port_state_in_3_3_5,
  input      [0:0]    port_state_in_3_3_6,
  input      [0:0]    port_state_in_3_3_7,
  input      [0:0]    port_state_in_4_0_0,
  input      [0:0]    port_state_in_4_0_1,
  input      [0:0]    port_state_in_4_0_2,
  input      [0:0]    port_state_in_4_0_3,
  input      [0:0]    port_state_in_4_0_4,
  input      [0:0]    port_state_in_4_0_5,
  input      [0:0]    port_state_in_4_0_6,
  input      [0:0]    port_state_in_4_0_7,
  input      [0:0]    port_state_in_4_1_0,
  input      [0:0]    port_state_in_4_1_1,
  input      [0:0]    port_state_in_4_1_2,
  input      [0:0]    port_state_in_4_1_3,
  input      [0:0]    port_state_in_4_1_4,
  input      [0:0]    port_state_in_4_1_5,
  input      [0:0]    port_state_in_4_1_6,
  input      [0:0]    port_state_in_4_1_7,
  input      [0:0]    port_state_in_4_2_0,
  input      [0:0]    port_state_in_4_2_1,
  input      [0:0]    port_state_in_4_2_2,
  input      [0:0]    port_state_in_4_2_3,
  input      [0:0]    port_state_in_4_2_4,
  input      [0:0]    port_state_in_4_2_5,
  input      [0:0]    port_state_in_4_2_6,
  input      [0:0]    port_state_in_4_2_7,
  input      [0:0]    port_state_in_4_3_0,
  input      [0:0]    port_state_in_4_3_1,
  input      [0:0]    port_state_in_4_3_2,
  input      [0:0]    port_state_in_4_3_3,
  input      [0:0]    port_state_in_4_3_4,
  input      [0:0]    port_state_in_4_3_5,
  input      [0:0]    port_state_in_4_3_6,
  input      [0:0]    port_state_in_4_3_7,
  input      [0:0]    port_state_in_5_0_0,
  input      [0:0]    port_state_in_5_0_1,
  input      [0:0]    port_state_in_5_0_2,
  input      [0:0]    port_state_in_5_0_3,
  input      [0:0]    port_state_in_5_0_4,
  input      [0:0]    port_state_in_5_0_5,
  input      [0:0]    port_state_in_5_0_6,
  input      [0:0]    port_state_in_5_0_7,
  input      [0:0]    port_state_in_5_1_0,
  input      [0:0]    port_state_in_5_1_1,
  input      [0:0]    port_state_in_5_1_2,
  input      [0:0]    port_state_in_5_1_3,
  input      [0:0]    port_state_in_5_1_4,
  input      [0:0]    port_state_in_5_1_5,
  input      [0:0]    port_state_in_5_1_6,
  input      [0:0]    port_state_in_5_1_7,
  input      [0:0]    port_state_in_5_2_0,
  input      [0:0]    port_state_in_5_2_1,
  input      [0:0]    port_state_in_5_2_2,
  input      [0:0]    port_state_in_5_2_3,
  input      [0:0]    port_state_in_5_2_4,
  input      [0:0]    port_state_in_5_2_5,
  input      [0:0]    port_state_in_5_2_6,
  input      [0:0]    port_state_in_5_2_7,
  input      [0:0]    port_state_in_5_3_0,
  input      [0:0]    port_state_in_5_3_1,
  input      [0:0]    port_state_in_5_3_2,
  input      [0:0]    port_state_in_5_3_3,
  input      [0:0]    port_state_in_5_3_4,
  input      [0:0]    port_state_in_5_3_5,
  input      [0:0]    port_state_in_5_3_6,
  input      [0:0]    port_state_in_5_3_7,
  input      [0:0]    port_state_in_6_0_0,
  input      [0:0]    port_state_in_6_0_1,
  input      [0:0]    port_state_in_6_0_2,
  input      [0:0]    port_state_in_6_0_3,
  input      [0:0]    port_state_in_6_0_4,
  input      [0:0]    port_state_in_6_0_5,
  input      [0:0]    port_state_in_6_0_6,
  input      [0:0]    port_state_in_6_0_7,
  input      [0:0]    port_state_in_6_1_0,
  input      [0:0]    port_state_in_6_1_1,
  input      [0:0]    port_state_in_6_1_2,
  input      [0:0]    port_state_in_6_1_3,
  input      [0:0]    port_state_in_6_1_4,
  input      [0:0]    port_state_in_6_1_5,
  input      [0:0]    port_state_in_6_1_6,
  input      [0:0]    port_state_in_6_1_7,
  input      [0:0]    port_state_in_6_2_0,
  input      [0:0]    port_state_in_6_2_1,
  input      [0:0]    port_state_in_6_2_2,
  input      [0:0]    port_state_in_6_2_3,
  input      [0:0]    port_state_in_6_2_4,
  input      [0:0]    port_state_in_6_2_5,
  input      [0:0]    port_state_in_6_2_6,
  input      [0:0]    port_state_in_6_2_7,
  input      [0:0]    port_state_in_6_3_0,
  input      [0:0]    port_state_in_6_3_1,
  input      [0:0]    port_state_in_6_3_2,
  input      [0:0]    port_state_in_6_3_3,
  input      [0:0]    port_state_in_6_3_4,
  input      [0:0]    port_state_in_6_3_5,
  input      [0:0]    port_state_in_6_3_6,
  input      [0:0]    port_state_in_6_3_7,
  input      [0:0]    port_state_in_7_0_0,
  input      [0:0]    port_state_in_7_0_1,
  input      [0:0]    port_state_in_7_0_2,
  input      [0:0]    port_state_in_7_0_3,
  input      [0:0]    port_state_in_7_0_4,
  input      [0:0]    port_state_in_7_0_5,
  input      [0:0]    port_state_in_7_0_6,
  input      [0:0]    port_state_in_7_0_7,
  input      [0:0]    port_state_in_7_1_0,
  input      [0:0]    port_state_in_7_1_1,
  input      [0:0]    port_state_in_7_1_2,
  input      [0:0]    port_state_in_7_1_3,
  input      [0:0]    port_state_in_7_1_4,
  input      [0:0]    port_state_in_7_1_5,
  input      [0:0]    port_state_in_7_1_6,
  input      [0:0]    port_state_in_7_1_7,
  input      [0:0]    port_state_in_7_2_0,
  input      [0:0]    port_state_in_7_2_1,
  input      [0:0]    port_state_in_7_2_2,
  input      [0:0]    port_state_in_7_2_3,
  input      [0:0]    port_state_in_7_2_4,
  input      [0:0]    port_state_in_7_2_5,
  input      [0:0]    port_state_in_7_2_6,
  input      [0:0]    port_state_in_7_2_7,
  input      [0:0]    port_state_in_7_3_0,
  input      [0:0]    port_state_in_7_3_1,
  input      [0:0]    port_state_in_7_3_2,
  input      [0:0]    port_state_in_7_3_3,
  input      [0:0]    port_state_in_7_3_4,
  input      [0:0]    port_state_in_7_3_5,
  input      [0:0]    port_state_in_7_3_6,
  input      [0:0]    port_state_in_7_3_7,
  input      [0:0]    port_state_in_8_0_0,
  input      [0:0]    port_state_in_8_0_1,
  input      [0:0]    port_state_in_8_0_2,
  input      [0:0]    port_state_in_8_0_3,
  input      [0:0]    port_state_in_8_0_4,
  input      [0:0]    port_state_in_8_0_5,
  input      [0:0]    port_state_in_8_0_6,
  input      [0:0]    port_state_in_8_0_7,
  input      [0:0]    port_state_in_8_1_0,
  input      [0:0]    port_state_in_8_1_1,
  input      [0:0]    port_state_in_8_1_2,
  input      [0:0]    port_state_in_8_1_3,
  input      [0:0]    port_state_in_8_1_4,
  input      [0:0]    port_state_in_8_1_5,
  input      [0:0]    port_state_in_8_1_6,
  input      [0:0]    port_state_in_8_1_7,
  input      [0:0]    port_state_in_8_2_0,
  input      [0:0]    port_state_in_8_2_1,
  input      [0:0]    port_state_in_8_2_2,
  input      [0:0]    port_state_in_8_2_3,
  input      [0:0]    port_state_in_8_2_4,
  input      [0:0]    port_state_in_8_2_5,
  input      [0:0]    port_state_in_8_2_6,
  input      [0:0]    port_state_in_8_2_7,
  input      [0:0]    port_state_in_8_3_0,
  input      [0:0]    port_state_in_8_3_1,
  input      [0:0]    port_state_in_8_3_2,
  input      [0:0]    port_state_in_8_3_3,
  input      [0:0]    port_state_in_8_3_4,
  input      [0:0]    port_state_in_8_3_5,
  input      [0:0]    port_state_in_8_3_6,
  input      [0:0]    port_state_in_8_3_7,
  input      [0:0]    port_state_in_9_0_0,
  input      [0:0]    port_state_in_9_0_1,
  input      [0:0]    port_state_in_9_0_2,
  input      [0:0]    port_state_in_9_0_3,
  input      [0:0]    port_state_in_9_0_4,
  input      [0:0]    port_state_in_9_0_5,
  input      [0:0]    port_state_in_9_0_6,
  input      [0:0]    port_state_in_9_0_7,
  input      [0:0]    port_state_in_9_1_0,
  input      [0:0]    port_state_in_9_1_1,
  input      [0:0]    port_state_in_9_1_2,
  input      [0:0]    port_state_in_9_1_3,
  input      [0:0]    port_state_in_9_1_4,
  input      [0:0]    port_state_in_9_1_5,
  input      [0:0]    port_state_in_9_1_6,
  input      [0:0]    port_state_in_9_1_7,
  input      [0:0]    port_state_in_9_2_0,
  input      [0:0]    port_state_in_9_2_1,
  input      [0:0]    port_state_in_9_2_2,
  input      [0:0]    port_state_in_9_2_3,
  input      [0:0]    port_state_in_9_2_4,
  input      [0:0]    port_state_in_9_2_5,
  input      [0:0]    port_state_in_9_2_6,
  input      [0:0]    port_state_in_9_2_7,
  input      [0:0]    port_state_in_9_3_0,
  input      [0:0]    port_state_in_9_3_1,
  input      [0:0]    port_state_in_9_3_2,
  input      [0:0]    port_state_in_9_3_3,
  input      [0:0]    port_state_in_9_3_4,
  input      [0:0]    port_state_in_9_3_5,
  input      [0:0]    port_state_in_9_3_6,
  input      [0:0]    port_state_in_9_3_7,
  input      [0:0]    port_state_in_10_0_0,
  input      [0:0]    port_state_in_10_0_1,
  input      [0:0]    port_state_in_10_0_2,
  input      [0:0]    port_state_in_10_0_3,
  input      [0:0]    port_state_in_10_0_4,
  input      [0:0]    port_state_in_10_0_5,
  input      [0:0]    port_state_in_10_0_6,
  input      [0:0]    port_state_in_10_0_7,
  input      [0:0]    port_state_in_10_1_0,
  input      [0:0]    port_state_in_10_1_1,
  input      [0:0]    port_state_in_10_1_2,
  input      [0:0]    port_state_in_10_1_3,
  input      [0:0]    port_state_in_10_1_4,
  input      [0:0]    port_state_in_10_1_5,
  input      [0:0]    port_state_in_10_1_6,
  input      [0:0]    port_state_in_10_1_7,
  input      [0:0]    port_state_in_10_2_0,
  input      [0:0]    port_state_in_10_2_1,
  input      [0:0]    port_state_in_10_2_2,
  input      [0:0]    port_state_in_10_2_3,
  input      [0:0]    port_state_in_10_2_4,
  input      [0:0]    port_state_in_10_2_5,
  input      [0:0]    port_state_in_10_2_6,
  input      [0:0]    port_state_in_10_2_7,
  input      [0:0]    port_state_in_10_3_0,
  input      [0:0]    port_state_in_10_3_1,
  input      [0:0]    port_state_in_10_3_2,
  input      [0:0]    port_state_in_10_3_3,
  input      [0:0]    port_state_in_10_3_4,
  input      [0:0]    port_state_in_10_3_5,
  input      [0:0]    port_state_in_10_3_6,
  input      [0:0]    port_state_in_10_3_7,
  input      [0:0]    port_state_in_11_0_0,
  input      [0:0]    port_state_in_11_0_1,
  input      [0:0]    port_state_in_11_0_2,
  input      [0:0]    port_state_in_11_0_3,
  input      [0:0]    port_state_in_11_0_4,
  input      [0:0]    port_state_in_11_0_5,
  input      [0:0]    port_state_in_11_0_6,
  input      [0:0]    port_state_in_11_0_7,
  input      [0:0]    port_state_in_11_1_0,
  input      [0:0]    port_state_in_11_1_1,
  input      [0:0]    port_state_in_11_1_2,
  input      [0:0]    port_state_in_11_1_3,
  input      [0:0]    port_state_in_11_1_4,
  input      [0:0]    port_state_in_11_1_5,
  input      [0:0]    port_state_in_11_1_6,
  input      [0:0]    port_state_in_11_1_7,
  input      [0:0]    port_state_in_11_2_0,
  input      [0:0]    port_state_in_11_2_1,
  input      [0:0]    port_state_in_11_2_2,
  input      [0:0]    port_state_in_11_2_3,
  input      [0:0]    port_state_in_11_2_4,
  input      [0:0]    port_state_in_11_2_5,
  input      [0:0]    port_state_in_11_2_6,
  input      [0:0]    port_state_in_11_2_7,
  input      [0:0]    port_state_in_11_3_0,
  input      [0:0]    port_state_in_11_3_1,
  input      [0:0]    port_state_in_11_3_2,
  input      [0:0]    port_state_in_11_3_3,
  input      [0:0]    port_state_in_11_3_4,
  input      [0:0]    port_state_in_11_3_5,
  input      [0:0]    port_state_in_11_3_6,
  input      [0:0]    port_state_in_11_3_7,
  input      [0:0]    port_state_in_12_0_0,
  input      [0:0]    port_state_in_12_0_1,
  input      [0:0]    port_state_in_12_0_2,
  input      [0:0]    port_state_in_12_0_3,
  input      [0:0]    port_state_in_12_0_4,
  input      [0:0]    port_state_in_12_0_5,
  input      [0:0]    port_state_in_12_0_6,
  input      [0:0]    port_state_in_12_0_7,
  input      [0:0]    port_state_in_12_1_0,
  input      [0:0]    port_state_in_12_1_1,
  input      [0:0]    port_state_in_12_1_2,
  input      [0:0]    port_state_in_12_1_3,
  input      [0:0]    port_state_in_12_1_4,
  input      [0:0]    port_state_in_12_1_5,
  input      [0:0]    port_state_in_12_1_6,
  input      [0:0]    port_state_in_12_1_7,
  input      [0:0]    port_state_in_12_2_0,
  input      [0:0]    port_state_in_12_2_1,
  input      [0:0]    port_state_in_12_2_2,
  input      [0:0]    port_state_in_12_2_3,
  input      [0:0]    port_state_in_12_2_4,
  input      [0:0]    port_state_in_12_2_5,
  input      [0:0]    port_state_in_12_2_6,
  input      [0:0]    port_state_in_12_2_7,
  input      [0:0]    port_state_in_12_3_0,
  input      [0:0]    port_state_in_12_3_1,
  input      [0:0]    port_state_in_12_3_2,
  input      [0:0]    port_state_in_12_3_3,
  input      [0:0]    port_state_in_12_3_4,
  input      [0:0]    port_state_in_12_3_5,
  input      [0:0]    port_state_in_12_3_6,
  input      [0:0]    port_state_in_12_3_7,
  input      [0:0]    port_state_in_13_0_0,
  input      [0:0]    port_state_in_13_0_1,
  input      [0:0]    port_state_in_13_0_2,
  input      [0:0]    port_state_in_13_0_3,
  input      [0:0]    port_state_in_13_0_4,
  input      [0:0]    port_state_in_13_0_5,
  input      [0:0]    port_state_in_13_0_6,
  input      [0:0]    port_state_in_13_0_7,
  input      [0:0]    port_state_in_13_1_0,
  input      [0:0]    port_state_in_13_1_1,
  input      [0:0]    port_state_in_13_1_2,
  input      [0:0]    port_state_in_13_1_3,
  input      [0:0]    port_state_in_13_1_4,
  input      [0:0]    port_state_in_13_1_5,
  input      [0:0]    port_state_in_13_1_6,
  input      [0:0]    port_state_in_13_1_7,
  input      [0:0]    port_state_in_13_2_0,
  input      [0:0]    port_state_in_13_2_1,
  input      [0:0]    port_state_in_13_2_2,
  input      [0:0]    port_state_in_13_2_3,
  input      [0:0]    port_state_in_13_2_4,
  input      [0:0]    port_state_in_13_2_5,
  input      [0:0]    port_state_in_13_2_6,
  input      [0:0]    port_state_in_13_2_7,
  input      [0:0]    port_state_in_13_3_0,
  input      [0:0]    port_state_in_13_3_1,
  input      [0:0]    port_state_in_13_3_2,
  input      [0:0]    port_state_in_13_3_3,
  input      [0:0]    port_state_in_13_3_4,
  input      [0:0]    port_state_in_13_3_5,
  input      [0:0]    port_state_in_13_3_6,
  input      [0:0]    port_state_in_13_3_7,
  input      [0:0]    port_state_in_14_0_0,
  input      [0:0]    port_state_in_14_0_1,
  input      [0:0]    port_state_in_14_0_2,
  input      [0:0]    port_state_in_14_0_3,
  input      [0:0]    port_state_in_14_0_4,
  input      [0:0]    port_state_in_14_0_5,
  input      [0:0]    port_state_in_14_0_6,
  input      [0:0]    port_state_in_14_0_7,
  input      [0:0]    port_state_in_14_1_0,
  input      [0:0]    port_state_in_14_1_1,
  input      [0:0]    port_state_in_14_1_2,
  input      [0:0]    port_state_in_14_1_3,
  input      [0:0]    port_state_in_14_1_4,
  input      [0:0]    port_state_in_14_1_5,
  input      [0:0]    port_state_in_14_1_6,
  input      [0:0]    port_state_in_14_1_7,
  input      [0:0]    port_state_in_14_2_0,
  input      [0:0]    port_state_in_14_2_1,
  input      [0:0]    port_state_in_14_2_2,
  input      [0:0]    port_state_in_14_2_3,
  input      [0:0]    port_state_in_14_2_4,
  input      [0:0]    port_state_in_14_2_5,
  input      [0:0]    port_state_in_14_2_6,
  input      [0:0]    port_state_in_14_2_7,
  input      [0:0]    port_state_in_14_3_0,
  input      [0:0]    port_state_in_14_3_1,
  input      [0:0]    port_state_in_14_3_2,
  input      [0:0]    port_state_in_14_3_3,
  input      [0:0]    port_state_in_14_3_4,
  input      [0:0]    port_state_in_14_3_5,
  input      [0:0]    port_state_in_14_3_6,
  input      [0:0]    port_state_in_14_3_7,
  input      [0:0]    port_state_in_15_0_0,
  input      [0:0]    port_state_in_15_0_1,
  input      [0:0]    port_state_in_15_0_2,
  input      [0:0]    port_state_in_15_0_3,
  input      [0:0]    port_state_in_15_0_4,
  input      [0:0]    port_state_in_15_0_5,
  input      [0:0]    port_state_in_15_0_6,
  input      [0:0]    port_state_in_15_0_7,
  input      [0:0]    port_state_in_15_1_0,
  input      [0:0]    port_state_in_15_1_1,
  input      [0:0]    port_state_in_15_1_2,
  input      [0:0]    port_state_in_15_1_3,
  input      [0:0]    port_state_in_15_1_4,
  input      [0:0]    port_state_in_15_1_5,
  input      [0:0]    port_state_in_15_1_6,
  input      [0:0]    port_state_in_15_1_7,
  input      [0:0]    port_state_in_15_2_0,
  input      [0:0]    port_state_in_15_2_1,
  input      [0:0]    port_state_in_15_2_2,
  input      [0:0]    port_state_in_15_2_3,
  input      [0:0]    port_state_in_15_2_4,
  input      [0:0]    port_state_in_15_2_5,
  input      [0:0]    port_state_in_15_2_6,
  input      [0:0]    port_state_in_15_2_7,
  input      [0:0]    port_state_in_15_3_0,
  input      [0:0]    port_state_in_15_3_1,
  input      [0:0]    port_state_in_15_3_2,
  input      [0:0]    port_state_in_15_3_3,
  input      [0:0]    port_state_in_15_3_4,
  input      [0:0]    port_state_in_15_3_5,
  input      [0:0]    port_state_in_15_3_6,
  input      [0:0]    port_state_in_15_3_7,
  output     [0:0]    port_state_out_0_0_0,
  output     [0:0]    port_state_out_0_0_1,
  output     [0:0]    port_state_out_0_0_2,
  output     [0:0]    port_state_out_0_0_3,
  output     [0:0]    port_state_out_0_0_4,
  output     [0:0]    port_state_out_0_0_5,
  output     [0:0]    port_state_out_0_0_6,
  output     [0:0]    port_state_out_0_0_7,
  output     [0:0]    port_state_out_0_1_0,
  output     [0:0]    port_state_out_0_1_1,
  output     [0:0]    port_state_out_0_1_2,
  output     [0:0]    port_state_out_0_1_3,
  output     [0:0]    port_state_out_0_1_4,
  output     [0:0]    port_state_out_0_1_5,
  output     [0:0]    port_state_out_0_1_6,
  output     [0:0]    port_state_out_0_1_7,
  output     [0:0]    port_state_out_0_2_0,
  output     [0:0]    port_state_out_0_2_1,
  output     [0:0]    port_state_out_0_2_2,
  output     [0:0]    port_state_out_0_2_3,
  output     [0:0]    port_state_out_0_2_4,
  output     [0:0]    port_state_out_0_2_5,
  output     [0:0]    port_state_out_0_2_6,
  output     [0:0]    port_state_out_0_2_7,
  output     [0:0]    port_state_out_0_3_0,
  output     [0:0]    port_state_out_0_3_1,
  output     [0:0]    port_state_out_0_3_2,
  output     [0:0]    port_state_out_0_3_3,
  output     [0:0]    port_state_out_0_3_4,
  output     [0:0]    port_state_out_0_3_5,
  output     [0:0]    port_state_out_0_3_6,
  output     [0:0]    port_state_out_0_3_7,
  output     [0:0]    port_state_out_1_0_0,
  output     [0:0]    port_state_out_1_0_1,
  output     [0:0]    port_state_out_1_0_2,
  output     [0:0]    port_state_out_1_0_3,
  output     [0:0]    port_state_out_1_0_4,
  output     [0:0]    port_state_out_1_0_5,
  output     [0:0]    port_state_out_1_0_6,
  output     [0:0]    port_state_out_1_0_7,
  output     [0:0]    port_state_out_1_1_0,
  output     [0:0]    port_state_out_1_1_1,
  output     [0:0]    port_state_out_1_1_2,
  output     [0:0]    port_state_out_1_1_3,
  output     [0:0]    port_state_out_1_1_4,
  output     [0:0]    port_state_out_1_1_5,
  output     [0:0]    port_state_out_1_1_6,
  output     [0:0]    port_state_out_1_1_7,
  output     [0:0]    port_state_out_1_2_0,
  output     [0:0]    port_state_out_1_2_1,
  output     [0:0]    port_state_out_1_2_2,
  output     [0:0]    port_state_out_1_2_3,
  output     [0:0]    port_state_out_1_2_4,
  output     [0:0]    port_state_out_1_2_5,
  output     [0:0]    port_state_out_1_2_6,
  output     [0:0]    port_state_out_1_2_7,
  output     [0:0]    port_state_out_1_3_0,
  output     [0:0]    port_state_out_1_3_1,
  output     [0:0]    port_state_out_1_3_2,
  output     [0:0]    port_state_out_1_3_3,
  output     [0:0]    port_state_out_1_3_4,
  output     [0:0]    port_state_out_1_3_5,
  output     [0:0]    port_state_out_1_3_6,
  output     [0:0]    port_state_out_1_3_7,
  output     [0:0]    port_state_out_2_0_0,
  output     [0:0]    port_state_out_2_0_1,
  output     [0:0]    port_state_out_2_0_2,
  output     [0:0]    port_state_out_2_0_3,
  output     [0:0]    port_state_out_2_0_4,
  output     [0:0]    port_state_out_2_0_5,
  output     [0:0]    port_state_out_2_0_6,
  output     [0:0]    port_state_out_2_0_7,
  output     [0:0]    port_state_out_2_1_0,
  output     [0:0]    port_state_out_2_1_1,
  output     [0:0]    port_state_out_2_1_2,
  output     [0:0]    port_state_out_2_1_3,
  output     [0:0]    port_state_out_2_1_4,
  output     [0:0]    port_state_out_2_1_5,
  output     [0:0]    port_state_out_2_1_6,
  output     [0:0]    port_state_out_2_1_7,
  output     [0:0]    port_state_out_2_2_0,
  output     [0:0]    port_state_out_2_2_1,
  output     [0:0]    port_state_out_2_2_2,
  output     [0:0]    port_state_out_2_2_3,
  output     [0:0]    port_state_out_2_2_4,
  output     [0:0]    port_state_out_2_2_5,
  output     [0:0]    port_state_out_2_2_6,
  output     [0:0]    port_state_out_2_2_7,
  output     [0:0]    port_state_out_2_3_0,
  output     [0:0]    port_state_out_2_3_1,
  output     [0:0]    port_state_out_2_3_2,
  output     [0:0]    port_state_out_2_3_3,
  output     [0:0]    port_state_out_2_3_4,
  output     [0:0]    port_state_out_2_3_5,
  output     [0:0]    port_state_out_2_3_6,
  output     [0:0]    port_state_out_2_3_7,
  output     [0:0]    port_state_out_3_0_0,
  output     [0:0]    port_state_out_3_0_1,
  output     [0:0]    port_state_out_3_0_2,
  output     [0:0]    port_state_out_3_0_3,
  output     [0:0]    port_state_out_3_0_4,
  output     [0:0]    port_state_out_3_0_5,
  output     [0:0]    port_state_out_3_0_6,
  output     [0:0]    port_state_out_3_0_7,
  output     [0:0]    port_state_out_3_1_0,
  output     [0:0]    port_state_out_3_1_1,
  output     [0:0]    port_state_out_3_1_2,
  output     [0:0]    port_state_out_3_1_3,
  output     [0:0]    port_state_out_3_1_4,
  output     [0:0]    port_state_out_3_1_5,
  output     [0:0]    port_state_out_3_1_6,
  output     [0:0]    port_state_out_3_1_7,
  output     [0:0]    port_state_out_3_2_0,
  output     [0:0]    port_state_out_3_2_1,
  output     [0:0]    port_state_out_3_2_2,
  output     [0:0]    port_state_out_3_2_3,
  output     [0:0]    port_state_out_3_2_4,
  output     [0:0]    port_state_out_3_2_5,
  output     [0:0]    port_state_out_3_2_6,
  output     [0:0]    port_state_out_3_2_7,
  output     [0:0]    port_state_out_3_3_0,
  output     [0:0]    port_state_out_3_3_1,
  output     [0:0]    port_state_out_3_3_2,
  output     [0:0]    port_state_out_3_3_3,
  output     [0:0]    port_state_out_3_3_4,
  output     [0:0]    port_state_out_3_3_5,
  output     [0:0]    port_state_out_3_3_6,
  output     [0:0]    port_state_out_3_3_7,
  output     [0:0]    port_state_out_4_0_0,
  output     [0:0]    port_state_out_4_0_1,
  output     [0:0]    port_state_out_4_0_2,
  output     [0:0]    port_state_out_4_0_3,
  output     [0:0]    port_state_out_4_0_4,
  output     [0:0]    port_state_out_4_0_5,
  output     [0:0]    port_state_out_4_0_6,
  output     [0:0]    port_state_out_4_0_7,
  output     [0:0]    port_state_out_4_1_0,
  output     [0:0]    port_state_out_4_1_1,
  output     [0:0]    port_state_out_4_1_2,
  output     [0:0]    port_state_out_4_1_3,
  output     [0:0]    port_state_out_4_1_4,
  output     [0:0]    port_state_out_4_1_5,
  output     [0:0]    port_state_out_4_1_6,
  output     [0:0]    port_state_out_4_1_7,
  output     [0:0]    port_state_out_4_2_0,
  output     [0:0]    port_state_out_4_2_1,
  output     [0:0]    port_state_out_4_2_2,
  output     [0:0]    port_state_out_4_2_3,
  output     [0:0]    port_state_out_4_2_4,
  output     [0:0]    port_state_out_4_2_5,
  output     [0:0]    port_state_out_4_2_6,
  output     [0:0]    port_state_out_4_2_7,
  output     [0:0]    port_state_out_4_3_0,
  output     [0:0]    port_state_out_4_3_1,
  output     [0:0]    port_state_out_4_3_2,
  output     [0:0]    port_state_out_4_3_3,
  output     [0:0]    port_state_out_4_3_4,
  output     [0:0]    port_state_out_4_3_5,
  output     [0:0]    port_state_out_4_3_6,
  output     [0:0]    port_state_out_4_3_7,
  output     [0:0]    port_state_out_5_0_0,
  output     [0:0]    port_state_out_5_0_1,
  output     [0:0]    port_state_out_5_0_2,
  output     [0:0]    port_state_out_5_0_3,
  output     [0:0]    port_state_out_5_0_4,
  output     [0:0]    port_state_out_5_0_5,
  output     [0:0]    port_state_out_5_0_6,
  output     [0:0]    port_state_out_5_0_7,
  output     [0:0]    port_state_out_5_1_0,
  output     [0:0]    port_state_out_5_1_1,
  output     [0:0]    port_state_out_5_1_2,
  output     [0:0]    port_state_out_5_1_3,
  output     [0:0]    port_state_out_5_1_4,
  output     [0:0]    port_state_out_5_1_5,
  output     [0:0]    port_state_out_5_1_6,
  output     [0:0]    port_state_out_5_1_7,
  output     [0:0]    port_state_out_5_2_0,
  output     [0:0]    port_state_out_5_2_1,
  output     [0:0]    port_state_out_5_2_2,
  output     [0:0]    port_state_out_5_2_3,
  output     [0:0]    port_state_out_5_2_4,
  output     [0:0]    port_state_out_5_2_5,
  output     [0:0]    port_state_out_5_2_6,
  output     [0:0]    port_state_out_5_2_7,
  output     [0:0]    port_state_out_5_3_0,
  output     [0:0]    port_state_out_5_3_1,
  output     [0:0]    port_state_out_5_3_2,
  output     [0:0]    port_state_out_5_3_3,
  output     [0:0]    port_state_out_5_3_4,
  output     [0:0]    port_state_out_5_3_5,
  output     [0:0]    port_state_out_5_3_6,
  output     [0:0]    port_state_out_5_3_7,
  output     [0:0]    port_state_out_6_0_0,
  output     [0:0]    port_state_out_6_0_1,
  output     [0:0]    port_state_out_6_0_2,
  output     [0:0]    port_state_out_6_0_3,
  output     [0:0]    port_state_out_6_0_4,
  output     [0:0]    port_state_out_6_0_5,
  output     [0:0]    port_state_out_6_0_6,
  output     [0:0]    port_state_out_6_0_7,
  output     [0:0]    port_state_out_6_1_0,
  output     [0:0]    port_state_out_6_1_1,
  output     [0:0]    port_state_out_6_1_2,
  output     [0:0]    port_state_out_6_1_3,
  output     [0:0]    port_state_out_6_1_4,
  output     [0:0]    port_state_out_6_1_5,
  output     [0:0]    port_state_out_6_1_6,
  output     [0:0]    port_state_out_6_1_7,
  output     [0:0]    port_state_out_6_2_0,
  output     [0:0]    port_state_out_6_2_1,
  output     [0:0]    port_state_out_6_2_2,
  output     [0:0]    port_state_out_6_2_3,
  output     [0:0]    port_state_out_6_2_4,
  output     [0:0]    port_state_out_6_2_5,
  output     [0:0]    port_state_out_6_2_6,
  output     [0:0]    port_state_out_6_2_7,
  output     [0:0]    port_state_out_6_3_0,
  output     [0:0]    port_state_out_6_3_1,
  output     [0:0]    port_state_out_6_3_2,
  output     [0:0]    port_state_out_6_3_3,
  output     [0:0]    port_state_out_6_3_4,
  output     [0:0]    port_state_out_6_3_5,
  output     [0:0]    port_state_out_6_3_6,
  output     [0:0]    port_state_out_6_3_7,
  output     [0:0]    port_state_out_7_0_0,
  output     [0:0]    port_state_out_7_0_1,
  output     [0:0]    port_state_out_7_0_2,
  output     [0:0]    port_state_out_7_0_3,
  output     [0:0]    port_state_out_7_0_4,
  output     [0:0]    port_state_out_7_0_5,
  output     [0:0]    port_state_out_7_0_6,
  output     [0:0]    port_state_out_7_0_7,
  output     [0:0]    port_state_out_7_1_0,
  output     [0:0]    port_state_out_7_1_1,
  output     [0:0]    port_state_out_7_1_2,
  output     [0:0]    port_state_out_7_1_3,
  output     [0:0]    port_state_out_7_1_4,
  output     [0:0]    port_state_out_7_1_5,
  output     [0:0]    port_state_out_7_1_6,
  output     [0:0]    port_state_out_7_1_7,
  output     [0:0]    port_state_out_7_2_0,
  output     [0:0]    port_state_out_7_2_1,
  output     [0:0]    port_state_out_7_2_2,
  output     [0:0]    port_state_out_7_2_3,
  output     [0:0]    port_state_out_7_2_4,
  output     [0:0]    port_state_out_7_2_5,
  output     [0:0]    port_state_out_7_2_6,
  output     [0:0]    port_state_out_7_2_7,
  output     [0:0]    port_state_out_7_3_0,
  output     [0:0]    port_state_out_7_3_1,
  output     [0:0]    port_state_out_7_3_2,
  output     [0:0]    port_state_out_7_3_3,
  output     [0:0]    port_state_out_7_3_4,
  output     [0:0]    port_state_out_7_3_5,
  output     [0:0]    port_state_out_7_3_6,
  output     [0:0]    port_state_out_7_3_7,
  output     [0:0]    port_state_out_8_0_0,
  output     [0:0]    port_state_out_8_0_1,
  output     [0:0]    port_state_out_8_0_2,
  output     [0:0]    port_state_out_8_0_3,
  output     [0:0]    port_state_out_8_0_4,
  output     [0:0]    port_state_out_8_0_5,
  output     [0:0]    port_state_out_8_0_6,
  output     [0:0]    port_state_out_8_0_7,
  output     [0:0]    port_state_out_8_1_0,
  output     [0:0]    port_state_out_8_1_1,
  output     [0:0]    port_state_out_8_1_2,
  output     [0:0]    port_state_out_8_1_3,
  output     [0:0]    port_state_out_8_1_4,
  output     [0:0]    port_state_out_8_1_5,
  output     [0:0]    port_state_out_8_1_6,
  output     [0:0]    port_state_out_8_1_7,
  output     [0:0]    port_state_out_8_2_0,
  output     [0:0]    port_state_out_8_2_1,
  output     [0:0]    port_state_out_8_2_2,
  output     [0:0]    port_state_out_8_2_3,
  output     [0:0]    port_state_out_8_2_4,
  output     [0:0]    port_state_out_8_2_5,
  output     [0:0]    port_state_out_8_2_6,
  output     [0:0]    port_state_out_8_2_7,
  output     [0:0]    port_state_out_8_3_0,
  output     [0:0]    port_state_out_8_3_1,
  output     [0:0]    port_state_out_8_3_2,
  output     [0:0]    port_state_out_8_3_3,
  output     [0:0]    port_state_out_8_3_4,
  output     [0:0]    port_state_out_8_3_5,
  output     [0:0]    port_state_out_8_3_6,
  output     [0:0]    port_state_out_8_3_7,
  output     [0:0]    port_state_out_9_0_0,
  output     [0:0]    port_state_out_9_0_1,
  output     [0:0]    port_state_out_9_0_2,
  output     [0:0]    port_state_out_9_0_3,
  output     [0:0]    port_state_out_9_0_4,
  output     [0:0]    port_state_out_9_0_5,
  output     [0:0]    port_state_out_9_0_6,
  output     [0:0]    port_state_out_9_0_7,
  output     [0:0]    port_state_out_9_1_0,
  output     [0:0]    port_state_out_9_1_1,
  output     [0:0]    port_state_out_9_1_2,
  output     [0:0]    port_state_out_9_1_3,
  output     [0:0]    port_state_out_9_1_4,
  output     [0:0]    port_state_out_9_1_5,
  output     [0:0]    port_state_out_9_1_6,
  output     [0:0]    port_state_out_9_1_7,
  output     [0:0]    port_state_out_9_2_0,
  output     [0:0]    port_state_out_9_2_1,
  output     [0:0]    port_state_out_9_2_2,
  output     [0:0]    port_state_out_9_2_3,
  output     [0:0]    port_state_out_9_2_4,
  output     [0:0]    port_state_out_9_2_5,
  output     [0:0]    port_state_out_9_2_6,
  output     [0:0]    port_state_out_9_2_7,
  output     [0:0]    port_state_out_9_3_0,
  output     [0:0]    port_state_out_9_3_1,
  output     [0:0]    port_state_out_9_3_2,
  output     [0:0]    port_state_out_9_3_3,
  output     [0:0]    port_state_out_9_3_4,
  output     [0:0]    port_state_out_9_3_5,
  output     [0:0]    port_state_out_9_3_6,
  output     [0:0]    port_state_out_9_3_7,
  output     [0:0]    port_state_out_10_0_0,
  output     [0:0]    port_state_out_10_0_1,
  output     [0:0]    port_state_out_10_0_2,
  output     [0:0]    port_state_out_10_0_3,
  output     [0:0]    port_state_out_10_0_4,
  output     [0:0]    port_state_out_10_0_5,
  output     [0:0]    port_state_out_10_0_6,
  output     [0:0]    port_state_out_10_0_7,
  output     [0:0]    port_state_out_10_1_0,
  output     [0:0]    port_state_out_10_1_1,
  output     [0:0]    port_state_out_10_1_2,
  output     [0:0]    port_state_out_10_1_3,
  output     [0:0]    port_state_out_10_1_4,
  output     [0:0]    port_state_out_10_1_5,
  output     [0:0]    port_state_out_10_1_6,
  output     [0:0]    port_state_out_10_1_7,
  output     [0:0]    port_state_out_10_2_0,
  output     [0:0]    port_state_out_10_2_1,
  output     [0:0]    port_state_out_10_2_2,
  output     [0:0]    port_state_out_10_2_3,
  output     [0:0]    port_state_out_10_2_4,
  output     [0:0]    port_state_out_10_2_5,
  output     [0:0]    port_state_out_10_2_6,
  output     [0:0]    port_state_out_10_2_7,
  output     [0:0]    port_state_out_10_3_0,
  output     [0:0]    port_state_out_10_3_1,
  output     [0:0]    port_state_out_10_3_2,
  output     [0:0]    port_state_out_10_3_3,
  output     [0:0]    port_state_out_10_3_4,
  output     [0:0]    port_state_out_10_3_5,
  output     [0:0]    port_state_out_10_3_6,
  output     [0:0]    port_state_out_10_3_7,
  output     [0:0]    port_state_out_11_0_0,
  output     [0:0]    port_state_out_11_0_1,
  output     [0:0]    port_state_out_11_0_2,
  output     [0:0]    port_state_out_11_0_3,
  output     [0:0]    port_state_out_11_0_4,
  output     [0:0]    port_state_out_11_0_5,
  output     [0:0]    port_state_out_11_0_6,
  output     [0:0]    port_state_out_11_0_7,
  output     [0:0]    port_state_out_11_1_0,
  output     [0:0]    port_state_out_11_1_1,
  output     [0:0]    port_state_out_11_1_2,
  output     [0:0]    port_state_out_11_1_3,
  output     [0:0]    port_state_out_11_1_4,
  output     [0:0]    port_state_out_11_1_5,
  output     [0:0]    port_state_out_11_1_6,
  output     [0:0]    port_state_out_11_1_7,
  output     [0:0]    port_state_out_11_2_0,
  output     [0:0]    port_state_out_11_2_1,
  output     [0:0]    port_state_out_11_2_2,
  output     [0:0]    port_state_out_11_2_3,
  output     [0:0]    port_state_out_11_2_4,
  output     [0:0]    port_state_out_11_2_5,
  output     [0:0]    port_state_out_11_2_6,
  output     [0:0]    port_state_out_11_2_7,
  output     [0:0]    port_state_out_11_3_0,
  output     [0:0]    port_state_out_11_3_1,
  output     [0:0]    port_state_out_11_3_2,
  output     [0:0]    port_state_out_11_3_3,
  output     [0:0]    port_state_out_11_3_4,
  output     [0:0]    port_state_out_11_3_5,
  output     [0:0]    port_state_out_11_3_6,
  output     [0:0]    port_state_out_11_3_7,
  output     [0:0]    port_state_out_12_0_0,
  output     [0:0]    port_state_out_12_0_1,
  output     [0:0]    port_state_out_12_0_2,
  output     [0:0]    port_state_out_12_0_3,
  output     [0:0]    port_state_out_12_0_4,
  output     [0:0]    port_state_out_12_0_5,
  output     [0:0]    port_state_out_12_0_6,
  output     [0:0]    port_state_out_12_0_7,
  output     [0:0]    port_state_out_12_1_0,
  output     [0:0]    port_state_out_12_1_1,
  output     [0:0]    port_state_out_12_1_2,
  output     [0:0]    port_state_out_12_1_3,
  output     [0:0]    port_state_out_12_1_4,
  output     [0:0]    port_state_out_12_1_5,
  output     [0:0]    port_state_out_12_1_6,
  output     [0:0]    port_state_out_12_1_7,
  output     [0:0]    port_state_out_12_2_0,
  output     [0:0]    port_state_out_12_2_1,
  output     [0:0]    port_state_out_12_2_2,
  output     [0:0]    port_state_out_12_2_3,
  output     [0:0]    port_state_out_12_2_4,
  output     [0:0]    port_state_out_12_2_5,
  output     [0:0]    port_state_out_12_2_6,
  output     [0:0]    port_state_out_12_2_7,
  output     [0:0]    port_state_out_12_3_0,
  output     [0:0]    port_state_out_12_3_1,
  output     [0:0]    port_state_out_12_3_2,
  output     [0:0]    port_state_out_12_3_3,
  output     [0:0]    port_state_out_12_3_4,
  output     [0:0]    port_state_out_12_3_5,
  output     [0:0]    port_state_out_12_3_6,
  output     [0:0]    port_state_out_12_3_7,
  output     [0:0]    port_state_out_13_0_0,
  output     [0:0]    port_state_out_13_0_1,
  output     [0:0]    port_state_out_13_0_2,
  output     [0:0]    port_state_out_13_0_3,
  output     [0:0]    port_state_out_13_0_4,
  output     [0:0]    port_state_out_13_0_5,
  output     [0:0]    port_state_out_13_0_6,
  output     [0:0]    port_state_out_13_0_7,
  output     [0:0]    port_state_out_13_1_0,
  output     [0:0]    port_state_out_13_1_1,
  output     [0:0]    port_state_out_13_1_2,
  output     [0:0]    port_state_out_13_1_3,
  output     [0:0]    port_state_out_13_1_4,
  output     [0:0]    port_state_out_13_1_5,
  output     [0:0]    port_state_out_13_1_6,
  output     [0:0]    port_state_out_13_1_7,
  output     [0:0]    port_state_out_13_2_0,
  output     [0:0]    port_state_out_13_2_1,
  output     [0:0]    port_state_out_13_2_2,
  output     [0:0]    port_state_out_13_2_3,
  output     [0:0]    port_state_out_13_2_4,
  output     [0:0]    port_state_out_13_2_5,
  output     [0:0]    port_state_out_13_2_6,
  output     [0:0]    port_state_out_13_2_7,
  output     [0:0]    port_state_out_13_3_0,
  output     [0:0]    port_state_out_13_3_1,
  output     [0:0]    port_state_out_13_3_2,
  output     [0:0]    port_state_out_13_3_3,
  output     [0:0]    port_state_out_13_3_4,
  output     [0:0]    port_state_out_13_3_5,
  output     [0:0]    port_state_out_13_3_6,
  output     [0:0]    port_state_out_13_3_7,
  output     [0:0]    port_state_out_14_0_0,
  output     [0:0]    port_state_out_14_0_1,
  output     [0:0]    port_state_out_14_0_2,
  output     [0:0]    port_state_out_14_0_3,
  output     [0:0]    port_state_out_14_0_4,
  output     [0:0]    port_state_out_14_0_5,
  output     [0:0]    port_state_out_14_0_6,
  output     [0:0]    port_state_out_14_0_7,
  output     [0:0]    port_state_out_14_1_0,
  output     [0:0]    port_state_out_14_1_1,
  output     [0:0]    port_state_out_14_1_2,
  output     [0:0]    port_state_out_14_1_3,
  output     [0:0]    port_state_out_14_1_4,
  output     [0:0]    port_state_out_14_1_5,
  output     [0:0]    port_state_out_14_1_6,
  output     [0:0]    port_state_out_14_1_7,
  output     [0:0]    port_state_out_14_2_0,
  output     [0:0]    port_state_out_14_2_1,
  output     [0:0]    port_state_out_14_2_2,
  output     [0:0]    port_state_out_14_2_3,
  output     [0:0]    port_state_out_14_2_4,
  output     [0:0]    port_state_out_14_2_5,
  output     [0:0]    port_state_out_14_2_6,
  output     [0:0]    port_state_out_14_2_7,
  output     [0:0]    port_state_out_14_3_0,
  output     [0:0]    port_state_out_14_3_1,
  output     [0:0]    port_state_out_14_3_2,
  output     [0:0]    port_state_out_14_3_3,
  output     [0:0]    port_state_out_14_3_4,
  output     [0:0]    port_state_out_14_3_5,
  output     [0:0]    port_state_out_14_3_6,
  output     [0:0]    port_state_out_14_3_7,
  output     [0:0]    port_state_out_15_0_0,
  output     [0:0]    port_state_out_15_0_1,
  output     [0:0]    port_state_out_15_0_2,
  output     [0:0]    port_state_out_15_0_3,
  output     [0:0]    port_state_out_15_0_4,
  output     [0:0]    port_state_out_15_0_5,
  output     [0:0]    port_state_out_15_0_6,
  output     [0:0]    port_state_out_15_0_7,
  output     [0:0]    port_state_out_15_1_0,
  output     [0:0]    port_state_out_15_1_1,
  output     [0:0]    port_state_out_15_1_2,
  output     [0:0]    port_state_out_15_1_3,
  output     [0:0]    port_state_out_15_1_4,
  output     [0:0]    port_state_out_15_1_5,
  output     [0:0]    port_state_out_15_1_6,
  output     [0:0]    port_state_out_15_1_7,
  output     [0:0]    port_state_out_15_2_0,
  output     [0:0]    port_state_out_15_2_1,
  output     [0:0]    port_state_out_15_2_2,
  output     [0:0]    port_state_out_15_2_3,
  output     [0:0]    port_state_out_15_2_4,
  output     [0:0]    port_state_out_15_2_5,
  output     [0:0]    port_state_out_15_2_6,
  output     [0:0]    port_state_out_15_2_7,
  output     [0:0]    port_state_out_15_3_0,
  output     [0:0]    port_state_out_15_3_1,
  output     [0:0]    port_state_out_15_3_2,
  output     [0:0]    port_state_out_15_3_3,
  output     [0:0]    port_state_out_15_3_4,
  output     [0:0]    port_state_out_15_3_5,
  output     [0:0]    port_state_out_15_3_6,
  output     [0:0]    port_state_out_15_3_7
);


  assign port_state_out_0_0_0 = port_state_in_0_0_0;
  assign port_state_out_0_0_1 = port_state_in_0_0_1;
  assign port_state_out_0_0_2 = port_state_in_0_0_2;
  assign port_state_out_0_0_3 = port_state_in_0_0_3;
  assign port_state_out_0_0_4 = port_state_in_0_0_4;
  assign port_state_out_0_0_5 = port_state_in_0_0_5;
  assign port_state_out_0_0_6 = port_state_in_0_0_6;
  assign port_state_out_0_0_7 = port_state_in_0_0_7;
  assign port_state_out_0_1_0 = port_state_in_0_1_0;
  assign port_state_out_0_1_1 = port_state_in_0_1_1;
  assign port_state_out_0_1_2 = port_state_in_0_1_2;
  assign port_state_out_0_1_3 = port_state_in_0_1_3;
  assign port_state_out_0_1_4 = port_state_in_0_1_4;
  assign port_state_out_0_1_5 = port_state_in_0_1_5;
  assign port_state_out_0_1_6 = port_state_in_0_1_6;
  assign port_state_out_0_1_7 = port_state_in_0_1_7;
  assign port_state_out_0_2_0 = port_state_in_0_2_0;
  assign port_state_out_0_2_1 = port_state_in_0_2_1;
  assign port_state_out_0_2_2 = port_state_in_0_2_2;
  assign port_state_out_0_2_3 = port_state_in_0_2_3;
  assign port_state_out_0_2_4 = port_state_in_0_2_4;
  assign port_state_out_0_2_5 = port_state_in_0_2_5;
  assign port_state_out_0_2_6 = port_state_in_0_2_6;
  assign port_state_out_0_2_7 = port_state_in_0_2_7;
  assign port_state_out_0_3_0 = port_state_in_0_3_0;
  assign port_state_out_0_3_1 = port_state_in_0_3_1;
  assign port_state_out_0_3_2 = port_state_in_0_3_2;
  assign port_state_out_0_3_3 = port_state_in_0_3_3;
  assign port_state_out_0_3_4 = port_state_in_0_3_4;
  assign port_state_out_0_3_5 = port_state_in_0_3_5;
  assign port_state_out_0_3_6 = port_state_in_0_3_6;
  assign port_state_out_0_3_7 = port_state_in_0_3_7;
  assign port_state_out_1_0_0 = port_state_in_5_0_0;
  assign port_state_out_1_0_1 = port_state_in_5_0_1;
  assign port_state_out_1_0_2 = port_state_in_5_0_2;
  assign port_state_out_1_0_3 = port_state_in_5_0_3;
  assign port_state_out_1_0_4 = port_state_in_5_0_4;
  assign port_state_out_1_0_5 = port_state_in_5_0_5;
  assign port_state_out_1_0_6 = port_state_in_5_0_6;
  assign port_state_out_1_0_7 = port_state_in_5_0_7;
  assign port_state_out_1_1_0 = port_state_in_5_1_0;
  assign port_state_out_1_1_1 = port_state_in_5_1_1;
  assign port_state_out_1_1_2 = port_state_in_5_1_2;
  assign port_state_out_1_1_3 = port_state_in_5_1_3;
  assign port_state_out_1_1_4 = port_state_in_5_1_4;
  assign port_state_out_1_1_5 = port_state_in_5_1_5;
  assign port_state_out_1_1_6 = port_state_in_5_1_6;
  assign port_state_out_1_1_7 = port_state_in_5_1_7;
  assign port_state_out_1_2_0 = port_state_in_5_2_0;
  assign port_state_out_1_2_1 = port_state_in_5_2_1;
  assign port_state_out_1_2_2 = port_state_in_5_2_2;
  assign port_state_out_1_2_3 = port_state_in_5_2_3;
  assign port_state_out_1_2_4 = port_state_in_5_2_4;
  assign port_state_out_1_2_5 = port_state_in_5_2_5;
  assign port_state_out_1_2_6 = port_state_in_5_2_6;
  assign port_state_out_1_2_7 = port_state_in_5_2_7;
  assign port_state_out_1_3_0 = port_state_in_5_3_0;
  assign port_state_out_1_3_1 = port_state_in_5_3_1;
  assign port_state_out_1_3_2 = port_state_in_5_3_2;
  assign port_state_out_1_3_3 = port_state_in_5_3_3;
  assign port_state_out_1_3_4 = port_state_in_5_3_4;
  assign port_state_out_1_3_5 = port_state_in_5_3_5;
  assign port_state_out_1_3_6 = port_state_in_5_3_6;
  assign port_state_out_1_3_7 = port_state_in_5_3_7;
  assign port_state_out_2_0_0 = port_state_in_10_0_0;
  assign port_state_out_2_0_1 = port_state_in_10_0_1;
  assign port_state_out_2_0_2 = port_state_in_10_0_2;
  assign port_state_out_2_0_3 = port_state_in_10_0_3;
  assign port_state_out_2_0_4 = port_state_in_10_0_4;
  assign port_state_out_2_0_5 = port_state_in_10_0_5;
  assign port_state_out_2_0_6 = port_state_in_10_0_6;
  assign port_state_out_2_0_7 = port_state_in_10_0_7;
  assign port_state_out_2_1_0 = port_state_in_10_1_0;
  assign port_state_out_2_1_1 = port_state_in_10_1_1;
  assign port_state_out_2_1_2 = port_state_in_10_1_2;
  assign port_state_out_2_1_3 = port_state_in_10_1_3;
  assign port_state_out_2_1_4 = port_state_in_10_1_4;
  assign port_state_out_2_1_5 = port_state_in_10_1_5;
  assign port_state_out_2_1_6 = port_state_in_10_1_6;
  assign port_state_out_2_1_7 = port_state_in_10_1_7;
  assign port_state_out_2_2_0 = port_state_in_10_2_0;
  assign port_state_out_2_2_1 = port_state_in_10_2_1;
  assign port_state_out_2_2_2 = port_state_in_10_2_2;
  assign port_state_out_2_2_3 = port_state_in_10_2_3;
  assign port_state_out_2_2_4 = port_state_in_10_2_4;
  assign port_state_out_2_2_5 = port_state_in_10_2_5;
  assign port_state_out_2_2_6 = port_state_in_10_2_6;
  assign port_state_out_2_2_7 = port_state_in_10_2_7;
  assign port_state_out_2_3_0 = port_state_in_10_3_0;
  assign port_state_out_2_3_1 = port_state_in_10_3_1;
  assign port_state_out_2_3_2 = port_state_in_10_3_2;
  assign port_state_out_2_3_3 = port_state_in_10_3_3;
  assign port_state_out_2_3_4 = port_state_in_10_3_4;
  assign port_state_out_2_3_5 = port_state_in_10_3_5;
  assign port_state_out_2_3_6 = port_state_in_10_3_6;
  assign port_state_out_2_3_7 = port_state_in_10_3_7;
  assign port_state_out_3_0_0 = port_state_in_15_0_0;
  assign port_state_out_3_0_1 = port_state_in_15_0_1;
  assign port_state_out_3_0_2 = port_state_in_15_0_2;
  assign port_state_out_3_0_3 = port_state_in_15_0_3;
  assign port_state_out_3_0_4 = port_state_in_15_0_4;
  assign port_state_out_3_0_5 = port_state_in_15_0_5;
  assign port_state_out_3_0_6 = port_state_in_15_0_6;
  assign port_state_out_3_0_7 = port_state_in_15_0_7;
  assign port_state_out_3_1_0 = port_state_in_15_1_0;
  assign port_state_out_3_1_1 = port_state_in_15_1_1;
  assign port_state_out_3_1_2 = port_state_in_15_1_2;
  assign port_state_out_3_1_3 = port_state_in_15_1_3;
  assign port_state_out_3_1_4 = port_state_in_15_1_4;
  assign port_state_out_3_1_5 = port_state_in_15_1_5;
  assign port_state_out_3_1_6 = port_state_in_15_1_6;
  assign port_state_out_3_1_7 = port_state_in_15_1_7;
  assign port_state_out_3_2_0 = port_state_in_15_2_0;
  assign port_state_out_3_2_1 = port_state_in_15_2_1;
  assign port_state_out_3_2_2 = port_state_in_15_2_2;
  assign port_state_out_3_2_3 = port_state_in_15_2_3;
  assign port_state_out_3_2_4 = port_state_in_15_2_4;
  assign port_state_out_3_2_5 = port_state_in_15_2_5;
  assign port_state_out_3_2_6 = port_state_in_15_2_6;
  assign port_state_out_3_2_7 = port_state_in_15_2_7;
  assign port_state_out_3_3_0 = port_state_in_15_3_0;
  assign port_state_out_3_3_1 = port_state_in_15_3_1;
  assign port_state_out_3_3_2 = port_state_in_15_3_2;
  assign port_state_out_3_3_3 = port_state_in_15_3_3;
  assign port_state_out_3_3_4 = port_state_in_15_3_4;
  assign port_state_out_3_3_5 = port_state_in_15_3_5;
  assign port_state_out_3_3_6 = port_state_in_15_3_6;
  assign port_state_out_3_3_7 = port_state_in_15_3_7;
  assign port_state_out_4_0_0 = port_state_in_4_0_0;
  assign port_state_out_4_0_1 = port_state_in_4_0_1;
  assign port_state_out_4_0_2 = port_state_in_4_0_2;
  assign port_state_out_4_0_3 = port_state_in_4_0_3;
  assign port_state_out_4_0_4 = port_state_in_4_0_4;
  assign port_state_out_4_0_5 = port_state_in_4_0_5;
  assign port_state_out_4_0_6 = port_state_in_4_0_6;
  assign port_state_out_4_0_7 = port_state_in_4_0_7;
  assign port_state_out_4_1_0 = port_state_in_4_1_0;
  assign port_state_out_4_1_1 = port_state_in_4_1_1;
  assign port_state_out_4_1_2 = port_state_in_4_1_2;
  assign port_state_out_4_1_3 = port_state_in_4_1_3;
  assign port_state_out_4_1_4 = port_state_in_4_1_4;
  assign port_state_out_4_1_5 = port_state_in_4_1_5;
  assign port_state_out_4_1_6 = port_state_in_4_1_6;
  assign port_state_out_4_1_7 = port_state_in_4_1_7;
  assign port_state_out_4_2_0 = port_state_in_4_2_0;
  assign port_state_out_4_2_1 = port_state_in_4_2_1;
  assign port_state_out_4_2_2 = port_state_in_4_2_2;
  assign port_state_out_4_2_3 = port_state_in_4_2_3;
  assign port_state_out_4_2_4 = port_state_in_4_2_4;
  assign port_state_out_4_2_5 = port_state_in_4_2_5;
  assign port_state_out_4_2_6 = port_state_in_4_2_6;
  assign port_state_out_4_2_7 = port_state_in_4_2_7;
  assign port_state_out_4_3_0 = port_state_in_4_3_0;
  assign port_state_out_4_3_1 = port_state_in_4_3_1;
  assign port_state_out_4_3_2 = port_state_in_4_3_2;
  assign port_state_out_4_3_3 = port_state_in_4_3_3;
  assign port_state_out_4_3_4 = port_state_in_4_3_4;
  assign port_state_out_4_3_5 = port_state_in_4_3_5;
  assign port_state_out_4_3_6 = port_state_in_4_3_6;
  assign port_state_out_4_3_7 = port_state_in_4_3_7;
  assign port_state_out_5_0_0 = port_state_in_9_0_0;
  assign port_state_out_5_0_1 = port_state_in_9_0_1;
  assign port_state_out_5_0_2 = port_state_in_9_0_2;
  assign port_state_out_5_0_3 = port_state_in_9_0_3;
  assign port_state_out_5_0_4 = port_state_in_9_0_4;
  assign port_state_out_5_0_5 = port_state_in_9_0_5;
  assign port_state_out_5_0_6 = port_state_in_9_0_6;
  assign port_state_out_5_0_7 = port_state_in_9_0_7;
  assign port_state_out_5_1_0 = port_state_in_9_1_0;
  assign port_state_out_5_1_1 = port_state_in_9_1_1;
  assign port_state_out_5_1_2 = port_state_in_9_1_2;
  assign port_state_out_5_1_3 = port_state_in_9_1_3;
  assign port_state_out_5_1_4 = port_state_in_9_1_4;
  assign port_state_out_5_1_5 = port_state_in_9_1_5;
  assign port_state_out_5_1_6 = port_state_in_9_1_6;
  assign port_state_out_5_1_7 = port_state_in_9_1_7;
  assign port_state_out_5_2_0 = port_state_in_9_2_0;
  assign port_state_out_5_2_1 = port_state_in_9_2_1;
  assign port_state_out_5_2_2 = port_state_in_9_2_2;
  assign port_state_out_5_2_3 = port_state_in_9_2_3;
  assign port_state_out_5_2_4 = port_state_in_9_2_4;
  assign port_state_out_5_2_5 = port_state_in_9_2_5;
  assign port_state_out_5_2_6 = port_state_in_9_2_6;
  assign port_state_out_5_2_7 = port_state_in_9_2_7;
  assign port_state_out_5_3_0 = port_state_in_9_3_0;
  assign port_state_out_5_3_1 = port_state_in_9_3_1;
  assign port_state_out_5_3_2 = port_state_in_9_3_2;
  assign port_state_out_5_3_3 = port_state_in_9_3_3;
  assign port_state_out_5_3_4 = port_state_in_9_3_4;
  assign port_state_out_5_3_5 = port_state_in_9_3_5;
  assign port_state_out_5_3_6 = port_state_in_9_3_6;
  assign port_state_out_5_3_7 = port_state_in_9_3_7;
  assign port_state_out_6_0_0 = port_state_in_14_0_0;
  assign port_state_out_6_0_1 = port_state_in_14_0_1;
  assign port_state_out_6_0_2 = port_state_in_14_0_2;
  assign port_state_out_6_0_3 = port_state_in_14_0_3;
  assign port_state_out_6_0_4 = port_state_in_14_0_4;
  assign port_state_out_6_0_5 = port_state_in_14_0_5;
  assign port_state_out_6_0_6 = port_state_in_14_0_6;
  assign port_state_out_6_0_7 = port_state_in_14_0_7;
  assign port_state_out_6_1_0 = port_state_in_14_1_0;
  assign port_state_out_6_1_1 = port_state_in_14_1_1;
  assign port_state_out_6_1_2 = port_state_in_14_1_2;
  assign port_state_out_6_1_3 = port_state_in_14_1_3;
  assign port_state_out_6_1_4 = port_state_in_14_1_4;
  assign port_state_out_6_1_5 = port_state_in_14_1_5;
  assign port_state_out_6_1_6 = port_state_in_14_1_6;
  assign port_state_out_6_1_7 = port_state_in_14_1_7;
  assign port_state_out_6_2_0 = port_state_in_14_2_0;
  assign port_state_out_6_2_1 = port_state_in_14_2_1;
  assign port_state_out_6_2_2 = port_state_in_14_2_2;
  assign port_state_out_6_2_3 = port_state_in_14_2_3;
  assign port_state_out_6_2_4 = port_state_in_14_2_4;
  assign port_state_out_6_2_5 = port_state_in_14_2_5;
  assign port_state_out_6_2_6 = port_state_in_14_2_6;
  assign port_state_out_6_2_7 = port_state_in_14_2_7;
  assign port_state_out_6_3_0 = port_state_in_14_3_0;
  assign port_state_out_6_3_1 = port_state_in_14_3_1;
  assign port_state_out_6_3_2 = port_state_in_14_3_2;
  assign port_state_out_6_3_3 = port_state_in_14_3_3;
  assign port_state_out_6_3_4 = port_state_in_14_3_4;
  assign port_state_out_6_3_5 = port_state_in_14_3_5;
  assign port_state_out_6_3_6 = port_state_in_14_3_6;
  assign port_state_out_6_3_7 = port_state_in_14_3_7;
  assign port_state_out_7_0_0 = port_state_in_3_0_0;
  assign port_state_out_7_0_1 = port_state_in_3_0_1;
  assign port_state_out_7_0_2 = port_state_in_3_0_2;
  assign port_state_out_7_0_3 = port_state_in_3_0_3;
  assign port_state_out_7_0_4 = port_state_in_3_0_4;
  assign port_state_out_7_0_5 = port_state_in_3_0_5;
  assign port_state_out_7_0_6 = port_state_in_3_0_6;
  assign port_state_out_7_0_7 = port_state_in_3_0_7;
  assign port_state_out_7_1_0 = port_state_in_3_1_0;
  assign port_state_out_7_1_1 = port_state_in_3_1_1;
  assign port_state_out_7_1_2 = port_state_in_3_1_2;
  assign port_state_out_7_1_3 = port_state_in_3_1_3;
  assign port_state_out_7_1_4 = port_state_in_3_1_4;
  assign port_state_out_7_1_5 = port_state_in_3_1_5;
  assign port_state_out_7_1_6 = port_state_in_3_1_6;
  assign port_state_out_7_1_7 = port_state_in_3_1_7;
  assign port_state_out_7_2_0 = port_state_in_3_2_0;
  assign port_state_out_7_2_1 = port_state_in_3_2_1;
  assign port_state_out_7_2_2 = port_state_in_3_2_2;
  assign port_state_out_7_2_3 = port_state_in_3_2_3;
  assign port_state_out_7_2_4 = port_state_in_3_2_4;
  assign port_state_out_7_2_5 = port_state_in_3_2_5;
  assign port_state_out_7_2_6 = port_state_in_3_2_6;
  assign port_state_out_7_2_7 = port_state_in_3_2_7;
  assign port_state_out_7_3_0 = port_state_in_3_3_0;
  assign port_state_out_7_3_1 = port_state_in_3_3_1;
  assign port_state_out_7_3_2 = port_state_in_3_3_2;
  assign port_state_out_7_3_3 = port_state_in_3_3_3;
  assign port_state_out_7_3_4 = port_state_in_3_3_4;
  assign port_state_out_7_3_5 = port_state_in_3_3_5;
  assign port_state_out_7_3_6 = port_state_in_3_3_6;
  assign port_state_out_7_3_7 = port_state_in_3_3_7;
  assign port_state_out_8_0_0 = port_state_in_8_0_0;
  assign port_state_out_8_0_1 = port_state_in_8_0_1;
  assign port_state_out_8_0_2 = port_state_in_8_0_2;
  assign port_state_out_8_0_3 = port_state_in_8_0_3;
  assign port_state_out_8_0_4 = port_state_in_8_0_4;
  assign port_state_out_8_0_5 = port_state_in_8_0_5;
  assign port_state_out_8_0_6 = port_state_in_8_0_6;
  assign port_state_out_8_0_7 = port_state_in_8_0_7;
  assign port_state_out_8_1_0 = port_state_in_8_1_0;
  assign port_state_out_8_1_1 = port_state_in_8_1_1;
  assign port_state_out_8_1_2 = port_state_in_8_1_2;
  assign port_state_out_8_1_3 = port_state_in_8_1_3;
  assign port_state_out_8_1_4 = port_state_in_8_1_4;
  assign port_state_out_8_1_5 = port_state_in_8_1_5;
  assign port_state_out_8_1_6 = port_state_in_8_1_6;
  assign port_state_out_8_1_7 = port_state_in_8_1_7;
  assign port_state_out_8_2_0 = port_state_in_8_2_0;
  assign port_state_out_8_2_1 = port_state_in_8_2_1;
  assign port_state_out_8_2_2 = port_state_in_8_2_2;
  assign port_state_out_8_2_3 = port_state_in_8_2_3;
  assign port_state_out_8_2_4 = port_state_in_8_2_4;
  assign port_state_out_8_2_5 = port_state_in_8_2_5;
  assign port_state_out_8_2_6 = port_state_in_8_2_6;
  assign port_state_out_8_2_7 = port_state_in_8_2_7;
  assign port_state_out_8_3_0 = port_state_in_8_3_0;
  assign port_state_out_8_3_1 = port_state_in_8_3_1;
  assign port_state_out_8_3_2 = port_state_in_8_3_2;
  assign port_state_out_8_3_3 = port_state_in_8_3_3;
  assign port_state_out_8_3_4 = port_state_in_8_3_4;
  assign port_state_out_8_3_5 = port_state_in_8_3_5;
  assign port_state_out_8_3_6 = port_state_in_8_3_6;
  assign port_state_out_8_3_7 = port_state_in_8_3_7;
  assign port_state_out_9_0_0 = port_state_in_13_0_0;
  assign port_state_out_9_0_1 = port_state_in_13_0_1;
  assign port_state_out_9_0_2 = port_state_in_13_0_2;
  assign port_state_out_9_0_3 = port_state_in_13_0_3;
  assign port_state_out_9_0_4 = port_state_in_13_0_4;
  assign port_state_out_9_0_5 = port_state_in_13_0_5;
  assign port_state_out_9_0_6 = port_state_in_13_0_6;
  assign port_state_out_9_0_7 = port_state_in_13_0_7;
  assign port_state_out_9_1_0 = port_state_in_13_1_0;
  assign port_state_out_9_1_1 = port_state_in_13_1_1;
  assign port_state_out_9_1_2 = port_state_in_13_1_2;
  assign port_state_out_9_1_3 = port_state_in_13_1_3;
  assign port_state_out_9_1_4 = port_state_in_13_1_4;
  assign port_state_out_9_1_5 = port_state_in_13_1_5;
  assign port_state_out_9_1_6 = port_state_in_13_1_6;
  assign port_state_out_9_1_7 = port_state_in_13_1_7;
  assign port_state_out_9_2_0 = port_state_in_13_2_0;
  assign port_state_out_9_2_1 = port_state_in_13_2_1;
  assign port_state_out_9_2_2 = port_state_in_13_2_2;
  assign port_state_out_9_2_3 = port_state_in_13_2_3;
  assign port_state_out_9_2_4 = port_state_in_13_2_4;
  assign port_state_out_9_2_5 = port_state_in_13_2_5;
  assign port_state_out_9_2_6 = port_state_in_13_2_6;
  assign port_state_out_9_2_7 = port_state_in_13_2_7;
  assign port_state_out_9_3_0 = port_state_in_13_3_0;
  assign port_state_out_9_3_1 = port_state_in_13_3_1;
  assign port_state_out_9_3_2 = port_state_in_13_3_2;
  assign port_state_out_9_3_3 = port_state_in_13_3_3;
  assign port_state_out_9_3_4 = port_state_in_13_3_4;
  assign port_state_out_9_3_5 = port_state_in_13_3_5;
  assign port_state_out_9_3_6 = port_state_in_13_3_6;
  assign port_state_out_9_3_7 = port_state_in_13_3_7;
  assign port_state_out_10_0_0 = port_state_in_2_0_0;
  assign port_state_out_10_0_1 = port_state_in_2_0_1;
  assign port_state_out_10_0_2 = port_state_in_2_0_2;
  assign port_state_out_10_0_3 = port_state_in_2_0_3;
  assign port_state_out_10_0_4 = port_state_in_2_0_4;
  assign port_state_out_10_0_5 = port_state_in_2_0_5;
  assign port_state_out_10_0_6 = port_state_in_2_0_6;
  assign port_state_out_10_0_7 = port_state_in_2_0_7;
  assign port_state_out_10_1_0 = port_state_in_2_1_0;
  assign port_state_out_10_1_1 = port_state_in_2_1_1;
  assign port_state_out_10_1_2 = port_state_in_2_1_2;
  assign port_state_out_10_1_3 = port_state_in_2_1_3;
  assign port_state_out_10_1_4 = port_state_in_2_1_4;
  assign port_state_out_10_1_5 = port_state_in_2_1_5;
  assign port_state_out_10_1_6 = port_state_in_2_1_6;
  assign port_state_out_10_1_7 = port_state_in_2_1_7;
  assign port_state_out_10_2_0 = port_state_in_2_2_0;
  assign port_state_out_10_2_1 = port_state_in_2_2_1;
  assign port_state_out_10_2_2 = port_state_in_2_2_2;
  assign port_state_out_10_2_3 = port_state_in_2_2_3;
  assign port_state_out_10_2_4 = port_state_in_2_2_4;
  assign port_state_out_10_2_5 = port_state_in_2_2_5;
  assign port_state_out_10_2_6 = port_state_in_2_2_6;
  assign port_state_out_10_2_7 = port_state_in_2_2_7;
  assign port_state_out_10_3_0 = port_state_in_2_3_0;
  assign port_state_out_10_3_1 = port_state_in_2_3_1;
  assign port_state_out_10_3_2 = port_state_in_2_3_2;
  assign port_state_out_10_3_3 = port_state_in_2_3_3;
  assign port_state_out_10_3_4 = port_state_in_2_3_4;
  assign port_state_out_10_3_5 = port_state_in_2_3_5;
  assign port_state_out_10_3_6 = port_state_in_2_3_6;
  assign port_state_out_10_3_7 = port_state_in_2_3_7;
  assign port_state_out_11_0_0 = port_state_in_7_0_0;
  assign port_state_out_11_0_1 = port_state_in_7_0_1;
  assign port_state_out_11_0_2 = port_state_in_7_0_2;
  assign port_state_out_11_0_3 = port_state_in_7_0_3;
  assign port_state_out_11_0_4 = port_state_in_7_0_4;
  assign port_state_out_11_0_5 = port_state_in_7_0_5;
  assign port_state_out_11_0_6 = port_state_in_7_0_6;
  assign port_state_out_11_0_7 = port_state_in_7_0_7;
  assign port_state_out_11_1_0 = port_state_in_7_1_0;
  assign port_state_out_11_1_1 = port_state_in_7_1_1;
  assign port_state_out_11_1_2 = port_state_in_7_1_2;
  assign port_state_out_11_1_3 = port_state_in_7_1_3;
  assign port_state_out_11_1_4 = port_state_in_7_1_4;
  assign port_state_out_11_1_5 = port_state_in_7_1_5;
  assign port_state_out_11_1_6 = port_state_in_7_1_6;
  assign port_state_out_11_1_7 = port_state_in_7_1_7;
  assign port_state_out_11_2_0 = port_state_in_7_2_0;
  assign port_state_out_11_2_1 = port_state_in_7_2_1;
  assign port_state_out_11_2_2 = port_state_in_7_2_2;
  assign port_state_out_11_2_3 = port_state_in_7_2_3;
  assign port_state_out_11_2_4 = port_state_in_7_2_4;
  assign port_state_out_11_2_5 = port_state_in_7_2_5;
  assign port_state_out_11_2_6 = port_state_in_7_2_6;
  assign port_state_out_11_2_7 = port_state_in_7_2_7;
  assign port_state_out_11_3_0 = port_state_in_7_3_0;
  assign port_state_out_11_3_1 = port_state_in_7_3_1;
  assign port_state_out_11_3_2 = port_state_in_7_3_2;
  assign port_state_out_11_3_3 = port_state_in_7_3_3;
  assign port_state_out_11_3_4 = port_state_in_7_3_4;
  assign port_state_out_11_3_5 = port_state_in_7_3_5;
  assign port_state_out_11_3_6 = port_state_in_7_3_6;
  assign port_state_out_11_3_7 = port_state_in_7_3_7;
  assign port_state_out_12_0_0 = port_state_in_12_0_0;
  assign port_state_out_12_0_1 = port_state_in_12_0_1;
  assign port_state_out_12_0_2 = port_state_in_12_0_2;
  assign port_state_out_12_0_3 = port_state_in_12_0_3;
  assign port_state_out_12_0_4 = port_state_in_12_0_4;
  assign port_state_out_12_0_5 = port_state_in_12_0_5;
  assign port_state_out_12_0_6 = port_state_in_12_0_6;
  assign port_state_out_12_0_7 = port_state_in_12_0_7;
  assign port_state_out_12_1_0 = port_state_in_12_1_0;
  assign port_state_out_12_1_1 = port_state_in_12_1_1;
  assign port_state_out_12_1_2 = port_state_in_12_1_2;
  assign port_state_out_12_1_3 = port_state_in_12_1_3;
  assign port_state_out_12_1_4 = port_state_in_12_1_4;
  assign port_state_out_12_1_5 = port_state_in_12_1_5;
  assign port_state_out_12_1_6 = port_state_in_12_1_6;
  assign port_state_out_12_1_7 = port_state_in_12_1_7;
  assign port_state_out_12_2_0 = port_state_in_12_2_0;
  assign port_state_out_12_2_1 = port_state_in_12_2_1;
  assign port_state_out_12_2_2 = port_state_in_12_2_2;
  assign port_state_out_12_2_3 = port_state_in_12_2_3;
  assign port_state_out_12_2_4 = port_state_in_12_2_4;
  assign port_state_out_12_2_5 = port_state_in_12_2_5;
  assign port_state_out_12_2_6 = port_state_in_12_2_6;
  assign port_state_out_12_2_7 = port_state_in_12_2_7;
  assign port_state_out_12_3_0 = port_state_in_12_3_0;
  assign port_state_out_12_3_1 = port_state_in_12_3_1;
  assign port_state_out_12_3_2 = port_state_in_12_3_2;
  assign port_state_out_12_3_3 = port_state_in_12_3_3;
  assign port_state_out_12_3_4 = port_state_in_12_3_4;
  assign port_state_out_12_3_5 = port_state_in_12_3_5;
  assign port_state_out_12_3_6 = port_state_in_12_3_6;
  assign port_state_out_12_3_7 = port_state_in_12_3_7;
  assign port_state_out_13_0_0 = port_state_in_1_0_0;
  assign port_state_out_13_0_1 = port_state_in_1_0_1;
  assign port_state_out_13_0_2 = port_state_in_1_0_2;
  assign port_state_out_13_0_3 = port_state_in_1_0_3;
  assign port_state_out_13_0_4 = port_state_in_1_0_4;
  assign port_state_out_13_0_5 = port_state_in_1_0_5;
  assign port_state_out_13_0_6 = port_state_in_1_0_6;
  assign port_state_out_13_0_7 = port_state_in_1_0_7;
  assign port_state_out_13_1_0 = port_state_in_1_1_0;
  assign port_state_out_13_1_1 = port_state_in_1_1_1;
  assign port_state_out_13_1_2 = port_state_in_1_1_2;
  assign port_state_out_13_1_3 = port_state_in_1_1_3;
  assign port_state_out_13_1_4 = port_state_in_1_1_4;
  assign port_state_out_13_1_5 = port_state_in_1_1_5;
  assign port_state_out_13_1_6 = port_state_in_1_1_6;
  assign port_state_out_13_1_7 = port_state_in_1_1_7;
  assign port_state_out_13_2_0 = port_state_in_1_2_0;
  assign port_state_out_13_2_1 = port_state_in_1_2_1;
  assign port_state_out_13_2_2 = port_state_in_1_2_2;
  assign port_state_out_13_2_3 = port_state_in_1_2_3;
  assign port_state_out_13_2_4 = port_state_in_1_2_4;
  assign port_state_out_13_2_5 = port_state_in_1_2_5;
  assign port_state_out_13_2_6 = port_state_in_1_2_6;
  assign port_state_out_13_2_7 = port_state_in_1_2_7;
  assign port_state_out_13_3_0 = port_state_in_1_3_0;
  assign port_state_out_13_3_1 = port_state_in_1_3_1;
  assign port_state_out_13_3_2 = port_state_in_1_3_2;
  assign port_state_out_13_3_3 = port_state_in_1_3_3;
  assign port_state_out_13_3_4 = port_state_in_1_3_4;
  assign port_state_out_13_3_5 = port_state_in_1_3_5;
  assign port_state_out_13_3_6 = port_state_in_1_3_6;
  assign port_state_out_13_3_7 = port_state_in_1_3_7;
  assign port_state_out_14_0_0 = port_state_in_6_0_0;
  assign port_state_out_14_0_1 = port_state_in_6_0_1;
  assign port_state_out_14_0_2 = port_state_in_6_0_2;
  assign port_state_out_14_0_3 = port_state_in_6_0_3;
  assign port_state_out_14_0_4 = port_state_in_6_0_4;
  assign port_state_out_14_0_5 = port_state_in_6_0_5;
  assign port_state_out_14_0_6 = port_state_in_6_0_6;
  assign port_state_out_14_0_7 = port_state_in_6_0_7;
  assign port_state_out_14_1_0 = port_state_in_6_1_0;
  assign port_state_out_14_1_1 = port_state_in_6_1_1;
  assign port_state_out_14_1_2 = port_state_in_6_1_2;
  assign port_state_out_14_1_3 = port_state_in_6_1_3;
  assign port_state_out_14_1_4 = port_state_in_6_1_4;
  assign port_state_out_14_1_5 = port_state_in_6_1_5;
  assign port_state_out_14_1_6 = port_state_in_6_1_6;
  assign port_state_out_14_1_7 = port_state_in_6_1_7;
  assign port_state_out_14_2_0 = port_state_in_6_2_0;
  assign port_state_out_14_2_1 = port_state_in_6_2_1;
  assign port_state_out_14_2_2 = port_state_in_6_2_2;
  assign port_state_out_14_2_3 = port_state_in_6_2_3;
  assign port_state_out_14_2_4 = port_state_in_6_2_4;
  assign port_state_out_14_2_5 = port_state_in_6_2_5;
  assign port_state_out_14_2_6 = port_state_in_6_2_6;
  assign port_state_out_14_2_7 = port_state_in_6_2_7;
  assign port_state_out_14_3_0 = port_state_in_6_3_0;
  assign port_state_out_14_3_1 = port_state_in_6_3_1;
  assign port_state_out_14_3_2 = port_state_in_6_3_2;
  assign port_state_out_14_3_3 = port_state_in_6_3_3;
  assign port_state_out_14_3_4 = port_state_in_6_3_4;
  assign port_state_out_14_3_5 = port_state_in_6_3_5;
  assign port_state_out_14_3_6 = port_state_in_6_3_6;
  assign port_state_out_14_3_7 = port_state_in_6_3_7;
  assign port_state_out_15_0_0 = port_state_in_11_0_0;
  assign port_state_out_15_0_1 = port_state_in_11_0_1;
  assign port_state_out_15_0_2 = port_state_in_11_0_2;
  assign port_state_out_15_0_3 = port_state_in_11_0_3;
  assign port_state_out_15_0_4 = port_state_in_11_0_4;
  assign port_state_out_15_0_5 = port_state_in_11_0_5;
  assign port_state_out_15_0_6 = port_state_in_11_0_6;
  assign port_state_out_15_0_7 = port_state_in_11_0_7;
  assign port_state_out_15_1_0 = port_state_in_11_1_0;
  assign port_state_out_15_1_1 = port_state_in_11_1_1;
  assign port_state_out_15_1_2 = port_state_in_11_1_2;
  assign port_state_out_15_1_3 = port_state_in_11_1_3;
  assign port_state_out_15_1_4 = port_state_in_11_1_4;
  assign port_state_out_15_1_5 = port_state_in_11_1_5;
  assign port_state_out_15_1_6 = port_state_in_11_1_6;
  assign port_state_out_15_1_7 = port_state_in_11_1_7;
  assign port_state_out_15_2_0 = port_state_in_11_2_0;
  assign port_state_out_15_2_1 = port_state_in_11_2_1;
  assign port_state_out_15_2_2 = port_state_in_11_2_2;
  assign port_state_out_15_2_3 = port_state_in_11_2_3;
  assign port_state_out_15_2_4 = port_state_in_11_2_4;
  assign port_state_out_15_2_5 = port_state_in_11_2_5;
  assign port_state_out_15_2_6 = port_state_in_11_2_6;
  assign port_state_out_15_2_7 = port_state_in_11_2_7;
  assign port_state_out_15_3_0 = port_state_in_11_3_0;
  assign port_state_out_15_3_1 = port_state_in_11_3_1;
  assign port_state_out_15_3_2 = port_state_in_11_3_2;
  assign port_state_out_15_3_3 = port_state_in_11_3_3;
  assign port_state_out_15_3_4 = port_state_in_11_3_4;
  assign port_state_out_15_3_5 = port_state_in_11_3_5;
  assign port_state_out_15_3_6 = port_state_in_11_3_6;
  assign port_state_out_15_3_7 = port_state_in_11_3_7;

endmodule

//Sbox_AES_BoyarPeralta replaced by Sbox_AES_BoyarPeralta

//Sbox_AES_BoyarPeralta replaced by Sbox_AES_BoyarPeralta

//Sbox_AES_BoyarPeralta replaced by Sbox_AES_BoyarPeralta

//Sbox_AES_BoyarPeralta replaced by Sbox_AES_BoyarPeralta

//Sbox_AES_BoyarPeralta replaced by Sbox_AES_BoyarPeralta

//Sbox_AES_BoyarPeralta replaced by Sbox_AES_BoyarPeralta

//Sbox_AES_BoyarPeralta replaced by Sbox_AES_BoyarPeralta

//Sbox_AES_BoyarPeralta replaced by Sbox_AES_BoyarPeralta

//Sbox_AES_BoyarPeralta replaced by Sbox_AES_BoyarPeralta

//Sbox_AES_BoyarPeralta replaced by Sbox_AES_BoyarPeralta

//Sbox_AES_BoyarPeralta replaced by Sbox_AES_BoyarPeralta

//Sbox_AES_BoyarPeralta replaced by Sbox_AES_BoyarPeralta

//Sbox_AES_BoyarPeralta replaced by Sbox_AES_BoyarPeralta

//Sbox_AES_BoyarPeralta replaced by Sbox_AES_BoyarPeralta

//Sbox_AES_BoyarPeralta replaced by Sbox_AES_BoyarPeralta

module Sbox_AES_BoyarPeralta (
  input      [0:0]    port_i_0_0,
  input      [0:0]    port_i_0_1,
  input      [0:0]    port_i_0_2,
  input      [0:0]    port_i_0_3,
  input      [0:0]    port_i_0_4,
  input      [0:0]    port_i_0_5,
  input      [0:0]    port_i_0_6,
  input      [0:0]    port_i_0_7,
  input      [0:0]    port_i_1_0,
  input      [0:0]    port_i_1_1,
  input      [0:0]    port_i_1_2,
  input      [0:0]    port_i_1_3,
  input      [0:0]    port_i_1_4,
  input      [0:0]    port_i_1_5,
  input      [0:0]    port_i_1_6,
  input      [0:0]    port_i_1_7,
  input      [0:0]    port_i_2_0,
  input      [0:0]    port_i_2_1,
  input      [0:0]    port_i_2_2,
  input      [0:0]    port_i_2_3,
  input      [0:0]    port_i_2_4,
  input      [0:0]    port_i_2_5,
  input      [0:0]    port_i_2_6,
  input      [0:0]    port_i_2_7,
  input      [0:0]    port_i_3_0,
  input      [0:0]    port_i_3_1,
  input      [0:0]    port_i_3_2,
  input      [0:0]    port_i_3_3,
  input      [0:0]    port_i_3_4,
  input      [0:0]    port_i_3_5,
  input      [0:0]    port_i_3_6,
  input      [0:0]    port_i_3_7,
  output     [0:0]    port_o_0_0,
  output     [0:0]    port_o_0_1,
  output     [0:0]    port_o_0_2,
  output     [0:0]    port_o_0_3,
  output     [0:0]    port_o_0_4,
  output     [0:0]    port_o_0_5,
  output     [0:0]    port_o_0_6,
  output     [0:0]    port_o_0_7,
  output     [0:0]    port_o_1_0,
  output     [0:0]    port_o_1_1,
  output     [0:0]    port_o_1_2,
  output     [0:0]    port_o_1_3,
  output     [0:0]    port_o_1_4,
  output     [0:0]    port_o_1_5,
  output     [0:0]    port_o_1_6,
  output     [0:0]    port_o_1_7,
  output     [0:0]    port_o_2_0,
  output     [0:0]    port_o_2_1,
  output     [0:0]    port_o_2_2,
  output     [0:0]    port_o_2_3,
  output     [0:0]    port_o_2_4,
  output     [0:0]    port_o_2_5,
  output     [0:0]    port_o_2_6,
  output     [0:0]    port_o_2_7,
  output     [0:0]    port_o_3_0,
  output     [0:0]    port_o_3_1,
  output     [0:0]    port_o_3_2,
  output     [0:0]    port_o_3_3,
  output     [0:0]    port_o_3_4,
  output     [0:0]    port_o_3_5,
  output     [0:0]    port_o_3_6,
  output     [0:0]    port_o_3_7,
  input               clk,
  input               reset
);

  wire       [0:0]    t1_xor_port_y_0;
  wire       [0:0]    t1_xor_port_y_1;
  wire       [0:0]    t1_xor_port_y_2;
  wire       [0:0]    t1_xor_port_y_3;
  wire       [0:0]    t2_xor_port_y_0;
  wire       [0:0]    t2_xor_port_y_1;
  wire       [0:0]    t2_xor_port_y_2;
  wire       [0:0]    t2_xor_port_y_3;
  wire       [0:0]    t3_xor_port_y_0;
  wire       [0:0]    t3_xor_port_y_1;
  wire       [0:0]    t3_xor_port_y_2;
  wire       [0:0]    t3_xor_port_y_3;
  wire       [0:0]    t4_xor_port_y_0;
  wire       [0:0]    t4_xor_port_y_1;
  wire       [0:0]    t4_xor_port_y_2;
  wire       [0:0]    t4_xor_port_y_3;
  wire       [0:0]    t5_xor_port_y_0;
  wire       [0:0]    t5_xor_port_y_1;
  wire       [0:0]    t5_xor_port_y_2;
  wire       [0:0]    t5_xor_port_y_3;
  wire       [0:0]    t6_xor_port_y_0;
  wire       [0:0]    t6_xor_port_y_1;
  wire       [0:0]    t6_xor_port_y_2;
  wire       [0:0]    t6_xor_port_y_3;
  wire       [0:0]    t7_xor_port_y_0;
  wire       [0:0]    t7_xor_port_y_1;
  wire       [0:0]    t7_xor_port_y_2;
  wire       [0:0]    t7_xor_port_y_3;
  wire       [0:0]    t8_xor_port_y_0;
  wire       [0:0]    t8_xor_port_y_1;
  wire       [0:0]    t8_xor_port_y_2;
  wire       [0:0]    t8_xor_port_y_3;
  wire       [0:0]    t9_xor_port_y_0;
  wire       [0:0]    t9_xor_port_y_1;
  wire       [0:0]    t9_xor_port_y_2;
  wire       [0:0]    t9_xor_port_y_3;
  wire       [0:0]    t10_xor_port_y_0;
  wire       [0:0]    t10_xor_port_y_1;
  wire       [0:0]    t10_xor_port_y_2;
  wire       [0:0]    t10_xor_port_y_3;
  wire       [0:0]    t11_xor_port_y_0;
  wire       [0:0]    t11_xor_port_y_1;
  wire       [0:0]    t11_xor_port_y_2;
  wire       [0:0]    t11_xor_port_y_3;
  wire       [0:0]    t12_xor_port_y_0;
  wire       [0:0]    t12_xor_port_y_1;
  wire       [0:0]    t12_xor_port_y_2;
  wire       [0:0]    t12_xor_port_y_3;
  wire       [0:0]    t13_xor_port_y_0;
  wire       [0:0]    t13_xor_port_y_1;
  wire       [0:0]    t13_xor_port_y_2;
  wire       [0:0]    t13_xor_port_y_3;
  wire       [0:0]    t14_xor_port_y_0;
  wire       [0:0]    t14_xor_port_y_1;
  wire       [0:0]    t14_xor_port_y_2;
  wire       [0:0]    t14_xor_port_y_3;
  wire       [0:0]    t15_xor_port_y_0;
  wire       [0:0]    t15_xor_port_y_1;
  wire       [0:0]    t15_xor_port_y_2;
  wire       [0:0]    t15_xor_port_y_3;
  wire       [0:0]    t16_xor_port_y_0;
  wire       [0:0]    t16_xor_port_y_1;
  wire       [0:0]    t16_xor_port_y_2;
  wire       [0:0]    t16_xor_port_y_3;
  wire       [0:0]    t17_xor_port_y_0;
  wire       [0:0]    t17_xor_port_y_1;
  wire       [0:0]    t17_xor_port_y_2;
  wire       [0:0]    t17_xor_port_y_3;
  wire       [0:0]    t18_xor_port_y_0;
  wire       [0:0]    t18_xor_port_y_1;
  wire       [0:0]    t18_xor_port_y_2;
  wire       [0:0]    t18_xor_port_y_3;
  wire       [0:0]    t19_xor_port_y_0;
  wire       [0:0]    t19_xor_port_y_1;
  wire       [0:0]    t19_xor_port_y_2;
  wire       [0:0]    t19_xor_port_y_3;
  wire       [0:0]    t20_xor_port_y_0;
  wire       [0:0]    t20_xor_port_y_1;
  wire       [0:0]    t20_xor_port_y_2;
  wire       [0:0]    t20_xor_port_y_3;
  wire       [0:0]    t21_xor_port_y_0;
  wire       [0:0]    t21_xor_port_y_1;
  wire       [0:0]    t21_xor_port_y_2;
  wire       [0:0]    t21_xor_port_y_3;
  wire       [0:0]    t22_xor_port_y_0;
  wire       [0:0]    t22_xor_port_y_1;
  wire       [0:0]    t22_xor_port_y_2;
  wire       [0:0]    t22_xor_port_y_3;
  wire       [0:0]    t23_xor_port_y_0;
  wire       [0:0]    t23_xor_port_y_1;
  wire       [0:0]    t23_xor_port_y_2;
  wire       [0:0]    t23_xor_port_y_3;
  wire       [0:0]    t24_xor_port_y_0;
  wire       [0:0]    t24_xor_port_y_1;
  wire       [0:0]    t24_xor_port_y_2;
  wire       [0:0]    t24_xor_port_y_3;
  wire       [0:0]    t25_xor_port_y_0;
  wire       [0:0]    t25_xor_port_y_1;
  wire       [0:0]    t25_xor_port_y_2;
  wire       [0:0]    t25_xor_port_y_3;
  wire       [0:0]    t26_xor_port_y_0;
  wire       [0:0]    t26_xor_port_y_1;
  wire       [0:0]    t26_xor_port_y_2;
  wire       [0:0]    t26_xor_port_y_3;
  wire       [0:0]    t27_xor_port_y_0;
  wire       [0:0]    t27_xor_port_y_1;
  wire       [0:0]    t27_xor_port_y_2;
  wire       [0:0]    t27_xor_port_y_3;
  wire       [0:0]    m1_port_y_0;
  wire       [0:0]    m1_port_y_1;
  wire       [0:0]    m1_port_y_2;
  wire       [0:0]    m1_port_y_3;
  wire       [0:0]    m2_port_y_0;
  wire       [0:0]    m2_port_y_1;
  wire       [0:0]    m2_port_y_2;
  wire       [0:0]    m2_port_y_3;
  wire       [0:0]    m4_port_y_0;
  wire       [0:0]    m4_port_y_1;
  wire       [0:0]    m4_port_y_2;
  wire       [0:0]    m4_port_y_3;
  wire       [0:0]    m6_port_y_0;
  wire       [0:0]    m6_port_y_1;
  wire       [0:0]    m6_port_y_2;
  wire       [0:0]    m6_port_y_3;
  wire       [0:0]    m7_port_y_0;
  wire       [0:0]    m7_port_y_1;
  wire       [0:0]    m7_port_y_2;
  wire       [0:0]    m7_port_y_3;
  wire       [0:0]    m9_port_y_0;
  wire       [0:0]    m9_port_y_1;
  wire       [0:0]    m9_port_y_2;
  wire       [0:0]    m9_port_y_3;
  wire       [0:0]    m11_port_y_0;
  wire       [0:0]    m11_port_y_1;
  wire       [0:0]    m11_port_y_2;
  wire       [0:0]    m11_port_y_3;
  wire       [0:0]    m12_port_y_0;
  wire       [0:0]    m12_port_y_1;
  wire       [0:0]    m12_port_y_2;
  wire       [0:0]    m12_port_y_3;
  wire       [0:0]    m14_port_y_0;
  wire       [0:0]    m14_port_y_1;
  wire       [0:0]    m14_port_y_2;
  wire       [0:0]    m14_port_y_3;
  wire       [0:0]    m3_xor_port_y_0;
  wire       [0:0]    m3_xor_port_y_1;
  wire       [0:0]    m3_xor_port_y_2;
  wire       [0:0]    m3_xor_port_y_3;
  wire       [0:0]    m5_xor_port_y_0;
  wire       [0:0]    m5_xor_port_y_1;
  wire       [0:0]    m5_xor_port_y_2;
  wire       [0:0]    m5_xor_port_y_3;
  wire       [0:0]    m8_xor_port_y_0;
  wire       [0:0]    m8_xor_port_y_1;
  wire       [0:0]    m8_xor_port_y_2;
  wire       [0:0]    m8_xor_port_y_3;
  wire       [0:0]    m10_xor_port_y_0;
  wire       [0:0]    m10_xor_port_y_1;
  wire       [0:0]    m10_xor_port_y_2;
  wire       [0:0]    m10_xor_port_y_3;
  wire       [0:0]    m13_xor_port_y_0;
  wire       [0:0]    m13_xor_port_y_1;
  wire       [0:0]    m13_xor_port_y_2;
  wire       [0:0]    m13_xor_port_y_3;
  wire       [0:0]    m15_xor_port_y_0;
  wire       [0:0]    m15_xor_port_y_1;
  wire       [0:0]    m15_xor_port_y_2;
  wire       [0:0]    m15_xor_port_y_3;
  wire       [0:0]    m16_xor_port_y_0;
  wire       [0:0]    m16_xor_port_y_1;
  wire       [0:0]    m16_xor_port_y_2;
  wire       [0:0]    m16_xor_port_y_3;
  wire       [0:0]    m17_xor_port_y_0;
  wire       [0:0]    m17_xor_port_y_1;
  wire       [0:0]    m17_xor_port_y_2;
  wire       [0:0]    m17_xor_port_y_3;
  wire       [0:0]    m18_xor_port_y_0;
  wire       [0:0]    m18_xor_port_y_1;
  wire       [0:0]    m18_xor_port_y_2;
  wire       [0:0]    m18_xor_port_y_3;
  wire       [0:0]    m19_xor_port_y_0;
  wire       [0:0]    m19_xor_port_y_1;
  wire       [0:0]    m19_xor_port_y_2;
  wire       [0:0]    m19_xor_port_y_3;
  wire       [0:0]    m20_xor_port_y_0;
  wire       [0:0]    m20_xor_port_y_1;
  wire       [0:0]    m20_xor_port_y_2;
  wire       [0:0]    m20_xor_port_y_3;
  wire       [0:0]    m21_xor_port_y_0;
  wire       [0:0]    m21_xor_port_y_1;
  wire       [0:0]    m21_xor_port_y_2;
  wire       [0:0]    m21_xor_port_y_3;
  wire       [0:0]    m22_xor_port_y_0;
  wire       [0:0]    m22_xor_port_y_1;
  wire       [0:0]    m22_xor_port_y_2;
  wire       [0:0]    m22_xor_port_y_3;
  wire       [0:0]    m23_xor_port_y_0;
  wire       [0:0]    m23_xor_port_y_1;
  wire       [0:0]    m23_xor_port_y_2;
  wire       [0:0]    m23_xor_port_y_3;
  wire       [0:0]    m24_xor_port_y_0;
  wire       [0:0]    m24_xor_port_y_1;
  wire       [0:0]    m24_xor_port_y_2;
  wire       [0:0]    m24_xor_port_y_3;
  wire       [0:0]    m25_port_y_0;
  wire       [0:0]    m25_port_y_1;
  wire       [0:0]    m25_port_y_2;
  wire       [0:0]    m25_port_y_3;
  wire       [0:0]    m27_xor_port_y_0;
  wire       [0:0]    m27_xor_port_y_1;
  wire       [0:0]    m27_xor_port_y_2;
  wire       [0:0]    m27_xor_port_y_3;
  wire       [0:0]    m31_port_y_0;
  wire       [0:0]    m31_port_y_1;
  wire       [0:0]    m31_port_y_2;
  wire       [0:0]    m31_port_y_3;
  wire       [0:0]    m34_port_y_0;
  wire       [0:0]    m34_port_y_1;
  wire       [0:0]    m34_port_y_2;
  wire       [0:0]    m34_port_y_3;
  wire       [0:0]    m26_xor_port_y_0;
  wire       [0:0]    m26_xor_port_y_1;
  wire       [0:0]    m26_xor_port_y_2;
  wire       [0:0]    m26_xor_port_y_3;
  wire       [0:0]    m28_xor_port_y_0;
  wire       [0:0]    m28_xor_port_y_1;
  wire       [0:0]    m28_xor_port_y_2;
  wire       [0:0]    m28_xor_port_y_3;
  wire       [0:0]    m29_port_y_0;
  wire       [0:0]    m29_port_y_1;
  wire       [0:0]    m29_port_y_2;
  wire       [0:0]    m29_port_y_3;
  wire       [0:0]    m30_port_y_0;
  wire       [0:0]    m30_port_y_1;
  wire       [0:0]    m30_port_y_2;
  wire       [0:0]    m30_port_y_3;
  wire       [0:0]    m32_port_y_0;
  wire       [0:0]    m32_port_y_1;
  wire       [0:0]    m32_port_y_2;
  wire       [0:0]    m32_port_y_3;
  wire       [0:0]    m33_xor_port_y_0;
  wire       [0:0]    m33_xor_port_y_1;
  wire       [0:0]    m33_xor_port_y_2;
  wire       [0:0]    m33_xor_port_y_3;
  wire       [0:0]    m35_port_y_0;
  wire       [0:0]    m35_port_y_1;
  wire       [0:0]    m35_port_y_2;
  wire       [0:0]    m35_port_y_3;
  wire       [0:0]    m36_xor_port_y_0;
  wire       [0:0]    m36_xor_port_y_1;
  wire       [0:0]    m36_xor_port_y_2;
  wire       [0:0]    m36_xor_port_y_3;
  wire       [0:0]    m37_xor_port_y_0;
  wire       [0:0]    m37_xor_port_y_1;
  wire       [0:0]    m37_xor_port_y_2;
  wire       [0:0]    m37_xor_port_y_3;
  wire       [0:0]    m38_xor_port_y_0;
  wire       [0:0]    m38_xor_port_y_1;
  wire       [0:0]    m38_xor_port_y_2;
  wire       [0:0]    m38_xor_port_y_3;
  wire       [0:0]    m39_xor_port_y_0;
  wire       [0:0]    m39_xor_port_y_1;
  wire       [0:0]    m39_xor_port_y_2;
  wire       [0:0]    m39_xor_port_y_3;
  wire       [0:0]    m40_xor_port_y_0;
  wire       [0:0]    m40_xor_port_y_1;
  wire       [0:0]    m40_xor_port_y_2;
  wire       [0:0]    m40_xor_port_y_3;
  wire       [0:0]    m41_xor_port_y_0;
  wire       [0:0]    m41_xor_port_y_1;
  wire       [0:0]    m41_xor_port_y_2;
  wire       [0:0]    m41_xor_port_y_3;
  wire       [0:0]    m42_xor_port_y_0;
  wire       [0:0]    m42_xor_port_y_1;
  wire       [0:0]    m42_xor_port_y_2;
  wire       [0:0]    m42_xor_port_y_3;
  wire       [0:0]    m43_xor_port_y_0;
  wire       [0:0]    m43_xor_port_y_1;
  wire       [0:0]    m43_xor_port_y_2;
  wire       [0:0]    m43_xor_port_y_3;
  wire       [0:0]    m44_xor_port_y_0;
  wire       [0:0]    m44_xor_port_y_1;
  wire       [0:0]    m44_xor_port_y_2;
  wire       [0:0]    m44_xor_port_y_3;
  wire       [0:0]    m45_xor_port_y_0;
  wire       [0:0]    m45_xor_port_y_1;
  wire       [0:0]    m45_xor_port_y_2;
  wire       [0:0]    m45_xor_port_y_3;
  wire       [0:0]    m46_mul_port_y_0;
  wire       [0:0]    m46_mul_port_y_1;
  wire       [0:0]    m46_mul_port_y_2;
  wire       [0:0]    m46_mul_port_y_3;
  wire       [0:0]    m47_mul_port_y_0;
  wire       [0:0]    m47_mul_port_y_1;
  wire       [0:0]    m47_mul_port_y_2;
  wire       [0:0]    m47_mul_port_y_3;
  wire       [0:0]    m48_mul_port_y_0;
  wire       [0:0]    m48_mul_port_y_1;
  wire       [0:0]    m48_mul_port_y_2;
  wire       [0:0]    m48_mul_port_y_3;
  wire       [0:0]    m49_mul_port_y_0;
  wire       [0:0]    m49_mul_port_y_1;
  wire       [0:0]    m49_mul_port_y_2;
  wire       [0:0]    m49_mul_port_y_3;
  wire       [0:0]    m50_mul_port_y_0;
  wire       [0:0]    m50_mul_port_y_1;
  wire       [0:0]    m50_mul_port_y_2;
  wire       [0:0]    m50_mul_port_y_3;
  wire       [0:0]    m51_mul_port_y_0;
  wire       [0:0]    m51_mul_port_y_1;
  wire       [0:0]    m51_mul_port_y_2;
  wire       [0:0]    m51_mul_port_y_3;
  wire       [0:0]    m52_mul_port_y_0;
  wire       [0:0]    m52_mul_port_y_1;
  wire       [0:0]    m52_mul_port_y_2;
  wire       [0:0]    m52_mul_port_y_3;
  wire       [0:0]    m53_mul_port_y_0;
  wire       [0:0]    m53_mul_port_y_1;
  wire       [0:0]    m53_mul_port_y_2;
  wire       [0:0]    m53_mul_port_y_3;
  wire       [0:0]    m54_mul_port_y_0;
  wire       [0:0]    m54_mul_port_y_1;
  wire       [0:0]    m54_mul_port_y_2;
  wire       [0:0]    m54_mul_port_y_3;
  wire       [0:0]    m55_mul_port_y_0;
  wire       [0:0]    m55_mul_port_y_1;
  wire       [0:0]    m55_mul_port_y_2;
  wire       [0:0]    m55_mul_port_y_3;
  wire       [0:0]    m56_mul_port_y_0;
  wire       [0:0]    m56_mul_port_y_1;
  wire       [0:0]    m56_mul_port_y_2;
  wire       [0:0]    m56_mul_port_y_3;
  wire       [0:0]    m57_mul_port_y_0;
  wire       [0:0]    m57_mul_port_y_1;
  wire       [0:0]    m57_mul_port_y_2;
  wire       [0:0]    m57_mul_port_y_3;
  wire       [0:0]    m58_mul_port_y_0;
  wire       [0:0]    m58_mul_port_y_1;
  wire       [0:0]    m58_mul_port_y_2;
  wire       [0:0]    m58_mul_port_y_3;
  wire       [0:0]    m59_mul_port_y_0;
  wire       [0:0]    m59_mul_port_y_1;
  wire       [0:0]    m59_mul_port_y_2;
  wire       [0:0]    m59_mul_port_y_3;
  wire       [0:0]    m60_mul_port_y_0;
  wire       [0:0]    m60_mul_port_y_1;
  wire       [0:0]    m60_mul_port_y_2;
  wire       [0:0]    m60_mul_port_y_3;
  wire       [0:0]    m61_mul_port_y_0;
  wire       [0:0]    m61_mul_port_y_1;
  wire       [0:0]    m61_mul_port_y_2;
  wire       [0:0]    m61_mul_port_y_3;
  wire       [0:0]    m62_mul_port_y_0;
  wire       [0:0]    m62_mul_port_y_1;
  wire       [0:0]    m62_mul_port_y_2;
  wire       [0:0]    m62_mul_port_y_3;
  wire       [0:0]    m63_mul_port_y_0;
  wire       [0:0]    m63_mul_port_y_1;
  wire       [0:0]    m63_mul_port_y_2;
  wire       [0:0]    m63_mul_port_y_3;
  wire       [0:0]    l0_xor_port_y_0;
  wire       [0:0]    l0_xor_port_y_1;
  wire       [0:0]    l0_xor_port_y_2;
  wire       [0:0]    l0_xor_port_y_3;
  wire       [0:0]    l1_xor_port_y_0;
  wire       [0:0]    l1_xor_port_y_1;
  wire       [0:0]    l1_xor_port_y_2;
  wire       [0:0]    l1_xor_port_y_3;
  wire       [0:0]    l2_xor_port_y_0;
  wire       [0:0]    l2_xor_port_y_1;
  wire       [0:0]    l2_xor_port_y_2;
  wire       [0:0]    l2_xor_port_y_3;
  wire       [0:0]    l3_xor_port_y_0;
  wire       [0:0]    l3_xor_port_y_1;
  wire       [0:0]    l3_xor_port_y_2;
  wire       [0:0]    l3_xor_port_y_3;
  wire       [0:0]    l4_xor_port_y_0;
  wire       [0:0]    l4_xor_port_y_1;
  wire       [0:0]    l4_xor_port_y_2;
  wire       [0:0]    l4_xor_port_y_3;
  wire       [0:0]    l5_xor_port_y_0;
  wire       [0:0]    l5_xor_port_y_1;
  wire       [0:0]    l5_xor_port_y_2;
  wire       [0:0]    l5_xor_port_y_3;
  wire       [0:0]    l6_xor_port_y_0;
  wire       [0:0]    l6_xor_port_y_1;
  wire       [0:0]    l6_xor_port_y_2;
  wire       [0:0]    l6_xor_port_y_3;
  wire       [0:0]    l7_xor_port_y_0;
  wire       [0:0]    l7_xor_port_y_1;
  wire       [0:0]    l7_xor_port_y_2;
  wire       [0:0]    l7_xor_port_y_3;
  wire       [0:0]    l8_xor_port_y_0;
  wire       [0:0]    l8_xor_port_y_1;
  wire       [0:0]    l8_xor_port_y_2;
  wire       [0:0]    l8_xor_port_y_3;
  wire       [0:0]    l9_xor_port_y_0;
  wire       [0:0]    l9_xor_port_y_1;
  wire       [0:0]    l9_xor_port_y_2;
  wire       [0:0]    l9_xor_port_y_3;
  wire       [0:0]    l10_xor_port_y_0;
  wire       [0:0]    l10_xor_port_y_1;
  wire       [0:0]    l10_xor_port_y_2;
  wire       [0:0]    l10_xor_port_y_3;
  wire       [0:0]    l11_xor_port_y_0;
  wire       [0:0]    l11_xor_port_y_1;
  wire       [0:0]    l11_xor_port_y_2;
  wire       [0:0]    l11_xor_port_y_3;
  wire       [0:0]    l12_xor_port_y_0;
  wire       [0:0]    l12_xor_port_y_1;
  wire       [0:0]    l12_xor_port_y_2;
  wire       [0:0]    l12_xor_port_y_3;
  wire       [0:0]    l13_xor_port_y_0;
  wire       [0:0]    l13_xor_port_y_1;
  wire       [0:0]    l13_xor_port_y_2;
  wire       [0:0]    l13_xor_port_y_3;
  wire       [0:0]    l14_xor_port_y_0;
  wire       [0:0]    l14_xor_port_y_1;
  wire       [0:0]    l14_xor_port_y_2;
  wire       [0:0]    l14_xor_port_y_3;
  wire       [0:0]    l15_xor_port_y_0;
  wire       [0:0]    l15_xor_port_y_1;
  wire       [0:0]    l15_xor_port_y_2;
  wire       [0:0]    l15_xor_port_y_3;
  wire       [0:0]    l16_xor_port_y_0;
  wire       [0:0]    l16_xor_port_y_1;
  wire       [0:0]    l16_xor_port_y_2;
  wire       [0:0]    l16_xor_port_y_3;
  wire       [0:0]    l17_xor_port_y_0;
  wire       [0:0]    l17_xor_port_y_1;
  wire       [0:0]    l17_xor_port_y_2;
  wire       [0:0]    l17_xor_port_y_3;
  wire       [0:0]    l18_xor_port_y_0;
  wire       [0:0]    l18_xor_port_y_1;
  wire       [0:0]    l18_xor_port_y_2;
  wire       [0:0]    l18_xor_port_y_3;
  wire       [0:0]    l19_xor_port_y_0;
  wire       [0:0]    l19_xor_port_y_1;
  wire       [0:0]    l19_xor_port_y_2;
  wire       [0:0]    l19_xor_port_y_3;
  wire       [0:0]    l20_xor_port_y_0;
  wire       [0:0]    l20_xor_port_y_1;
  wire       [0:0]    l20_xor_port_y_2;
  wire       [0:0]    l20_xor_port_y_3;
  wire       [0:0]    l21_xor_port_y_0;
  wire       [0:0]    l21_xor_port_y_1;
  wire       [0:0]    l21_xor_port_y_2;
  wire       [0:0]    l21_xor_port_y_3;
  wire       [0:0]    l22_xor_port_y_0;
  wire       [0:0]    l22_xor_port_y_1;
  wire       [0:0]    l22_xor_port_y_2;
  wire       [0:0]    l22_xor_port_y_3;
  wire       [0:0]    l23_xor_port_y_0;
  wire       [0:0]    l23_xor_port_y_1;
  wire       [0:0]    l23_xor_port_y_2;
  wire       [0:0]    l23_xor_port_y_3;
  wire       [0:0]    l24_xor_port_y_0;
  wire       [0:0]    l24_xor_port_y_1;
  wire       [0:0]    l24_xor_port_y_2;
  wire       [0:0]    l24_xor_port_y_3;
  wire       [0:0]    l25_xor_port_y_0;
  wire       [0:0]    l25_xor_port_y_1;
  wire       [0:0]    l25_xor_port_y_2;
  wire       [0:0]    l25_xor_port_y_3;
  wire       [0:0]    l26_xor_port_y_0;
  wire       [0:0]    l26_xor_port_y_1;
  wire       [0:0]    l26_xor_port_y_2;
  wire       [0:0]    l26_xor_port_y_3;
  wire       [0:0]    l27_xor_port_y_0;
  wire       [0:0]    l27_xor_port_y_1;
  wire       [0:0]    l27_xor_port_y_2;
  wire       [0:0]    l27_xor_port_y_3;
  wire       [0:0]    l28_xor_port_y_0;
  wire       [0:0]    l28_xor_port_y_1;
  wire       [0:0]    l28_xor_port_y_2;
  wire       [0:0]    l28_xor_port_y_3;
  wire       [0:0]    l29_xor_port_y_0;
  wire       [0:0]    l29_xor_port_y_1;
  wire       [0:0]    l29_xor_port_y_2;
  wire       [0:0]    l29_xor_port_y_3;
  wire       [0:0]    s0_port_y_0;
  wire       [0:0]    s0_port_y_1;
  wire       [0:0]    s0_port_y_2;
  wire       [0:0]    s0_port_y_3;
  wire       [0:0]    s1_port_y_0;
  wire       [0:0]    s1_port_y_1;
  wire       [0:0]    s1_port_y_2;
  wire       [0:0]    s1_port_y_3;
  wire       [0:0]    s2_port_y_0;
  wire       [0:0]    s2_port_y_1;
  wire       [0:0]    s2_port_y_2;
  wire       [0:0]    s2_port_y_3;
  wire       [0:0]    s3_port_y_0;
  wire       [0:0]    s3_port_y_1;
  wire       [0:0]    s3_port_y_2;
  wire       [0:0]    s3_port_y_3;
  wire       [0:0]    s4_port_y_0;
  wire       [0:0]    s4_port_y_1;
  wire       [0:0]    s4_port_y_2;
  wire       [0:0]    s4_port_y_3;
  wire       [0:0]    s5_port_y_0;
  wire       [0:0]    s5_port_y_1;
  wire       [0:0]    s5_port_y_2;
  wire       [0:0]    s5_port_y_3;
  wire       [0:0]    s6_port_y_0;
  wire       [0:0]    s6_port_y_1;
  wire       [0:0]    s6_port_y_2;
  wire       [0:0]    s6_port_y_3;
  wire       [0:0]    s7_port_y_0;
  wire       [0:0]    s7_port_y_1;
  wire       [0:0]    s7_port_y_2;
  wire       [0:0]    s7_port_y_3;
  wire       [0:0]    in_x0_0;
  wire       [0:0]    in_x0_1;
  wire       [0:0]    in_x0_2;
  wire       [0:0]    in_x0_3;
  wire       [0:0]    in_x1_0;
  wire       [0:0]    in_x1_1;
  wire       [0:0]    in_x1_2;
  wire       [0:0]    in_x1_3;
  wire       [0:0]    in_x2_0;
  wire       [0:0]    in_x2_1;
  wire       [0:0]    in_x2_2;
  wire       [0:0]    in_x2_3;
  wire       [0:0]    in_x3_0;
  wire       [0:0]    in_x3_1;
  wire       [0:0]    in_x3_2;
  wire       [0:0]    in_x3_3;
  wire       [0:0]    in_x4_0;
  wire       [0:0]    in_x4_1;
  wire       [0:0]    in_x4_2;
  wire       [0:0]    in_x4_3;
  wire       [0:0]    in_x5_0;
  wire       [0:0]    in_x5_1;
  wire       [0:0]    in_x5_2;
  wire       [0:0]    in_x5_3;
  wire       [0:0]    in_x6_0;
  wire       [0:0]    in_x6_1;
  wire       [0:0]    in_x6_2;
  wire       [0:0]    in_x6_3;
  wire       [0:0]    in_x7_0;
  wire       [0:0]    in_x7_1;
  wire       [0:0]    in_x7_2;
  wire       [0:0]    in_x7_3;
  wire       [0:0]    out_y0_0;
  wire       [0:0]    out_y0_1;
  wire       [0:0]    out_y0_2;
  wire       [0:0]    out_y0_3;
  wire       [0:0]    out_y1_0;
  wire       [0:0]    out_y1_1;
  wire       [0:0]    out_y1_2;
  wire       [0:0]    out_y1_3;
  wire       [0:0]    out_y2_0;
  wire       [0:0]    out_y2_1;
  wire       [0:0]    out_y2_2;
  wire       [0:0]    out_y2_3;
  wire       [0:0]    out_y3_0;
  wire       [0:0]    out_y3_1;
  wire       [0:0]    out_y3_2;
  wire       [0:0]    out_y3_3;
  wire       [0:0]    out_y4_0;
  wire       [0:0]    out_y4_1;
  wire       [0:0]    out_y4_2;
  wire       [0:0]    out_y4_3;
  wire       [0:0]    out_y5_0;
  wire       [0:0]    out_y5_1;
  wire       [0:0]    out_y5_2;
  wire       [0:0]    out_y5_3;
  wire       [0:0]    out_y6_0;
  wire       [0:0]    out_y6_1;
  wire       [0:0]    out_y6_2;
  wire       [0:0]    out_y6_3;
  wire       [0:0]    out_y7_0;
  wire       [0:0]    out_y7_1;
  wire       [0:0]    out_y7_2;
  wire       [0:0]    out_y7_3;
  reg        [0:0]    x7_0;
  reg        [0:0]    x7_1;
  reg        [0:0]    x7_2;
  reg        [0:0]    x7_3;
  reg        [0:0]    t1_0;
  reg        [0:0]    t1_1;
  reg        [0:0]    t1_2;
  reg        [0:0]    t1_3;
  reg        [0:0]    t2_0;
  reg        [0:0]    t2_1;
  reg        [0:0]    t2_2;
  reg        [0:0]    t2_3;
  reg        [0:0]    t3_0;
  reg        [0:0]    t3_1;
  reg        [0:0]    t3_2;
  reg        [0:0]    t3_3;
  reg        [0:0]    t4_0;
  reg        [0:0]    t4_1;
  reg        [0:0]    t4_2;
  reg        [0:0]    t4_3;
  reg        [0:0]    t6_0;
  reg        [0:0]    t6_1;
  reg        [0:0]    t6_2;
  reg        [0:0]    t6_3;
  reg        [0:0]    t7_0;
  reg        [0:0]    t7_1;
  reg        [0:0]    t7_2;
  reg        [0:0]    t7_3;
  reg        [0:0]    t8_0;
  reg        [0:0]    t8_1;
  reg        [0:0]    t8_2;
  reg        [0:0]    t8_3;
  reg        [0:0]    t9_0;
  reg        [0:0]    t9_1;
  reg        [0:0]    t9_2;
  reg        [0:0]    t9_3;
  reg        [0:0]    t10_0;
  reg        [0:0]    t10_1;
  reg        [0:0]    t10_2;
  reg        [0:0]    t10_3;
  reg        [0:0]    t13_0;
  reg        [0:0]    t13_1;
  reg        [0:0]    t13_2;
  reg        [0:0]    t13_3;
  reg        [0:0]    t14_0;
  reg        [0:0]    t14_1;
  reg        [0:0]    t14_2;
  reg        [0:0]    t14_3;
  reg        [0:0]    t15_0;
  reg        [0:0]    t15_1;
  reg        [0:0]    t15_2;
  reg        [0:0]    t15_3;
  reg        [0:0]    t16_0;
  reg        [0:0]    t16_1;
  reg        [0:0]    t16_2;
  reg        [0:0]    t16_3;
  reg        [0:0]    t17_0;
  reg        [0:0]    t17_1;
  reg        [0:0]    t17_2;
  reg        [0:0]    t17_3;
  reg        [0:0]    t19_0;
  reg        [0:0]    t19_1;
  reg        [0:0]    t19_2;
  reg        [0:0]    t19_3;
  reg        [0:0]    t20_0;
  reg        [0:0]    t20_1;
  reg        [0:0]    t20_2;
  reg        [0:0]    t20_3;
  reg        [0:0]    t22_0;
  reg        [0:0]    t22_1;
  reg        [0:0]    t22_2;
  reg        [0:0]    t22_3;
  reg        [0:0]    t23_0;
  reg        [0:0]    t23_1;
  reg        [0:0]    t23_2;
  reg        [0:0]    t23_3;
  reg        [0:0]    t24_0;
  reg        [0:0]    t24_1;
  reg        [0:0]    t24_2;
  reg        [0:0]    t24_3;
  reg        [0:0]    t25_0;
  reg        [0:0]    t25_1;
  reg        [0:0]    t25_2;
  reg        [0:0]    t25_3;
  reg        [0:0]    t26_0;
  reg        [0:0]    t26_1;
  reg        [0:0]    t26_2;
  reg        [0:0]    t26_3;
  reg        [0:0]    t27_0;
  reg        [0:0]    t27_1;
  reg        [0:0]    t27_2;
  reg        [0:0]    t27_3;
  reg        [0:0]    x7_1_0;
  reg        [0:0]    x7_1_1;
  reg        [0:0]    x7_1_2;
  reg        [0:0]    x7_1_3;
  reg        [0:0]    t1_1_0;
  reg        [0:0]    t1_1_1;
  reg        [0:0]    t1_1_2;
  reg        [0:0]    t1_1_3;
  reg        [0:0]    t2_1_0;
  reg        [0:0]    t2_1_1;
  reg        [0:0]    t2_1_2;
  reg        [0:0]    t2_1_3;
  reg        [0:0]    t3_1_0;
  reg        [0:0]    t3_1_1;
  reg        [0:0]    t3_1_2;
  reg        [0:0]    t3_1_3;
  reg        [0:0]    t4_1_0;
  reg        [0:0]    t4_1_1;
  reg        [0:0]    t4_1_2;
  reg        [0:0]    t4_1_3;
  reg        [0:0]    t6_1_0;
  reg        [0:0]    t6_1_1;
  reg        [0:0]    t6_1_2;
  reg        [0:0]    t6_1_3;
  reg        [0:0]    t8_1_0;
  reg        [0:0]    t8_1_1;
  reg        [0:0]    t8_1_2;
  reg        [0:0]    t8_1_3;
  reg        [0:0]    t9_1_0;
  reg        [0:0]    t9_1_1;
  reg        [0:0]    t9_1_2;
  reg        [0:0]    t9_1_3;
  reg        [0:0]    t10_1_0;
  reg        [0:0]    t10_1_1;
  reg        [0:0]    t10_1_2;
  reg        [0:0]    t10_1_3;
  reg        [0:0]    t13_1_0;
  reg        [0:0]    t13_1_1;
  reg        [0:0]    t13_1_2;
  reg        [0:0]    t13_1_3;
  reg        [0:0]    t15_1_0;
  reg        [0:0]    t15_1_1;
  reg        [0:0]    t15_1_2;
  reg        [0:0]    t15_1_3;
  reg        [0:0]    t16_1_0;
  reg        [0:0]    t16_1_1;
  reg        [0:0]    t16_1_2;
  reg        [0:0]    t16_1_3;
  reg        [0:0]    t17_1_0;
  reg        [0:0]    t17_1_1;
  reg        [0:0]    t17_1_2;
  reg        [0:0]    t17_1_3;
  reg        [0:0]    t19_1_0;
  reg        [0:0]    t19_1_1;
  reg        [0:0]    t19_1_2;
  reg        [0:0]    t19_1_3;
  reg        [0:0]    t20_1_0;
  reg        [0:0]    t20_1_1;
  reg        [0:0]    t20_1_2;
  reg        [0:0]    t20_1_3;
  reg        [0:0]    t22_1_0;
  reg        [0:0]    t22_1_1;
  reg        [0:0]    t22_1_2;
  reg        [0:0]    t22_1_3;
  reg        [0:0]    t23_1_0;
  reg        [0:0]    t23_1_1;
  reg        [0:0]    t23_1_2;
  reg        [0:0]    t23_1_3;
  reg        [0:0]    t27_1_0;
  reg        [0:0]    t27_1_1;
  reg        [0:0]    t27_1_2;
  reg        [0:0]    t27_1_3;
  reg        [0:0]    m21_0;
  reg        [0:0]    m21_1;
  reg        [0:0]    m21_2;
  reg        [0:0]    m21_3;
  reg        [0:0]    m23_0;
  reg        [0:0]    m23_1;
  reg        [0:0]    m23_2;
  reg        [0:0]    m23_3;
  reg        [0:0]    m24_0;
  reg        [0:0]    m24_1;
  reg        [0:0]    m24_2;
  reg        [0:0]    m24_3;
  reg        [0:0]    m27_0;
  reg        [0:0]    m27_1;
  reg        [0:0]    m27_2;
  reg        [0:0]    m27_3;
  reg        [0:0]    x7_2_0;
  reg        [0:0]    x7_2_1;
  reg        [0:0]    x7_2_2;
  reg        [0:0]    x7_2_3;
  reg        [0:0]    t1_2_0;
  reg        [0:0]    t1_2_1;
  reg        [0:0]    t1_2_2;
  reg        [0:0]    t1_2_3;
  reg        [0:0]    t2_2_0;
  reg        [0:0]    t2_2_1;
  reg        [0:0]    t2_2_2;
  reg        [0:0]    t2_2_3;
  reg        [0:0]    t3_2_0;
  reg        [0:0]    t3_2_1;
  reg        [0:0]    t3_2_2;
  reg        [0:0]    t3_2_3;
  reg        [0:0]    t4_2_0;
  reg        [0:0]    t4_2_1;
  reg        [0:0]    t4_2_2;
  reg        [0:0]    t4_2_3;
  reg        [0:0]    t6_2_0;
  reg        [0:0]    t6_2_1;
  reg        [0:0]    t6_2_2;
  reg        [0:0]    t6_2_3;
  reg        [0:0]    t8_2_0;
  reg        [0:0]    t8_2_1;
  reg        [0:0]    t8_2_2;
  reg        [0:0]    t8_2_3;
  reg        [0:0]    t9_2_0;
  reg        [0:0]    t9_2_1;
  reg        [0:0]    t9_2_2;
  reg        [0:0]    t9_2_3;
  reg        [0:0]    t10_2_0;
  reg        [0:0]    t10_2_1;
  reg        [0:0]    t10_2_2;
  reg        [0:0]    t10_2_3;
  reg        [0:0]    t13_2_0;
  reg        [0:0]    t13_2_1;
  reg        [0:0]    t13_2_2;
  reg        [0:0]    t13_2_3;
  reg        [0:0]    t15_2_0;
  reg        [0:0]    t15_2_1;
  reg        [0:0]    t15_2_2;
  reg        [0:0]    t15_2_3;
  reg        [0:0]    t16_2_0;
  reg        [0:0]    t16_2_1;
  reg        [0:0]    t16_2_2;
  reg        [0:0]    t16_2_3;
  reg        [0:0]    t17_2_0;
  reg        [0:0]    t17_2_1;
  reg        [0:0]    t17_2_2;
  reg        [0:0]    t17_2_3;
  reg        [0:0]    t19_2_0;
  reg        [0:0]    t19_2_1;
  reg        [0:0]    t19_2_2;
  reg        [0:0]    t19_2_3;
  reg        [0:0]    t20_2_0;
  reg        [0:0]    t20_2_1;
  reg        [0:0]    t20_2_2;
  reg        [0:0]    t20_2_3;
  reg        [0:0]    t22_2_0;
  reg        [0:0]    t22_2_1;
  reg        [0:0]    t22_2_2;
  reg        [0:0]    t22_2_3;
  reg        [0:0]    t23_2_0;
  reg        [0:0]    t23_2_1;
  reg        [0:0]    t23_2_2;
  reg        [0:0]    t23_2_3;
  reg        [0:0]    t27_2_0;
  reg        [0:0]    t27_2_1;
  reg        [0:0]    t27_2_2;
  reg        [0:0]    t27_2_3;
  reg        [0:0]    m21_1_0;
  reg        [0:0]    m21_1_1;
  reg        [0:0]    m21_1_2;
  reg        [0:0]    m21_1_3;
  reg        [0:0]    m23_1_0;
  reg        [0:0]    m23_1_1;
  reg        [0:0]    m23_1_2;
  reg        [0:0]    m23_1_3;
  reg        [0:0]    m33_0;
  reg        [0:0]    m33_1;
  reg        [0:0]    m33_2;
  reg        [0:0]    m33_3;
  reg        [0:0]    m36_0;
  reg        [0:0]    m36_1;
  reg        [0:0]    m36_2;
  reg        [0:0]    m36_3;

  Addition_TI t1_xor (
    .port_x0_0 (in_x0_0        ), //i
    .port_x0_1 (in_x0_1        ), //i
    .port_x0_2 (in_x0_2        ), //i
    .port_x0_3 (in_x0_3        ), //i
    .port_x1_0 (in_x3_0        ), //i
    .port_x1_1 (in_x3_1        ), //i
    .port_x1_2 (in_x3_2        ), //i
    .port_x1_3 (in_x3_3        ), //i
    .port_y_0  (t1_xor_port_y_0), //o
    .port_y_1  (t1_xor_port_y_1), //o
    .port_y_2  (t1_xor_port_y_2), //o
    .port_y_3  (t1_xor_port_y_3)  //o
  );
  Addition_TI t2_xor (
    .port_x0_0 (in_x0_0        ), //i
    .port_x0_1 (in_x0_1        ), //i
    .port_x0_2 (in_x0_2        ), //i
    .port_x0_3 (in_x0_3        ), //i
    .port_x1_0 (in_x5_0        ), //i
    .port_x1_1 (in_x5_1        ), //i
    .port_x1_2 (in_x5_2        ), //i
    .port_x1_3 (in_x5_3        ), //i
    .port_y_0  (t2_xor_port_y_0), //o
    .port_y_1  (t2_xor_port_y_1), //o
    .port_y_2  (t2_xor_port_y_2), //o
    .port_y_3  (t2_xor_port_y_3)  //o
  );
  Addition_TI t3_xor (
    .port_x0_0 (in_x0_0        ), //i
    .port_x0_1 (in_x0_1        ), //i
    .port_x0_2 (in_x0_2        ), //i
    .port_x0_3 (in_x0_3        ), //i
    .port_x1_0 (in_x6_0        ), //i
    .port_x1_1 (in_x6_1        ), //i
    .port_x1_2 (in_x6_2        ), //i
    .port_x1_3 (in_x6_3        ), //i
    .port_y_0  (t3_xor_port_y_0), //o
    .port_y_1  (t3_xor_port_y_1), //o
    .port_y_2  (t3_xor_port_y_2), //o
    .port_y_3  (t3_xor_port_y_3)  //o
  );
  Addition_TI t4_xor (
    .port_x0_0 (in_x3_0        ), //i
    .port_x0_1 (in_x3_1        ), //i
    .port_x0_2 (in_x3_2        ), //i
    .port_x0_3 (in_x3_3        ), //i
    .port_x1_0 (in_x5_0        ), //i
    .port_x1_1 (in_x5_1        ), //i
    .port_x1_2 (in_x5_2        ), //i
    .port_x1_3 (in_x5_3        ), //i
    .port_y_0  (t4_xor_port_y_0), //o
    .port_y_1  (t4_xor_port_y_1), //o
    .port_y_2  (t4_xor_port_y_2), //o
    .port_y_3  (t4_xor_port_y_3)  //o
  );
  Addition_TI t5_xor (
    .port_x0_0 (in_x4_0        ), //i
    .port_x0_1 (in_x4_1        ), //i
    .port_x0_2 (in_x4_2        ), //i
    .port_x0_3 (in_x4_3        ), //i
    .port_x1_0 (in_x6_0        ), //i
    .port_x1_1 (in_x6_1        ), //i
    .port_x1_2 (in_x6_2        ), //i
    .port_x1_3 (in_x6_3        ), //i
    .port_y_0  (t5_xor_port_y_0), //o
    .port_y_1  (t5_xor_port_y_1), //o
    .port_y_2  (t5_xor_port_y_2), //o
    .port_y_3  (t5_xor_port_y_3)  //o
  );
  Addition_TI t6_xor (
    .port_x0_0 (t1_xor_port_y_0), //i
    .port_x0_1 (t1_xor_port_y_1), //i
    .port_x0_2 (t1_xor_port_y_2), //i
    .port_x0_3 (t1_xor_port_y_3), //i
    .port_x1_0 (t5_xor_port_y_0), //i
    .port_x1_1 (t5_xor_port_y_1), //i
    .port_x1_2 (t5_xor_port_y_2), //i
    .port_x1_3 (t5_xor_port_y_3), //i
    .port_y_0  (t6_xor_port_y_0), //o
    .port_y_1  (t6_xor_port_y_1), //o
    .port_y_2  (t6_xor_port_y_2), //o
    .port_y_3  (t6_xor_port_y_3)  //o
  );
  Addition_TI t7_xor (
    .port_x0_0 (in_x1_0        ), //i
    .port_x0_1 (in_x1_1        ), //i
    .port_x0_2 (in_x1_2        ), //i
    .port_x0_3 (in_x1_3        ), //i
    .port_x1_0 (in_x2_0        ), //i
    .port_x1_1 (in_x2_1        ), //i
    .port_x1_2 (in_x2_2        ), //i
    .port_x1_3 (in_x2_3        ), //i
    .port_y_0  (t7_xor_port_y_0), //o
    .port_y_1  (t7_xor_port_y_1), //o
    .port_y_2  (t7_xor_port_y_2), //o
    .port_y_3  (t7_xor_port_y_3)  //o
  );
  Addition_TI t8_xor (
    .port_x0_0 (in_x7_0        ), //i
    .port_x0_1 (in_x7_1        ), //i
    .port_x0_2 (in_x7_2        ), //i
    .port_x0_3 (in_x7_3        ), //i
    .port_x1_0 (t6_xor_port_y_0), //i
    .port_x1_1 (t6_xor_port_y_1), //i
    .port_x1_2 (t6_xor_port_y_2), //i
    .port_x1_3 (t6_xor_port_y_3), //i
    .port_y_0  (t8_xor_port_y_0), //o
    .port_y_1  (t8_xor_port_y_1), //o
    .port_y_2  (t8_xor_port_y_2), //o
    .port_y_3  (t8_xor_port_y_3)  //o
  );
  Addition_TI t9_xor (
    .port_x0_0 (in_x7_0        ), //i
    .port_x0_1 (in_x7_1        ), //i
    .port_x0_2 (in_x7_2        ), //i
    .port_x0_3 (in_x7_3        ), //i
    .port_x1_0 (t7_xor_port_y_0), //i
    .port_x1_1 (t7_xor_port_y_1), //i
    .port_x1_2 (t7_xor_port_y_2), //i
    .port_x1_3 (t7_xor_port_y_3), //i
    .port_y_0  (t9_xor_port_y_0), //o
    .port_y_1  (t9_xor_port_y_1), //o
    .port_y_2  (t9_xor_port_y_2), //o
    .port_y_3  (t9_xor_port_y_3)  //o
  );
  Addition_TI t10_xor (
    .port_x0_0 (t6_xor_port_y_0 ), //i
    .port_x0_1 (t6_xor_port_y_1 ), //i
    .port_x0_2 (t6_xor_port_y_2 ), //i
    .port_x0_3 (t6_xor_port_y_3 ), //i
    .port_x1_0 (t7_xor_port_y_0 ), //i
    .port_x1_1 (t7_xor_port_y_1 ), //i
    .port_x1_2 (t7_xor_port_y_2 ), //i
    .port_x1_3 (t7_xor_port_y_3 ), //i
    .port_y_0  (t10_xor_port_y_0), //o
    .port_y_1  (t10_xor_port_y_1), //o
    .port_y_2  (t10_xor_port_y_2), //o
    .port_y_3  (t10_xor_port_y_3)  //o
  );
  Addition_TI t11_xor (
    .port_x0_0 (in_x1_0         ), //i
    .port_x0_1 (in_x1_1         ), //i
    .port_x0_2 (in_x1_2         ), //i
    .port_x0_3 (in_x1_3         ), //i
    .port_x1_0 (in_x5_0         ), //i
    .port_x1_1 (in_x5_1         ), //i
    .port_x1_2 (in_x5_2         ), //i
    .port_x1_3 (in_x5_3         ), //i
    .port_y_0  (t11_xor_port_y_0), //o
    .port_y_1  (t11_xor_port_y_1), //o
    .port_y_2  (t11_xor_port_y_2), //o
    .port_y_3  (t11_xor_port_y_3)  //o
  );
  Addition_TI t12_xor (
    .port_x0_0 (in_x2_0         ), //i
    .port_x0_1 (in_x2_1         ), //i
    .port_x0_2 (in_x2_2         ), //i
    .port_x0_3 (in_x2_3         ), //i
    .port_x1_0 (in_x5_0         ), //i
    .port_x1_1 (in_x5_1         ), //i
    .port_x1_2 (in_x5_2         ), //i
    .port_x1_3 (in_x5_3         ), //i
    .port_y_0  (t12_xor_port_y_0), //o
    .port_y_1  (t12_xor_port_y_1), //o
    .port_y_2  (t12_xor_port_y_2), //o
    .port_y_3  (t12_xor_port_y_3)  //o
  );
  Addition_TI t13_xor (
    .port_x0_0 (t3_xor_port_y_0 ), //i
    .port_x0_1 (t3_xor_port_y_1 ), //i
    .port_x0_2 (t3_xor_port_y_2 ), //i
    .port_x0_3 (t3_xor_port_y_3 ), //i
    .port_x1_0 (t4_xor_port_y_0 ), //i
    .port_x1_1 (t4_xor_port_y_1 ), //i
    .port_x1_2 (t4_xor_port_y_2 ), //i
    .port_x1_3 (t4_xor_port_y_3 ), //i
    .port_y_0  (t13_xor_port_y_0), //o
    .port_y_1  (t13_xor_port_y_1), //o
    .port_y_2  (t13_xor_port_y_2), //o
    .port_y_3  (t13_xor_port_y_3)  //o
  );
  Addition_TI t14_xor (
    .port_x0_0 (t6_xor_port_y_0 ), //i
    .port_x0_1 (t6_xor_port_y_1 ), //i
    .port_x0_2 (t6_xor_port_y_2 ), //i
    .port_x0_3 (t6_xor_port_y_3 ), //i
    .port_x1_0 (t11_xor_port_y_0), //i
    .port_x1_1 (t11_xor_port_y_1), //i
    .port_x1_2 (t11_xor_port_y_2), //i
    .port_x1_3 (t11_xor_port_y_3), //i
    .port_y_0  (t14_xor_port_y_0), //o
    .port_y_1  (t14_xor_port_y_1), //o
    .port_y_2  (t14_xor_port_y_2), //o
    .port_y_3  (t14_xor_port_y_3)  //o
  );
  Addition_TI t15_xor (
    .port_x0_0 (t5_xor_port_y_0 ), //i
    .port_x0_1 (t5_xor_port_y_1 ), //i
    .port_x0_2 (t5_xor_port_y_2 ), //i
    .port_x0_3 (t5_xor_port_y_3 ), //i
    .port_x1_0 (t11_xor_port_y_0), //i
    .port_x1_1 (t11_xor_port_y_1), //i
    .port_x1_2 (t11_xor_port_y_2), //i
    .port_x1_3 (t11_xor_port_y_3), //i
    .port_y_0  (t15_xor_port_y_0), //o
    .port_y_1  (t15_xor_port_y_1), //o
    .port_y_2  (t15_xor_port_y_2), //o
    .port_y_3  (t15_xor_port_y_3)  //o
  );
  Addition_TI t16_xor (
    .port_x0_0 (t5_xor_port_y_0 ), //i
    .port_x0_1 (t5_xor_port_y_1 ), //i
    .port_x0_2 (t5_xor_port_y_2 ), //i
    .port_x0_3 (t5_xor_port_y_3 ), //i
    .port_x1_0 (t12_xor_port_y_0), //i
    .port_x1_1 (t12_xor_port_y_1), //i
    .port_x1_2 (t12_xor_port_y_2), //i
    .port_x1_3 (t12_xor_port_y_3), //i
    .port_y_0  (t16_xor_port_y_0), //o
    .port_y_1  (t16_xor_port_y_1), //o
    .port_y_2  (t16_xor_port_y_2), //o
    .port_y_3  (t16_xor_port_y_3)  //o
  );
  Addition_TI t17_xor (
    .port_x0_0 (t9_xor_port_y_0 ), //i
    .port_x0_1 (t9_xor_port_y_1 ), //i
    .port_x0_2 (t9_xor_port_y_2 ), //i
    .port_x0_3 (t9_xor_port_y_3 ), //i
    .port_x1_0 (t16_xor_port_y_0), //i
    .port_x1_1 (t16_xor_port_y_1), //i
    .port_x1_2 (t16_xor_port_y_2), //i
    .port_x1_3 (t16_xor_port_y_3), //i
    .port_y_0  (t17_xor_port_y_0), //o
    .port_y_1  (t17_xor_port_y_1), //o
    .port_y_2  (t17_xor_port_y_2), //o
    .port_y_3  (t17_xor_port_y_3)  //o
  );
  Addition_TI t18_xor (
    .port_x0_0 (in_x3_0         ), //i
    .port_x0_1 (in_x3_1         ), //i
    .port_x0_2 (in_x3_2         ), //i
    .port_x0_3 (in_x3_3         ), //i
    .port_x1_0 (in_x7_0         ), //i
    .port_x1_1 (in_x7_1         ), //i
    .port_x1_2 (in_x7_2         ), //i
    .port_x1_3 (in_x7_3         ), //i
    .port_y_0  (t18_xor_port_y_0), //o
    .port_y_1  (t18_xor_port_y_1), //o
    .port_y_2  (t18_xor_port_y_2), //o
    .port_y_3  (t18_xor_port_y_3)  //o
  );
  Addition_TI t19_xor (
    .port_x0_0 (t7_xor_port_y_0 ), //i
    .port_x0_1 (t7_xor_port_y_1 ), //i
    .port_x0_2 (t7_xor_port_y_2 ), //i
    .port_x0_3 (t7_xor_port_y_3 ), //i
    .port_x1_0 (t18_xor_port_y_0), //i
    .port_x1_1 (t18_xor_port_y_1), //i
    .port_x1_2 (t18_xor_port_y_2), //i
    .port_x1_3 (t18_xor_port_y_3), //i
    .port_y_0  (t19_xor_port_y_0), //o
    .port_y_1  (t19_xor_port_y_1), //o
    .port_y_2  (t19_xor_port_y_2), //o
    .port_y_3  (t19_xor_port_y_3)  //o
  );
  Addition_TI t20_xor (
    .port_x0_0 (t1_xor_port_y_0 ), //i
    .port_x0_1 (t1_xor_port_y_1 ), //i
    .port_x0_2 (t1_xor_port_y_2 ), //i
    .port_x0_3 (t1_xor_port_y_3 ), //i
    .port_x1_0 (t19_xor_port_y_0), //i
    .port_x1_1 (t19_xor_port_y_1), //i
    .port_x1_2 (t19_xor_port_y_2), //i
    .port_x1_3 (t19_xor_port_y_3), //i
    .port_y_0  (t20_xor_port_y_0), //o
    .port_y_1  (t20_xor_port_y_1), //o
    .port_y_2  (t20_xor_port_y_2), //o
    .port_y_3  (t20_xor_port_y_3)  //o
  );
  Addition_TI t21_xor (
    .port_x0_0 (in_x6_0         ), //i
    .port_x0_1 (in_x6_1         ), //i
    .port_x0_2 (in_x6_2         ), //i
    .port_x0_3 (in_x6_3         ), //i
    .port_x1_0 (in_x7_0         ), //i
    .port_x1_1 (in_x7_1         ), //i
    .port_x1_2 (in_x7_2         ), //i
    .port_x1_3 (in_x7_3         ), //i
    .port_y_0  (t21_xor_port_y_0), //o
    .port_y_1  (t21_xor_port_y_1), //o
    .port_y_2  (t21_xor_port_y_2), //o
    .port_y_3  (t21_xor_port_y_3)  //o
  );
  Addition_TI t22_xor (
    .port_x0_0 (t7_xor_port_y_0 ), //i
    .port_x0_1 (t7_xor_port_y_1 ), //i
    .port_x0_2 (t7_xor_port_y_2 ), //i
    .port_x0_3 (t7_xor_port_y_3 ), //i
    .port_x1_0 (t21_xor_port_y_0), //i
    .port_x1_1 (t21_xor_port_y_1), //i
    .port_x1_2 (t21_xor_port_y_2), //i
    .port_x1_3 (t21_xor_port_y_3), //i
    .port_y_0  (t22_xor_port_y_0), //o
    .port_y_1  (t22_xor_port_y_1), //o
    .port_y_2  (t22_xor_port_y_2), //o
    .port_y_3  (t22_xor_port_y_3)  //o
  );
  Addition_TI t23_xor (
    .port_x0_0 (t2_xor_port_y_0 ), //i
    .port_x0_1 (t2_xor_port_y_1 ), //i
    .port_x0_2 (t2_xor_port_y_2 ), //i
    .port_x0_3 (t2_xor_port_y_3 ), //i
    .port_x1_0 (t22_xor_port_y_0), //i
    .port_x1_1 (t22_xor_port_y_1), //i
    .port_x1_2 (t22_xor_port_y_2), //i
    .port_x1_3 (t22_xor_port_y_3), //i
    .port_y_0  (t23_xor_port_y_0), //o
    .port_y_1  (t23_xor_port_y_1), //o
    .port_y_2  (t23_xor_port_y_2), //o
    .port_y_3  (t23_xor_port_y_3)  //o
  );
  Addition_TI t24_xor (
    .port_x0_0 (t2_xor_port_y_0 ), //i
    .port_x0_1 (t2_xor_port_y_1 ), //i
    .port_x0_2 (t2_xor_port_y_2 ), //i
    .port_x0_3 (t2_xor_port_y_3 ), //i
    .port_x1_0 (t10_xor_port_y_0), //i
    .port_x1_1 (t10_xor_port_y_1), //i
    .port_x1_2 (t10_xor_port_y_2), //i
    .port_x1_3 (t10_xor_port_y_3), //i
    .port_y_0  (t24_xor_port_y_0), //o
    .port_y_1  (t24_xor_port_y_1), //o
    .port_y_2  (t24_xor_port_y_2), //o
    .port_y_3  (t24_xor_port_y_3)  //o
  );
  Addition_TI t25_xor (
    .port_x0_0 (t20_xor_port_y_0), //i
    .port_x0_1 (t20_xor_port_y_1), //i
    .port_x0_2 (t20_xor_port_y_2), //i
    .port_x0_3 (t20_xor_port_y_3), //i
    .port_x1_0 (t17_xor_port_y_0), //i
    .port_x1_1 (t17_xor_port_y_1), //i
    .port_x1_2 (t17_xor_port_y_2), //i
    .port_x1_3 (t17_xor_port_y_3), //i
    .port_y_0  (t25_xor_port_y_0), //o
    .port_y_1  (t25_xor_port_y_1), //o
    .port_y_2  (t25_xor_port_y_2), //o
    .port_y_3  (t25_xor_port_y_3)  //o
  );
  Addition_TI t26_xor (
    .port_x0_0 (t3_xor_port_y_0 ), //i
    .port_x0_1 (t3_xor_port_y_1 ), //i
    .port_x0_2 (t3_xor_port_y_2 ), //i
    .port_x0_3 (t3_xor_port_y_3 ), //i
    .port_x1_0 (t16_xor_port_y_0), //i
    .port_x1_1 (t16_xor_port_y_1), //i
    .port_x1_2 (t16_xor_port_y_2), //i
    .port_x1_3 (t16_xor_port_y_3), //i
    .port_y_0  (t26_xor_port_y_0), //o
    .port_y_1  (t26_xor_port_y_1), //o
    .port_y_2  (t26_xor_port_y_2), //o
    .port_y_3  (t26_xor_port_y_3)  //o
  );
  Addition_TI t27_xor (
    .port_x0_0 (t1_xor_port_y_0 ), //i
    .port_x0_1 (t1_xor_port_y_1 ), //i
    .port_x0_2 (t1_xor_port_y_2 ), //i
    .port_x0_3 (t1_xor_port_y_3 ), //i
    .port_x1_0 (t12_xor_port_y_0), //i
    .port_x1_1 (t12_xor_port_y_1), //i
    .port_x1_2 (t12_xor_port_y_2), //i
    .port_x1_3 (t12_xor_port_y_3), //i
    .port_y_0  (t27_xor_port_y_0), //o
    .port_y_1  (t27_xor_port_y_1), //o
    .port_y_2  (t27_xor_port_y_2), //o
    .port_y_3  (t27_xor_port_y_3)  //o
  );
  Multiplication_TI m1 (
    .port_x0_0 (t13_xor_port_y_0), //i
    .port_x0_1 (t13_xor_port_y_1), //i
    .port_x0_2 (t13_xor_port_y_2), //i
    .port_x0_3 (t13_xor_port_y_3), //i
    .port_x1_0 (t6_xor_port_y_0 ), //i
    .port_x1_1 (t6_xor_port_y_1 ), //i
    .port_x1_2 (t6_xor_port_y_2 ), //i
    .port_x1_3 (t6_xor_port_y_3 ), //i
    .port_y_0  (m1_port_y_0     ), //o
    .port_y_1  (m1_port_y_1     ), //o
    .port_y_2  (m1_port_y_2     ), //o
    .port_y_3  (m1_port_y_3     ), //o
    .clk       (clk             ), //i
    .reset     (reset           )  //i
  );
  Multiplication_TI m2 (
    .port_x0_0 (t23_xor_port_y_0), //i
    .port_x0_1 (t23_xor_port_y_1), //i
    .port_x0_2 (t23_xor_port_y_2), //i
    .port_x0_3 (t23_xor_port_y_3), //i
    .port_x1_0 (t8_xor_port_y_0 ), //i
    .port_x1_1 (t8_xor_port_y_1 ), //i
    .port_x1_2 (t8_xor_port_y_2 ), //i
    .port_x1_3 (t8_xor_port_y_3 ), //i
    .port_y_0  (m2_port_y_0     ), //o
    .port_y_1  (m2_port_y_1     ), //o
    .port_y_2  (m2_port_y_2     ), //o
    .port_y_3  (m2_port_y_3     ), //o
    .clk       (clk             ), //i
    .reset     (reset           )  //i
  );
  Multiplication_TI m4 (
    .port_x0_0 (t19_xor_port_y_0), //i
    .port_x0_1 (t19_xor_port_y_1), //i
    .port_x0_2 (t19_xor_port_y_2), //i
    .port_x0_3 (t19_xor_port_y_3), //i
    .port_x1_0 (in_x7_0         ), //i
    .port_x1_1 (in_x7_1         ), //i
    .port_x1_2 (in_x7_2         ), //i
    .port_x1_3 (in_x7_3         ), //i
    .port_y_0  (m4_port_y_0     ), //o
    .port_y_1  (m4_port_y_1     ), //o
    .port_y_2  (m4_port_y_2     ), //o
    .port_y_3  (m4_port_y_3     ), //o
    .clk       (clk             ), //i
    .reset     (reset           )  //i
  );
  Multiplication_TI m6 (
    .port_x0_0 (t3_xor_port_y_0 ), //i
    .port_x0_1 (t3_xor_port_y_1 ), //i
    .port_x0_2 (t3_xor_port_y_2 ), //i
    .port_x0_3 (t3_xor_port_y_3 ), //i
    .port_x1_0 (t16_xor_port_y_0), //i
    .port_x1_1 (t16_xor_port_y_1), //i
    .port_x1_2 (t16_xor_port_y_2), //i
    .port_x1_3 (t16_xor_port_y_3), //i
    .port_y_0  (m6_port_y_0     ), //o
    .port_y_1  (m6_port_y_1     ), //o
    .port_y_2  (m6_port_y_2     ), //o
    .port_y_3  (m6_port_y_3     ), //o
    .clk       (clk             ), //i
    .reset     (reset           )  //i
  );
  Multiplication_TI m7 (
    .port_x0_0 (t22_xor_port_y_0), //i
    .port_x0_1 (t22_xor_port_y_1), //i
    .port_x0_2 (t22_xor_port_y_2), //i
    .port_x0_3 (t22_xor_port_y_3), //i
    .port_x1_0 (t9_xor_port_y_0 ), //i
    .port_x1_1 (t9_xor_port_y_1 ), //i
    .port_x1_2 (t9_xor_port_y_2 ), //i
    .port_x1_3 (t9_xor_port_y_3 ), //i
    .port_y_0  (m7_port_y_0     ), //o
    .port_y_1  (m7_port_y_1     ), //o
    .port_y_2  (m7_port_y_2     ), //o
    .port_y_3  (m7_port_y_3     ), //o
    .clk       (clk             ), //i
    .reset     (reset           )  //i
  );
  Multiplication_TI m9 (
    .port_x0_0 (t20_xor_port_y_0), //i
    .port_x0_1 (t20_xor_port_y_1), //i
    .port_x0_2 (t20_xor_port_y_2), //i
    .port_x0_3 (t20_xor_port_y_3), //i
    .port_x1_0 (t17_xor_port_y_0), //i
    .port_x1_1 (t17_xor_port_y_1), //i
    .port_x1_2 (t17_xor_port_y_2), //i
    .port_x1_3 (t17_xor_port_y_3), //i
    .port_y_0  (m9_port_y_0     ), //o
    .port_y_1  (m9_port_y_1     ), //o
    .port_y_2  (m9_port_y_2     ), //o
    .port_y_3  (m9_port_y_3     ), //o
    .clk       (clk             ), //i
    .reset     (reset           )  //i
  );
  Multiplication_TI m11 (
    .port_x0_0 (t1_xor_port_y_0 ), //i
    .port_x0_1 (t1_xor_port_y_1 ), //i
    .port_x0_2 (t1_xor_port_y_2 ), //i
    .port_x0_3 (t1_xor_port_y_3 ), //i
    .port_x1_0 (t15_xor_port_y_0), //i
    .port_x1_1 (t15_xor_port_y_1), //i
    .port_x1_2 (t15_xor_port_y_2), //i
    .port_x1_3 (t15_xor_port_y_3), //i
    .port_y_0  (m11_port_y_0    ), //o
    .port_y_1  (m11_port_y_1    ), //o
    .port_y_2  (m11_port_y_2    ), //o
    .port_y_3  (m11_port_y_3    ), //o
    .clk       (clk             ), //i
    .reset     (reset           )  //i
  );
  Multiplication_TI m12 (
    .port_x0_0 (t4_xor_port_y_0 ), //i
    .port_x0_1 (t4_xor_port_y_1 ), //i
    .port_x0_2 (t4_xor_port_y_2 ), //i
    .port_x0_3 (t4_xor_port_y_3 ), //i
    .port_x1_0 (t27_xor_port_y_0), //i
    .port_x1_1 (t27_xor_port_y_1), //i
    .port_x1_2 (t27_xor_port_y_2), //i
    .port_x1_3 (t27_xor_port_y_3), //i
    .port_y_0  (m12_port_y_0    ), //o
    .port_y_1  (m12_port_y_1    ), //o
    .port_y_2  (m12_port_y_2    ), //o
    .port_y_3  (m12_port_y_3    ), //o
    .clk       (clk             ), //i
    .reset     (reset           )  //i
  );
  Multiplication_TI m14 (
    .port_x0_0 (t2_xor_port_y_0 ), //i
    .port_x0_1 (t2_xor_port_y_1 ), //i
    .port_x0_2 (t2_xor_port_y_2 ), //i
    .port_x0_3 (t2_xor_port_y_3 ), //i
    .port_x1_0 (t10_xor_port_y_0), //i
    .port_x1_1 (t10_xor_port_y_1), //i
    .port_x1_2 (t10_xor_port_y_2), //i
    .port_x1_3 (t10_xor_port_y_3), //i
    .port_y_0  (m14_port_y_0    ), //o
    .port_y_1  (m14_port_y_1    ), //o
    .port_y_2  (m14_port_y_2    ), //o
    .port_y_3  (m14_port_y_3    ), //o
    .clk       (clk             ), //i
    .reset     (reset           )  //i
  );
  Addition_TI m3_xor (
    .port_x0_0 (t14_0          ), //i
    .port_x0_1 (t14_1          ), //i
    .port_x0_2 (t14_2          ), //i
    .port_x0_3 (t14_3          ), //i
    .port_x1_0 (m1_port_y_0    ), //i
    .port_x1_1 (m1_port_y_1    ), //i
    .port_x1_2 (m1_port_y_2    ), //i
    .port_x1_3 (m1_port_y_3    ), //i
    .port_y_0  (m3_xor_port_y_0), //o
    .port_y_1  (m3_xor_port_y_1), //o
    .port_y_2  (m3_xor_port_y_2), //o
    .port_y_3  (m3_xor_port_y_3)  //o
  );
  Addition_TI m5_xor (
    .port_x0_0 (m4_port_y_0    ), //i
    .port_x0_1 (m4_port_y_1    ), //i
    .port_x0_2 (m4_port_y_2    ), //i
    .port_x0_3 (m4_port_y_3    ), //i
    .port_x1_0 (m1_port_y_0    ), //i
    .port_x1_1 (m1_port_y_1    ), //i
    .port_x1_2 (m1_port_y_2    ), //i
    .port_x1_3 (m1_port_y_3    ), //i
    .port_y_0  (m5_xor_port_y_0), //o
    .port_y_1  (m5_xor_port_y_1), //o
    .port_y_2  (m5_xor_port_y_2), //o
    .port_y_3  (m5_xor_port_y_3)  //o
  );
  Addition_TI m8_xor (
    .port_x0_0 (t26_0          ), //i
    .port_x0_1 (t26_1          ), //i
    .port_x0_2 (t26_2          ), //i
    .port_x0_3 (t26_3          ), //i
    .port_x1_0 (m6_port_y_0    ), //i
    .port_x1_1 (m6_port_y_1    ), //i
    .port_x1_2 (m6_port_y_2    ), //i
    .port_x1_3 (m6_port_y_3    ), //i
    .port_y_0  (m8_xor_port_y_0), //o
    .port_y_1  (m8_xor_port_y_1), //o
    .port_y_2  (m8_xor_port_y_2), //o
    .port_y_3  (m8_xor_port_y_3)  //o
  );
  Addition_TI m10_xor (
    .port_x0_0 (m9_port_y_0     ), //i
    .port_x0_1 (m9_port_y_1     ), //i
    .port_x0_2 (m9_port_y_2     ), //i
    .port_x0_3 (m9_port_y_3     ), //i
    .port_x1_0 (m6_port_y_0     ), //i
    .port_x1_1 (m6_port_y_1     ), //i
    .port_x1_2 (m6_port_y_2     ), //i
    .port_x1_3 (m6_port_y_3     ), //i
    .port_y_0  (m10_xor_port_y_0), //o
    .port_y_1  (m10_xor_port_y_1), //o
    .port_y_2  (m10_xor_port_y_2), //o
    .port_y_3  (m10_xor_port_y_3)  //o
  );
  Addition_TI m13_xor (
    .port_x0_0 (m12_port_y_0    ), //i
    .port_x0_1 (m12_port_y_1    ), //i
    .port_x0_2 (m12_port_y_2    ), //i
    .port_x0_3 (m12_port_y_3    ), //i
    .port_x1_0 (m11_port_y_0    ), //i
    .port_x1_1 (m11_port_y_1    ), //i
    .port_x1_2 (m11_port_y_2    ), //i
    .port_x1_3 (m11_port_y_3    ), //i
    .port_y_0  (m13_xor_port_y_0), //o
    .port_y_1  (m13_xor_port_y_1), //o
    .port_y_2  (m13_xor_port_y_2), //o
    .port_y_3  (m13_xor_port_y_3)  //o
  );
  Addition_TI m15_xor (
    .port_x0_0 (m14_port_y_0    ), //i
    .port_x0_1 (m14_port_y_1    ), //i
    .port_x0_2 (m14_port_y_2    ), //i
    .port_x0_3 (m14_port_y_3    ), //i
    .port_x1_0 (m11_port_y_0    ), //i
    .port_x1_1 (m11_port_y_1    ), //i
    .port_x1_2 (m11_port_y_2    ), //i
    .port_x1_3 (m11_port_y_3    ), //i
    .port_y_0  (m15_xor_port_y_0), //o
    .port_y_1  (m15_xor_port_y_1), //o
    .port_y_2  (m15_xor_port_y_2), //o
    .port_y_3  (m15_xor_port_y_3)  //o
  );
  Addition_TI m16_xor (
    .port_x0_0 (m3_xor_port_y_0 ), //i
    .port_x0_1 (m3_xor_port_y_1 ), //i
    .port_x0_2 (m3_xor_port_y_2 ), //i
    .port_x0_3 (m3_xor_port_y_3 ), //i
    .port_x1_0 (m2_port_y_0     ), //i
    .port_x1_1 (m2_port_y_1     ), //i
    .port_x1_2 (m2_port_y_2     ), //i
    .port_x1_3 (m2_port_y_3     ), //i
    .port_y_0  (m16_xor_port_y_0), //o
    .port_y_1  (m16_xor_port_y_1), //o
    .port_y_2  (m16_xor_port_y_2), //o
    .port_y_3  (m16_xor_port_y_3)  //o
  );
  Addition_TI m17_xor (
    .port_x0_0 (m5_xor_port_y_0 ), //i
    .port_x0_1 (m5_xor_port_y_1 ), //i
    .port_x0_2 (m5_xor_port_y_2 ), //i
    .port_x0_3 (m5_xor_port_y_3 ), //i
    .port_x1_0 (t24_0           ), //i
    .port_x1_1 (t24_1           ), //i
    .port_x1_2 (t24_2           ), //i
    .port_x1_3 (t24_3           ), //i
    .port_y_0  (m17_xor_port_y_0), //o
    .port_y_1  (m17_xor_port_y_1), //o
    .port_y_2  (m17_xor_port_y_2), //o
    .port_y_3  (m17_xor_port_y_3)  //o
  );
  Addition_TI m18_xor (
    .port_x0_0 (m8_xor_port_y_0 ), //i
    .port_x0_1 (m8_xor_port_y_1 ), //i
    .port_x0_2 (m8_xor_port_y_2 ), //i
    .port_x0_3 (m8_xor_port_y_3 ), //i
    .port_x1_0 (m7_port_y_0     ), //i
    .port_x1_1 (m7_port_y_1     ), //i
    .port_x1_2 (m7_port_y_2     ), //i
    .port_x1_3 (m7_port_y_3     ), //i
    .port_y_0  (m18_xor_port_y_0), //o
    .port_y_1  (m18_xor_port_y_1), //o
    .port_y_2  (m18_xor_port_y_2), //o
    .port_y_3  (m18_xor_port_y_3)  //o
  );
  Addition_TI m19_xor (
    .port_x0_0 (m10_xor_port_y_0), //i
    .port_x0_1 (m10_xor_port_y_1), //i
    .port_x0_2 (m10_xor_port_y_2), //i
    .port_x0_3 (m10_xor_port_y_3), //i
    .port_x1_0 (m15_xor_port_y_0), //i
    .port_x1_1 (m15_xor_port_y_1), //i
    .port_x1_2 (m15_xor_port_y_2), //i
    .port_x1_3 (m15_xor_port_y_3), //i
    .port_y_0  (m19_xor_port_y_0), //o
    .port_y_1  (m19_xor_port_y_1), //o
    .port_y_2  (m19_xor_port_y_2), //o
    .port_y_3  (m19_xor_port_y_3)  //o
  );
  Addition_TI m20_xor (
    .port_x0_0 (m16_xor_port_y_0), //i
    .port_x0_1 (m16_xor_port_y_1), //i
    .port_x0_2 (m16_xor_port_y_2), //i
    .port_x0_3 (m16_xor_port_y_3), //i
    .port_x1_0 (m13_xor_port_y_0), //i
    .port_x1_1 (m13_xor_port_y_1), //i
    .port_x1_2 (m13_xor_port_y_2), //i
    .port_x1_3 (m13_xor_port_y_3), //i
    .port_y_0  (m20_xor_port_y_0), //o
    .port_y_1  (m20_xor_port_y_1), //o
    .port_y_2  (m20_xor_port_y_2), //o
    .port_y_3  (m20_xor_port_y_3)  //o
  );
  Addition_TI m21_xor (
    .port_x0_0 (m17_xor_port_y_0), //i
    .port_x0_1 (m17_xor_port_y_1), //i
    .port_x0_2 (m17_xor_port_y_2), //i
    .port_x0_3 (m17_xor_port_y_3), //i
    .port_x1_0 (m15_xor_port_y_0), //i
    .port_x1_1 (m15_xor_port_y_1), //i
    .port_x1_2 (m15_xor_port_y_2), //i
    .port_x1_3 (m15_xor_port_y_3), //i
    .port_y_0  (m21_xor_port_y_0), //o
    .port_y_1  (m21_xor_port_y_1), //o
    .port_y_2  (m21_xor_port_y_2), //o
    .port_y_3  (m21_xor_port_y_3)  //o
  );
  Addition_TI m22_xor (
    .port_x0_0 (m18_xor_port_y_0), //i
    .port_x0_1 (m18_xor_port_y_1), //i
    .port_x0_2 (m18_xor_port_y_2), //i
    .port_x0_3 (m18_xor_port_y_3), //i
    .port_x1_0 (m13_xor_port_y_0), //i
    .port_x1_1 (m13_xor_port_y_1), //i
    .port_x1_2 (m13_xor_port_y_2), //i
    .port_x1_3 (m13_xor_port_y_3), //i
    .port_y_0  (m22_xor_port_y_0), //o
    .port_y_1  (m22_xor_port_y_1), //o
    .port_y_2  (m22_xor_port_y_2), //o
    .port_y_3  (m22_xor_port_y_3)  //o
  );
  Addition_TI m23_xor (
    .port_x0_0 (m19_xor_port_y_0), //i
    .port_x0_1 (m19_xor_port_y_1), //i
    .port_x0_2 (m19_xor_port_y_2), //i
    .port_x0_3 (m19_xor_port_y_3), //i
    .port_x1_0 (t25_0           ), //i
    .port_x1_1 (t25_1           ), //i
    .port_x1_2 (t25_2           ), //i
    .port_x1_3 (t25_3           ), //i
    .port_y_0  (m23_xor_port_y_0), //o
    .port_y_1  (m23_xor_port_y_1), //o
    .port_y_2  (m23_xor_port_y_2), //o
    .port_y_3  (m23_xor_port_y_3)  //o
  );
  Addition_TI m24_xor (
    .port_x0_0 (m22_xor_port_y_0), //i
    .port_x0_1 (m22_xor_port_y_1), //i
    .port_x0_2 (m22_xor_port_y_2), //i
    .port_x0_3 (m22_xor_port_y_3), //i
    .port_x1_0 (m23_xor_port_y_0), //i
    .port_x1_1 (m23_xor_port_y_1), //i
    .port_x1_2 (m23_xor_port_y_2), //i
    .port_x1_3 (m23_xor_port_y_3), //i
    .port_y_0  (m24_xor_port_y_0), //o
    .port_y_1  (m24_xor_port_y_1), //o
    .port_y_2  (m24_xor_port_y_2), //o
    .port_y_3  (m24_xor_port_y_3)  //o
  );
  Multiplication_TI m25 (
    .port_x0_0 (m22_xor_port_y_0), //i
    .port_x0_1 (m22_xor_port_y_1), //i
    .port_x0_2 (m22_xor_port_y_2), //i
    .port_x0_3 (m22_xor_port_y_3), //i
    .port_x1_0 (m20_xor_port_y_0), //i
    .port_x1_1 (m20_xor_port_y_1), //i
    .port_x1_2 (m20_xor_port_y_2), //i
    .port_x1_3 (m20_xor_port_y_3), //i
    .port_y_0  (m25_port_y_0    ), //o
    .port_y_1  (m25_port_y_1    ), //o
    .port_y_2  (m25_port_y_2    ), //o
    .port_y_3  (m25_port_y_3    ), //o
    .clk       (clk             ), //i
    .reset     (reset           )  //i
  );
  Addition_TI m27_xor (
    .port_x0_0 (m20_xor_port_y_0), //i
    .port_x0_1 (m20_xor_port_y_1), //i
    .port_x0_2 (m20_xor_port_y_2), //i
    .port_x0_3 (m20_xor_port_y_3), //i
    .port_x1_0 (m21_xor_port_y_0), //i
    .port_x1_1 (m21_xor_port_y_1), //i
    .port_x1_2 (m21_xor_port_y_2), //i
    .port_x1_3 (m21_xor_port_y_3), //i
    .port_y_0  (m27_xor_port_y_0), //o
    .port_y_1  (m27_xor_port_y_1), //o
    .port_y_2  (m27_xor_port_y_2), //o
    .port_y_3  (m27_xor_port_y_3)  //o
  );
  Multiplication_TI m31 (
    .port_x0_0 (m20_xor_port_y_0), //i
    .port_x0_1 (m20_xor_port_y_1), //i
    .port_x0_2 (m20_xor_port_y_2), //i
    .port_x0_3 (m20_xor_port_y_3), //i
    .port_x1_0 (m23_xor_port_y_0), //i
    .port_x1_1 (m23_xor_port_y_1), //i
    .port_x1_2 (m23_xor_port_y_2), //i
    .port_x1_3 (m23_xor_port_y_3), //i
    .port_y_0  (m31_port_y_0    ), //o
    .port_y_1  (m31_port_y_1    ), //o
    .port_y_2  (m31_port_y_2    ), //o
    .port_y_3  (m31_port_y_3    ), //o
    .clk       (clk             ), //i
    .reset     (reset           )  //i
  );
  Multiplication_TI m34 (
    .port_x0_0 (m21_xor_port_y_0), //i
    .port_x0_1 (m21_xor_port_y_1), //i
    .port_x0_2 (m21_xor_port_y_2), //i
    .port_x0_3 (m21_xor_port_y_3), //i
    .port_x1_0 (m22_xor_port_y_0), //i
    .port_x1_1 (m22_xor_port_y_1), //i
    .port_x1_2 (m22_xor_port_y_2), //i
    .port_x1_3 (m22_xor_port_y_3), //i
    .port_y_0  (m34_port_y_0    ), //o
    .port_y_1  (m34_port_y_1    ), //o
    .port_y_2  (m34_port_y_2    ), //o
    .port_y_3  (m34_port_y_3    ), //o
    .clk       (clk             ), //i
    .reset     (reset           )  //i
  );
  Addition_TI m26_xor (
    .port_x0_0 (m21_0           ), //i
    .port_x0_1 (m21_1           ), //i
    .port_x0_2 (m21_2           ), //i
    .port_x0_3 (m21_3           ), //i
    .port_x1_0 (m25_port_y_0    ), //i
    .port_x1_1 (m25_port_y_1    ), //i
    .port_x1_2 (m25_port_y_2    ), //i
    .port_x1_3 (m25_port_y_3    ), //i
    .port_y_0  (m26_xor_port_y_0), //o
    .port_y_1  (m26_xor_port_y_1), //o
    .port_y_2  (m26_xor_port_y_2), //o
    .port_y_3  (m26_xor_port_y_3)  //o
  );
  Addition_TI m28_xor (
    .port_x0_0 (m23_0           ), //i
    .port_x0_1 (m23_1           ), //i
    .port_x0_2 (m23_2           ), //i
    .port_x0_3 (m23_3           ), //i
    .port_x1_0 (m25_port_y_0    ), //i
    .port_x1_1 (m25_port_y_1    ), //i
    .port_x1_2 (m25_port_y_2    ), //i
    .port_x1_3 (m25_port_y_3    ), //i
    .port_y_0  (m28_xor_port_y_0), //o
    .port_y_1  (m28_xor_port_y_1), //o
    .port_y_2  (m28_xor_port_y_2), //o
    .port_y_3  (m28_xor_port_y_3)  //o
  );
  Multiplication_TI m29 (
    .port_x0_0 (m28_xor_port_y_0), //i
    .port_x0_1 (m28_xor_port_y_1), //i
    .port_x0_2 (m28_xor_port_y_2), //i
    .port_x0_3 (m28_xor_port_y_3), //i
    .port_x1_0 (m27_0           ), //i
    .port_x1_1 (m27_1           ), //i
    .port_x1_2 (m27_2           ), //i
    .port_x1_3 (m27_3           ), //i
    .port_y_0  (m29_port_y_0    ), //o
    .port_y_1  (m29_port_y_1    ), //o
    .port_y_2  (m29_port_y_2    ), //o
    .port_y_3  (m29_port_y_3    ), //o
    .clk       (clk             ), //i
    .reset     (reset           )  //i
  );
  Multiplication_TI m30 (
    .port_x0_0 (m26_xor_port_y_0), //i
    .port_x0_1 (m26_xor_port_y_1), //i
    .port_x0_2 (m26_xor_port_y_2), //i
    .port_x0_3 (m26_xor_port_y_3), //i
    .port_x1_0 (m24_0           ), //i
    .port_x1_1 (m24_1           ), //i
    .port_x1_2 (m24_2           ), //i
    .port_x1_3 (m24_3           ), //i
    .port_y_0  (m30_port_y_0    ), //o
    .port_y_1  (m30_port_y_1    ), //o
    .port_y_2  (m30_port_y_2    ), //o
    .port_y_3  (m30_port_y_3    ), //o
    .clk       (clk             ), //i
    .reset     (reset           )  //i
  );
  Multiplication_TI m32 (
    .port_x0_0 (m27_0       ), //i
    .port_x0_1 (m27_1       ), //i
    .port_x0_2 (m27_2       ), //i
    .port_x0_3 (m27_3       ), //i
    .port_x1_0 (m31_port_y_0), //i
    .port_x1_1 (m31_port_y_1), //i
    .port_x1_2 (m31_port_y_2), //i
    .port_x1_3 (m31_port_y_3), //i
    .port_y_0  (m32_port_y_0), //o
    .port_y_1  (m32_port_y_1), //o
    .port_y_2  (m32_port_y_2), //o
    .port_y_3  (m32_port_y_3), //o
    .clk       (clk         ), //i
    .reset     (reset       )  //i
  );
  Addition_TI m33_xor (
    .port_x0_0 (m27_0           ), //i
    .port_x0_1 (m27_1           ), //i
    .port_x0_2 (m27_2           ), //i
    .port_x0_3 (m27_3           ), //i
    .port_x1_0 (m25_port_y_0    ), //i
    .port_x1_1 (m25_port_y_1    ), //i
    .port_x1_2 (m25_port_y_2    ), //i
    .port_x1_3 (m25_port_y_3    ), //i
    .port_y_0  (m33_xor_port_y_0), //o
    .port_y_1  (m33_xor_port_y_1), //o
    .port_y_2  (m33_xor_port_y_2), //o
    .port_y_3  (m33_xor_port_y_3)  //o
  );
  Multiplication_TI m35 (
    .port_x0_0 (m24_0       ), //i
    .port_x0_1 (m24_1       ), //i
    .port_x0_2 (m24_2       ), //i
    .port_x0_3 (m24_3       ), //i
    .port_x1_0 (m34_port_y_0), //i
    .port_x1_1 (m34_port_y_1), //i
    .port_x1_2 (m34_port_y_2), //i
    .port_x1_3 (m34_port_y_3), //i
    .port_y_0  (m35_port_y_0), //o
    .port_y_1  (m35_port_y_1), //o
    .port_y_2  (m35_port_y_2), //o
    .port_y_3  (m35_port_y_3), //o
    .clk       (clk         ), //i
    .reset     (reset       )  //i
  );
  Addition_TI m36_xor (
    .port_x0_0 (m24_0           ), //i
    .port_x0_1 (m24_1           ), //i
    .port_x0_2 (m24_2           ), //i
    .port_x0_3 (m24_3           ), //i
    .port_x1_0 (m25_port_y_0    ), //i
    .port_x1_1 (m25_port_y_1    ), //i
    .port_x1_2 (m25_port_y_2    ), //i
    .port_x1_3 (m25_port_y_3    ), //i
    .port_y_0  (m36_xor_port_y_0), //o
    .port_y_1  (m36_xor_port_y_1), //o
    .port_y_2  (m36_xor_port_y_2), //o
    .port_y_3  (m36_xor_port_y_3)  //o
  );
  Addition_TI m37_xor (
    .port_x0_0 (m21_1_0         ), //i
    .port_x0_1 (m21_1_1         ), //i
    .port_x0_2 (m21_1_2         ), //i
    .port_x0_3 (m21_1_3         ), //i
    .port_x1_0 (m29_port_y_0    ), //i
    .port_x1_1 (m29_port_y_1    ), //i
    .port_x1_2 (m29_port_y_2    ), //i
    .port_x1_3 (m29_port_y_3    ), //i
    .port_y_0  (m37_xor_port_y_0), //o
    .port_y_1  (m37_xor_port_y_1), //o
    .port_y_2  (m37_xor_port_y_2), //o
    .port_y_3  (m37_xor_port_y_3)  //o
  );
  Addition_TI m38_xor (
    .port_x0_0 (m32_port_y_0    ), //i
    .port_x0_1 (m32_port_y_1    ), //i
    .port_x0_2 (m32_port_y_2    ), //i
    .port_x0_3 (m32_port_y_3    ), //i
    .port_x1_0 (m33_0           ), //i
    .port_x1_1 (m33_1           ), //i
    .port_x1_2 (m33_2           ), //i
    .port_x1_3 (m33_3           ), //i
    .port_y_0  (m38_xor_port_y_0), //o
    .port_y_1  (m38_xor_port_y_1), //o
    .port_y_2  (m38_xor_port_y_2), //o
    .port_y_3  (m38_xor_port_y_3)  //o
  );
  Addition_TI m39_xor (
    .port_x0_0 (m23_1_0         ), //i
    .port_x0_1 (m23_1_1         ), //i
    .port_x0_2 (m23_1_2         ), //i
    .port_x0_3 (m23_1_3         ), //i
    .port_x1_0 (m30_port_y_0    ), //i
    .port_x1_1 (m30_port_y_1    ), //i
    .port_x1_2 (m30_port_y_2    ), //i
    .port_x1_3 (m30_port_y_3    ), //i
    .port_y_0  (m39_xor_port_y_0), //o
    .port_y_1  (m39_xor_port_y_1), //o
    .port_y_2  (m39_xor_port_y_2), //o
    .port_y_3  (m39_xor_port_y_3)  //o
  );
  Addition_TI m40_xor (
    .port_x0_0 (m35_port_y_0    ), //i
    .port_x0_1 (m35_port_y_1    ), //i
    .port_x0_2 (m35_port_y_2    ), //i
    .port_x0_3 (m35_port_y_3    ), //i
    .port_x1_0 (m36_0           ), //i
    .port_x1_1 (m36_1           ), //i
    .port_x1_2 (m36_2           ), //i
    .port_x1_3 (m36_3           ), //i
    .port_y_0  (m40_xor_port_y_0), //o
    .port_y_1  (m40_xor_port_y_1), //o
    .port_y_2  (m40_xor_port_y_2), //o
    .port_y_3  (m40_xor_port_y_3)  //o
  );
  Addition_TI m41_xor (
    .port_x0_0 (m38_xor_port_y_0), //i
    .port_x0_1 (m38_xor_port_y_1), //i
    .port_x0_2 (m38_xor_port_y_2), //i
    .port_x0_3 (m38_xor_port_y_3), //i
    .port_x1_0 (m40_xor_port_y_0), //i
    .port_x1_1 (m40_xor_port_y_1), //i
    .port_x1_2 (m40_xor_port_y_2), //i
    .port_x1_3 (m40_xor_port_y_3), //i
    .port_y_0  (m41_xor_port_y_0), //o
    .port_y_1  (m41_xor_port_y_1), //o
    .port_y_2  (m41_xor_port_y_2), //o
    .port_y_3  (m41_xor_port_y_3)  //o
  );
  Addition_TI m42_xor (
    .port_x0_0 (m37_xor_port_y_0), //i
    .port_x0_1 (m37_xor_port_y_1), //i
    .port_x0_2 (m37_xor_port_y_2), //i
    .port_x0_3 (m37_xor_port_y_3), //i
    .port_x1_0 (m39_xor_port_y_0), //i
    .port_x1_1 (m39_xor_port_y_1), //i
    .port_x1_2 (m39_xor_port_y_2), //i
    .port_x1_3 (m39_xor_port_y_3), //i
    .port_y_0  (m42_xor_port_y_0), //o
    .port_y_1  (m42_xor_port_y_1), //o
    .port_y_2  (m42_xor_port_y_2), //o
    .port_y_3  (m42_xor_port_y_3)  //o
  );
  Addition_TI m43_xor (
    .port_x0_0 (m37_xor_port_y_0), //i
    .port_x0_1 (m37_xor_port_y_1), //i
    .port_x0_2 (m37_xor_port_y_2), //i
    .port_x0_3 (m37_xor_port_y_3), //i
    .port_x1_0 (m38_xor_port_y_0), //i
    .port_x1_1 (m38_xor_port_y_1), //i
    .port_x1_2 (m38_xor_port_y_2), //i
    .port_x1_3 (m38_xor_port_y_3), //i
    .port_y_0  (m43_xor_port_y_0), //o
    .port_y_1  (m43_xor_port_y_1), //o
    .port_y_2  (m43_xor_port_y_2), //o
    .port_y_3  (m43_xor_port_y_3)  //o
  );
  Addition_TI m44_xor (
    .port_x0_0 (m39_xor_port_y_0), //i
    .port_x0_1 (m39_xor_port_y_1), //i
    .port_x0_2 (m39_xor_port_y_2), //i
    .port_x0_3 (m39_xor_port_y_3), //i
    .port_x1_0 (m40_xor_port_y_0), //i
    .port_x1_1 (m40_xor_port_y_1), //i
    .port_x1_2 (m40_xor_port_y_2), //i
    .port_x1_3 (m40_xor_port_y_3), //i
    .port_y_0  (m44_xor_port_y_0), //o
    .port_y_1  (m44_xor_port_y_1), //o
    .port_y_2  (m44_xor_port_y_2), //o
    .port_y_3  (m44_xor_port_y_3)  //o
  );
  Addition_TI m45_xor (
    .port_x0_0 (m42_xor_port_y_0), //i
    .port_x0_1 (m42_xor_port_y_1), //i
    .port_x0_2 (m42_xor_port_y_2), //i
    .port_x0_3 (m42_xor_port_y_3), //i
    .port_x1_0 (m41_xor_port_y_0), //i
    .port_x1_1 (m41_xor_port_y_1), //i
    .port_x1_2 (m41_xor_port_y_2), //i
    .port_x1_3 (m41_xor_port_y_3), //i
    .port_y_0  (m45_xor_port_y_0), //o
    .port_y_1  (m45_xor_port_y_1), //o
    .port_y_2  (m45_xor_port_y_2), //o
    .port_y_3  (m45_xor_port_y_3)  //o
  );
  Multiplication_TI_noReg m46_mul (
    .port_x0_0 (m44_xor_port_y_0), //i
    .port_x0_1 (m44_xor_port_y_1), //i
    .port_x0_2 (m44_xor_port_y_2), //i
    .port_x0_3 (m44_xor_port_y_3), //i
    .port_x1_0 (t6_2_0          ), //i
    .port_x1_1 (t6_2_1          ), //i
    .port_x1_2 (t6_2_2          ), //i
    .port_x1_3 (t6_2_3          ), //i
    .port_y_0  (m46_mul_port_y_0), //o
    .port_y_1  (m46_mul_port_y_1), //o
    .port_y_2  (m46_mul_port_y_2), //o
    .port_y_3  (m46_mul_port_y_3)  //o
  );
  Multiplication_TI_noReg m47_mul (
    .port_x0_0 (m40_xor_port_y_0), //i
    .port_x0_1 (m40_xor_port_y_1), //i
    .port_x0_2 (m40_xor_port_y_2), //i
    .port_x0_3 (m40_xor_port_y_3), //i
    .port_x1_0 (t8_2_0          ), //i
    .port_x1_1 (t8_2_1          ), //i
    .port_x1_2 (t8_2_2          ), //i
    .port_x1_3 (t8_2_3          ), //i
    .port_y_0  (m47_mul_port_y_0), //o
    .port_y_1  (m47_mul_port_y_1), //o
    .port_y_2  (m47_mul_port_y_2), //o
    .port_y_3  (m47_mul_port_y_3)  //o
  );
  Multiplication_TI_noReg m48_mul (
    .port_x0_0 (m39_xor_port_y_0), //i
    .port_x0_1 (m39_xor_port_y_1), //i
    .port_x0_2 (m39_xor_port_y_2), //i
    .port_x0_3 (m39_xor_port_y_3), //i
    .port_x1_0 (x7_2_0          ), //i
    .port_x1_1 (x7_2_1          ), //i
    .port_x1_2 (x7_2_2          ), //i
    .port_x1_3 (x7_2_3          ), //i
    .port_y_0  (m48_mul_port_y_0), //o
    .port_y_1  (m48_mul_port_y_1), //o
    .port_y_2  (m48_mul_port_y_2), //o
    .port_y_3  (m48_mul_port_y_3)  //o
  );
  Multiplication_TI_noReg m49_mul (
    .port_x0_0 (m43_xor_port_y_0), //i
    .port_x0_1 (m43_xor_port_y_1), //i
    .port_x0_2 (m43_xor_port_y_2), //i
    .port_x0_3 (m43_xor_port_y_3), //i
    .port_x1_0 (t16_1_0         ), //i
    .port_x1_1 (t16_1_1         ), //i
    .port_x1_2 (t16_1_2         ), //i
    .port_x1_3 (t16_1_3         ), //i
    .port_y_0  (m49_mul_port_y_0), //o
    .port_y_1  (m49_mul_port_y_1), //o
    .port_y_2  (m49_mul_port_y_2), //o
    .port_y_3  (m49_mul_port_y_3)  //o
  );
  Multiplication_TI_noReg m50_mul (
    .port_x0_0 (m38_xor_port_y_0), //i
    .port_x0_1 (m38_xor_port_y_1), //i
    .port_x0_2 (m38_xor_port_y_2), //i
    .port_x0_3 (m38_xor_port_y_3), //i
    .port_x1_0 (t9_2_0          ), //i
    .port_x1_1 (t9_2_1          ), //i
    .port_x1_2 (t9_2_2          ), //i
    .port_x1_3 (t9_2_3          ), //i
    .port_y_0  (m50_mul_port_y_0), //o
    .port_y_1  (m50_mul_port_y_1), //o
    .port_y_2  (m50_mul_port_y_2), //o
    .port_y_3  (m50_mul_port_y_3)  //o
  );
  Multiplication_TI_noReg m51_mul (
    .port_x0_0 (m37_xor_port_y_0), //i
    .port_x0_1 (m37_xor_port_y_1), //i
    .port_x0_2 (m37_xor_port_y_2), //i
    .port_x0_3 (m37_xor_port_y_3), //i
    .port_x1_0 (t17_2_0         ), //i
    .port_x1_1 (t17_2_1         ), //i
    .port_x1_2 (t17_2_2         ), //i
    .port_x1_3 (t17_2_3         ), //i
    .port_y_0  (m51_mul_port_y_0), //o
    .port_y_1  (m51_mul_port_y_1), //o
    .port_y_2  (m51_mul_port_y_2), //o
    .port_y_3  (m51_mul_port_y_3)  //o
  );
  Multiplication_TI_noReg m52_mul (
    .port_x0_0 (m42_xor_port_y_0), //i
    .port_x0_1 (m42_xor_port_y_1), //i
    .port_x0_2 (m42_xor_port_y_2), //i
    .port_x0_3 (m42_xor_port_y_3), //i
    .port_x1_0 (t15_2_0         ), //i
    .port_x1_1 (t15_2_1         ), //i
    .port_x1_2 (t15_2_2         ), //i
    .port_x1_3 (t15_2_3         ), //i
    .port_y_0  (m52_mul_port_y_0), //o
    .port_y_1  (m52_mul_port_y_1), //o
    .port_y_2  (m52_mul_port_y_2), //o
    .port_y_3  (m52_mul_port_y_3)  //o
  );
  Multiplication_TI_noReg m53_mul (
    .port_x0_0 (m45_xor_port_y_0), //i
    .port_x0_1 (m45_xor_port_y_1), //i
    .port_x0_2 (m45_xor_port_y_2), //i
    .port_x0_3 (m45_xor_port_y_3), //i
    .port_x1_0 (t27_2_0         ), //i
    .port_x1_1 (t27_2_1         ), //i
    .port_x1_2 (t27_2_2         ), //i
    .port_x1_3 (t27_2_3         ), //i
    .port_y_0  (m53_mul_port_y_0), //o
    .port_y_1  (m53_mul_port_y_1), //o
    .port_y_2  (m53_mul_port_y_2), //o
    .port_y_3  (m53_mul_port_y_3)  //o
  );
  Multiplication_TI_noReg m54_mul (
    .port_x0_0 (m41_xor_port_y_0), //i
    .port_x0_1 (m41_xor_port_y_1), //i
    .port_x0_2 (m41_xor_port_y_2), //i
    .port_x0_3 (m41_xor_port_y_3), //i
    .port_x1_0 (t10_2_0         ), //i
    .port_x1_1 (t10_2_1         ), //i
    .port_x1_2 (t10_2_2         ), //i
    .port_x1_3 (t10_2_3         ), //i
    .port_y_0  (m54_mul_port_y_0), //o
    .port_y_1  (m54_mul_port_y_1), //o
    .port_y_2  (m54_mul_port_y_2), //o
    .port_y_3  (m54_mul_port_y_3)  //o
  );
  Multiplication_TI_noReg m55_mul (
    .port_x0_0 (m44_xor_port_y_0), //i
    .port_x0_1 (m44_xor_port_y_1), //i
    .port_x0_2 (m44_xor_port_y_2), //i
    .port_x0_3 (m44_xor_port_y_3), //i
    .port_x1_0 (t13_2_0         ), //i
    .port_x1_1 (t13_2_1         ), //i
    .port_x1_2 (t13_2_2         ), //i
    .port_x1_3 (t13_2_3         ), //i
    .port_y_0  (m55_mul_port_y_0), //o
    .port_y_1  (m55_mul_port_y_1), //o
    .port_y_2  (m55_mul_port_y_2), //o
    .port_y_3  (m55_mul_port_y_3)  //o
  );
  Multiplication_TI_noReg m56_mul (
    .port_x0_0 (m40_xor_port_y_0), //i
    .port_x0_1 (m40_xor_port_y_1), //i
    .port_x0_2 (m40_xor_port_y_2), //i
    .port_x0_3 (m40_xor_port_y_3), //i
    .port_x1_0 (t23_2_0         ), //i
    .port_x1_1 (t23_2_1         ), //i
    .port_x1_2 (t23_2_2         ), //i
    .port_x1_3 (t23_2_3         ), //i
    .port_y_0  (m56_mul_port_y_0), //o
    .port_y_1  (m56_mul_port_y_1), //o
    .port_y_2  (m56_mul_port_y_2), //o
    .port_y_3  (m56_mul_port_y_3)  //o
  );
  Multiplication_TI_noReg m57_mul (
    .port_x0_0 (m39_xor_port_y_0), //i
    .port_x0_1 (m39_xor_port_y_1), //i
    .port_x0_2 (m39_xor_port_y_2), //i
    .port_x0_3 (m39_xor_port_y_3), //i
    .port_x1_0 (t19_2_0         ), //i
    .port_x1_1 (t19_2_1         ), //i
    .port_x1_2 (t19_2_2         ), //i
    .port_x1_3 (t19_2_3         ), //i
    .port_y_0  (m57_mul_port_y_0), //o
    .port_y_1  (m57_mul_port_y_1), //o
    .port_y_2  (m57_mul_port_y_2), //o
    .port_y_3  (m57_mul_port_y_3)  //o
  );
  Multiplication_TI_noReg m58_mul (
    .port_x0_0 (m43_xor_port_y_0), //i
    .port_x0_1 (m43_xor_port_y_1), //i
    .port_x0_2 (m43_xor_port_y_2), //i
    .port_x0_3 (m43_xor_port_y_3), //i
    .port_x1_0 (t3_2_0          ), //i
    .port_x1_1 (t3_2_1          ), //i
    .port_x1_2 (t3_2_2          ), //i
    .port_x1_3 (t3_2_3          ), //i
    .port_y_0  (m58_mul_port_y_0), //o
    .port_y_1  (m58_mul_port_y_1), //o
    .port_y_2  (m58_mul_port_y_2), //o
    .port_y_3  (m58_mul_port_y_3)  //o
  );
  Multiplication_TI_noReg m59_mul (
    .port_x0_0 (m38_xor_port_y_0), //i
    .port_x0_1 (m38_xor_port_y_1), //i
    .port_x0_2 (m38_xor_port_y_2), //i
    .port_x0_3 (m38_xor_port_y_3), //i
    .port_x1_0 (t22_2_0         ), //i
    .port_x1_1 (t22_2_1         ), //i
    .port_x1_2 (t22_2_2         ), //i
    .port_x1_3 (t22_2_3         ), //i
    .port_y_0  (m59_mul_port_y_0), //o
    .port_y_1  (m59_mul_port_y_1), //o
    .port_y_2  (m59_mul_port_y_2), //o
    .port_y_3  (m59_mul_port_y_3)  //o
  );
  Multiplication_TI_noReg m60_mul (
    .port_x0_0 (m37_xor_port_y_0), //i
    .port_x0_1 (m37_xor_port_y_1), //i
    .port_x0_2 (m37_xor_port_y_2), //i
    .port_x0_3 (m37_xor_port_y_3), //i
    .port_x1_0 (t20_2_0         ), //i
    .port_x1_1 (t20_2_1         ), //i
    .port_x1_2 (t20_2_2         ), //i
    .port_x1_3 (t20_2_3         ), //i
    .port_y_0  (m60_mul_port_y_0), //o
    .port_y_1  (m60_mul_port_y_1), //o
    .port_y_2  (m60_mul_port_y_2), //o
    .port_y_3  (m60_mul_port_y_3)  //o
  );
  Multiplication_TI_noReg m61_mul (
    .port_x0_0 (m42_xor_port_y_0), //i
    .port_x0_1 (m42_xor_port_y_1), //i
    .port_x0_2 (m42_xor_port_y_2), //i
    .port_x0_3 (m42_xor_port_y_3), //i
    .port_x1_0 (t1_2_0          ), //i
    .port_x1_1 (t1_2_1          ), //i
    .port_x1_2 (t1_2_2          ), //i
    .port_x1_3 (t1_2_3          ), //i
    .port_y_0  (m61_mul_port_y_0), //o
    .port_y_1  (m61_mul_port_y_1), //o
    .port_y_2  (m61_mul_port_y_2), //o
    .port_y_3  (m61_mul_port_y_3)  //o
  );
  Multiplication_TI_noReg m62_mul (
    .port_x0_0 (m45_xor_port_y_0), //i
    .port_x0_1 (m45_xor_port_y_1), //i
    .port_x0_2 (m45_xor_port_y_2), //i
    .port_x0_3 (m45_xor_port_y_3), //i
    .port_x1_0 (t4_2_0          ), //i
    .port_x1_1 (t4_2_1          ), //i
    .port_x1_2 (t4_2_2          ), //i
    .port_x1_3 (t4_2_3          ), //i
    .port_y_0  (m62_mul_port_y_0), //o
    .port_y_1  (m62_mul_port_y_1), //o
    .port_y_2  (m62_mul_port_y_2), //o
    .port_y_3  (m62_mul_port_y_3)  //o
  );
  Multiplication_TI_noReg m63_mul (
    .port_x0_0 (m41_xor_port_y_0), //i
    .port_x0_1 (m41_xor_port_y_1), //i
    .port_x0_2 (m41_xor_port_y_2), //i
    .port_x0_3 (m41_xor_port_y_3), //i
    .port_x1_0 (t2_2_0          ), //i
    .port_x1_1 (t2_2_1          ), //i
    .port_x1_2 (t2_2_2          ), //i
    .port_x1_3 (t2_2_3          ), //i
    .port_y_0  (m63_mul_port_y_0), //o
    .port_y_1  (m63_mul_port_y_1), //o
    .port_y_2  (m63_mul_port_y_2), //o
    .port_y_3  (m63_mul_port_y_3)  //o
  );
  Addition_TI l0_xor (
    .port_x0_0 (m61_mul_port_y_0), //i
    .port_x0_1 (m61_mul_port_y_1), //i
    .port_x0_2 (m61_mul_port_y_2), //i
    .port_x0_3 (m61_mul_port_y_3), //i
    .port_x1_0 (m62_mul_port_y_0), //i
    .port_x1_1 (m62_mul_port_y_1), //i
    .port_x1_2 (m62_mul_port_y_2), //i
    .port_x1_3 (m62_mul_port_y_3), //i
    .port_y_0  (l0_xor_port_y_0 ), //o
    .port_y_1  (l0_xor_port_y_1 ), //o
    .port_y_2  (l0_xor_port_y_2 ), //o
    .port_y_3  (l0_xor_port_y_3 )  //o
  );
  Addition_TI l1_xor (
    .port_x0_0 (m50_mul_port_y_0), //i
    .port_x0_1 (m50_mul_port_y_1), //i
    .port_x0_2 (m50_mul_port_y_2), //i
    .port_x0_3 (m50_mul_port_y_3), //i
    .port_x1_0 (m56_mul_port_y_0), //i
    .port_x1_1 (m56_mul_port_y_1), //i
    .port_x1_2 (m56_mul_port_y_2), //i
    .port_x1_3 (m56_mul_port_y_3), //i
    .port_y_0  (l1_xor_port_y_0 ), //o
    .port_y_1  (l1_xor_port_y_1 ), //o
    .port_y_2  (l1_xor_port_y_2 ), //o
    .port_y_3  (l1_xor_port_y_3 )  //o
  );
  Addition_TI l2_xor (
    .port_x0_0 (m46_mul_port_y_0), //i
    .port_x0_1 (m46_mul_port_y_1), //i
    .port_x0_2 (m46_mul_port_y_2), //i
    .port_x0_3 (m46_mul_port_y_3), //i
    .port_x1_0 (m48_mul_port_y_0), //i
    .port_x1_1 (m48_mul_port_y_1), //i
    .port_x1_2 (m48_mul_port_y_2), //i
    .port_x1_3 (m48_mul_port_y_3), //i
    .port_y_0  (l2_xor_port_y_0 ), //o
    .port_y_1  (l2_xor_port_y_1 ), //o
    .port_y_2  (l2_xor_port_y_2 ), //o
    .port_y_3  (l2_xor_port_y_3 )  //o
  );
  Addition_TI l3_xor (
    .port_x0_0 (m47_mul_port_y_0), //i
    .port_x0_1 (m47_mul_port_y_1), //i
    .port_x0_2 (m47_mul_port_y_2), //i
    .port_x0_3 (m47_mul_port_y_3), //i
    .port_x1_0 (m55_mul_port_y_0), //i
    .port_x1_1 (m55_mul_port_y_1), //i
    .port_x1_2 (m55_mul_port_y_2), //i
    .port_x1_3 (m55_mul_port_y_3), //i
    .port_y_0  (l3_xor_port_y_0 ), //o
    .port_y_1  (l3_xor_port_y_1 ), //o
    .port_y_2  (l3_xor_port_y_2 ), //o
    .port_y_3  (l3_xor_port_y_3 )  //o
  );
  Addition_TI l4_xor (
    .port_x0_0 (m54_mul_port_y_0), //i
    .port_x0_1 (m54_mul_port_y_1), //i
    .port_x0_2 (m54_mul_port_y_2), //i
    .port_x0_3 (m54_mul_port_y_3), //i
    .port_x1_0 (m58_mul_port_y_0), //i
    .port_x1_1 (m58_mul_port_y_1), //i
    .port_x1_2 (m58_mul_port_y_2), //i
    .port_x1_3 (m58_mul_port_y_3), //i
    .port_y_0  (l4_xor_port_y_0 ), //o
    .port_y_1  (l4_xor_port_y_1 ), //o
    .port_y_2  (l4_xor_port_y_2 ), //o
    .port_y_3  (l4_xor_port_y_3 )  //o
  );
  Addition_TI l5_xor (
    .port_x0_0 (m49_mul_port_y_0), //i
    .port_x0_1 (m49_mul_port_y_1), //i
    .port_x0_2 (m49_mul_port_y_2), //i
    .port_x0_3 (m49_mul_port_y_3), //i
    .port_x1_0 (m61_mul_port_y_0), //i
    .port_x1_1 (m61_mul_port_y_1), //i
    .port_x1_2 (m61_mul_port_y_2), //i
    .port_x1_3 (m61_mul_port_y_3), //i
    .port_y_0  (l5_xor_port_y_0 ), //o
    .port_y_1  (l5_xor_port_y_1 ), //o
    .port_y_2  (l5_xor_port_y_2 ), //o
    .port_y_3  (l5_xor_port_y_3 )  //o
  );
  Addition_TI l6_xor (
    .port_x0_0 (m62_mul_port_y_0), //i
    .port_x0_1 (m62_mul_port_y_1), //i
    .port_x0_2 (m62_mul_port_y_2), //i
    .port_x0_3 (m62_mul_port_y_3), //i
    .port_x1_0 (l5_xor_port_y_0 ), //i
    .port_x1_1 (l5_xor_port_y_1 ), //i
    .port_x1_2 (l5_xor_port_y_2 ), //i
    .port_x1_3 (l5_xor_port_y_3 ), //i
    .port_y_0  (l6_xor_port_y_0 ), //o
    .port_y_1  (l6_xor_port_y_1 ), //o
    .port_y_2  (l6_xor_port_y_2 ), //o
    .port_y_3  (l6_xor_port_y_3 )  //o
  );
  Addition_TI l7_xor (
    .port_x0_0 (m46_mul_port_y_0), //i
    .port_x0_1 (m46_mul_port_y_1), //i
    .port_x0_2 (m46_mul_port_y_2), //i
    .port_x0_3 (m46_mul_port_y_3), //i
    .port_x1_0 (l3_xor_port_y_0 ), //i
    .port_x1_1 (l3_xor_port_y_1 ), //i
    .port_x1_2 (l3_xor_port_y_2 ), //i
    .port_x1_3 (l3_xor_port_y_3 ), //i
    .port_y_0  (l7_xor_port_y_0 ), //o
    .port_y_1  (l7_xor_port_y_1 ), //o
    .port_y_2  (l7_xor_port_y_2 ), //o
    .port_y_3  (l7_xor_port_y_3 )  //o
  );
  Addition_TI l8_xor (
    .port_x0_0 (m51_mul_port_y_0), //i
    .port_x0_1 (m51_mul_port_y_1), //i
    .port_x0_2 (m51_mul_port_y_2), //i
    .port_x0_3 (m51_mul_port_y_3), //i
    .port_x1_0 (m59_mul_port_y_0), //i
    .port_x1_1 (m59_mul_port_y_1), //i
    .port_x1_2 (m59_mul_port_y_2), //i
    .port_x1_3 (m59_mul_port_y_3), //i
    .port_y_0  (l8_xor_port_y_0 ), //o
    .port_y_1  (l8_xor_port_y_1 ), //o
    .port_y_2  (l8_xor_port_y_2 ), //o
    .port_y_3  (l8_xor_port_y_3 )  //o
  );
  Addition_TI l9_xor (
    .port_x0_0 (m52_mul_port_y_0), //i
    .port_x0_1 (m52_mul_port_y_1), //i
    .port_x0_2 (m52_mul_port_y_2), //i
    .port_x0_3 (m52_mul_port_y_3), //i
    .port_x1_0 (m53_mul_port_y_0), //i
    .port_x1_1 (m53_mul_port_y_1), //i
    .port_x1_2 (m53_mul_port_y_2), //i
    .port_x1_3 (m53_mul_port_y_3), //i
    .port_y_0  (l9_xor_port_y_0 ), //o
    .port_y_1  (l9_xor_port_y_1 ), //o
    .port_y_2  (l9_xor_port_y_2 ), //o
    .port_y_3  (l9_xor_port_y_3 )  //o
  );
  Addition_TI l10_xor (
    .port_x0_0 (m53_mul_port_y_0), //i
    .port_x0_1 (m53_mul_port_y_1), //i
    .port_x0_2 (m53_mul_port_y_2), //i
    .port_x0_3 (m53_mul_port_y_3), //i
    .port_x1_0 (l4_xor_port_y_0 ), //i
    .port_x1_1 (l4_xor_port_y_1 ), //i
    .port_x1_2 (l4_xor_port_y_2 ), //i
    .port_x1_3 (l4_xor_port_y_3 ), //i
    .port_y_0  (l10_xor_port_y_0), //o
    .port_y_1  (l10_xor_port_y_1), //o
    .port_y_2  (l10_xor_port_y_2), //o
    .port_y_3  (l10_xor_port_y_3)  //o
  );
  Addition_TI l11_xor (
    .port_x0_0 (m60_mul_port_y_0), //i
    .port_x0_1 (m60_mul_port_y_1), //i
    .port_x0_2 (m60_mul_port_y_2), //i
    .port_x0_3 (m60_mul_port_y_3), //i
    .port_x1_0 (l2_xor_port_y_0 ), //i
    .port_x1_1 (l2_xor_port_y_1 ), //i
    .port_x1_2 (l2_xor_port_y_2 ), //i
    .port_x1_3 (l2_xor_port_y_3 ), //i
    .port_y_0  (l11_xor_port_y_0), //o
    .port_y_1  (l11_xor_port_y_1), //o
    .port_y_2  (l11_xor_port_y_2), //o
    .port_y_3  (l11_xor_port_y_3)  //o
  );
  Addition_TI l12_xor (
    .port_x0_0 (m48_mul_port_y_0), //i
    .port_x0_1 (m48_mul_port_y_1), //i
    .port_x0_2 (m48_mul_port_y_2), //i
    .port_x0_3 (m48_mul_port_y_3), //i
    .port_x1_0 (m51_mul_port_y_0), //i
    .port_x1_1 (m51_mul_port_y_1), //i
    .port_x1_2 (m51_mul_port_y_2), //i
    .port_x1_3 (m51_mul_port_y_3), //i
    .port_y_0  (l12_xor_port_y_0), //o
    .port_y_1  (l12_xor_port_y_1), //o
    .port_y_2  (l12_xor_port_y_2), //o
    .port_y_3  (l12_xor_port_y_3)  //o
  );
  Addition_TI l13_xor (
    .port_x0_0 (m50_mul_port_y_0), //i
    .port_x0_1 (m50_mul_port_y_1), //i
    .port_x0_2 (m50_mul_port_y_2), //i
    .port_x0_3 (m50_mul_port_y_3), //i
    .port_x1_0 (l0_xor_port_y_0 ), //i
    .port_x1_1 (l0_xor_port_y_1 ), //i
    .port_x1_2 (l0_xor_port_y_2 ), //i
    .port_x1_3 (l0_xor_port_y_3 ), //i
    .port_y_0  (l13_xor_port_y_0), //o
    .port_y_1  (l13_xor_port_y_1), //o
    .port_y_2  (l13_xor_port_y_2), //o
    .port_y_3  (l13_xor_port_y_3)  //o
  );
  Addition_TI l14_xor (
    .port_x0_0 (m52_mul_port_y_0), //i
    .port_x0_1 (m52_mul_port_y_1), //i
    .port_x0_2 (m52_mul_port_y_2), //i
    .port_x0_3 (m52_mul_port_y_3), //i
    .port_x1_0 (m61_mul_port_y_0), //i
    .port_x1_1 (m61_mul_port_y_1), //i
    .port_x1_2 (m61_mul_port_y_2), //i
    .port_x1_3 (m61_mul_port_y_3), //i
    .port_y_0  (l14_xor_port_y_0), //o
    .port_y_1  (l14_xor_port_y_1), //o
    .port_y_2  (l14_xor_port_y_2), //o
    .port_y_3  (l14_xor_port_y_3)  //o
  );
  Addition_TI l15_xor (
    .port_x0_0 (m55_mul_port_y_0), //i
    .port_x0_1 (m55_mul_port_y_1), //i
    .port_x0_2 (m55_mul_port_y_2), //i
    .port_x0_3 (m55_mul_port_y_3), //i
    .port_x1_0 (l1_xor_port_y_0 ), //i
    .port_x1_1 (l1_xor_port_y_1 ), //i
    .port_x1_2 (l1_xor_port_y_2 ), //i
    .port_x1_3 (l1_xor_port_y_3 ), //i
    .port_y_0  (l15_xor_port_y_0), //o
    .port_y_1  (l15_xor_port_y_1), //o
    .port_y_2  (l15_xor_port_y_2), //o
    .port_y_3  (l15_xor_port_y_3)  //o
  );
  Addition_TI l16_xor (
    .port_x0_0 (m56_mul_port_y_0), //i
    .port_x0_1 (m56_mul_port_y_1), //i
    .port_x0_2 (m56_mul_port_y_2), //i
    .port_x0_3 (m56_mul_port_y_3), //i
    .port_x1_0 (l0_xor_port_y_0 ), //i
    .port_x1_1 (l0_xor_port_y_1 ), //i
    .port_x1_2 (l0_xor_port_y_2 ), //i
    .port_x1_3 (l0_xor_port_y_3 ), //i
    .port_y_0  (l16_xor_port_y_0), //o
    .port_y_1  (l16_xor_port_y_1), //o
    .port_y_2  (l16_xor_port_y_2), //o
    .port_y_3  (l16_xor_port_y_3)  //o
  );
  Addition_TI l17_xor (
    .port_x0_0 (m57_mul_port_y_0), //i
    .port_x0_1 (m57_mul_port_y_1), //i
    .port_x0_2 (m57_mul_port_y_2), //i
    .port_x0_3 (m57_mul_port_y_3), //i
    .port_x1_0 (l1_xor_port_y_0 ), //i
    .port_x1_1 (l1_xor_port_y_1 ), //i
    .port_x1_2 (l1_xor_port_y_2 ), //i
    .port_x1_3 (l1_xor_port_y_3 ), //i
    .port_y_0  (l17_xor_port_y_0), //o
    .port_y_1  (l17_xor_port_y_1), //o
    .port_y_2  (l17_xor_port_y_2), //o
    .port_y_3  (l17_xor_port_y_3)  //o
  );
  Addition_TI l18_xor (
    .port_x0_0 (m58_mul_port_y_0), //i
    .port_x0_1 (m58_mul_port_y_1), //i
    .port_x0_2 (m58_mul_port_y_2), //i
    .port_x0_3 (m58_mul_port_y_3), //i
    .port_x1_0 (l8_xor_port_y_0 ), //i
    .port_x1_1 (l8_xor_port_y_1 ), //i
    .port_x1_2 (l8_xor_port_y_2 ), //i
    .port_x1_3 (l8_xor_port_y_3 ), //i
    .port_y_0  (l18_xor_port_y_0), //o
    .port_y_1  (l18_xor_port_y_1), //o
    .port_y_2  (l18_xor_port_y_2), //o
    .port_y_3  (l18_xor_port_y_3)  //o
  );
  Addition_TI l19_xor (
    .port_x0_0 (m63_mul_port_y_0), //i
    .port_x0_1 (m63_mul_port_y_1), //i
    .port_x0_2 (m63_mul_port_y_2), //i
    .port_x0_3 (m63_mul_port_y_3), //i
    .port_x1_0 (l4_xor_port_y_0 ), //i
    .port_x1_1 (l4_xor_port_y_1 ), //i
    .port_x1_2 (l4_xor_port_y_2 ), //i
    .port_x1_3 (l4_xor_port_y_3 ), //i
    .port_y_0  (l19_xor_port_y_0), //o
    .port_y_1  (l19_xor_port_y_1), //o
    .port_y_2  (l19_xor_port_y_2), //o
    .port_y_3  (l19_xor_port_y_3)  //o
  );
  Addition_TI l20_xor (
    .port_x0_0 (l0_xor_port_y_0 ), //i
    .port_x0_1 (l0_xor_port_y_1 ), //i
    .port_x0_2 (l0_xor_port_y_2 ), //i
    .port_x0_3 (l0_xor_port_y_3 ), //i
    .port_x1_0 (l1_xor_port_y_0 ), //i
    .port_x1_1 (l1_xor_port_y_1 ), //i
    .port_x1_2 (l1_xor_port_y_2 ), //i
    .port_x1_3 (l1_xor_port_y_3 ), //i
    .port_y_0  (l20_xor_port_y_0), //o
    .port_y_1  (l20_xor_port_y_1), //o
    .port_y_2  (l20_xor_port_y_2), //o
    .port_y_3  (l20_xor_port_y_3)  //o
  );
  Addition_TI l21_xor (
    .port_x0_0 (l1_xor_port_y_0 ), //i
    .port_x0_1 (l1_xor_port_y_1 ), //i
    .port_x0_2 (l1_xor_port_y_2 ), //i
    .port_x0_3 (l1_xor_port_y_3 ), //i
    .port_x1_0 (l7_xor_port_y_0 ), //i
    .port_x1_1 (l7_xor_port_y_1 ), //i
    .port_x1_2 (l7_xor_port_y_2 ), //i
    .port_x1_3 (l7_xor_port_y_3 ), //i
    .port_y_0  (l21_xor_port_y_0), //o
    .port_y_1  (l21_xor_port_y_1), //o
    .port_y_2  (l21_xor_port_y_2), //o
    .port_y_3  (l21_xor_port_y_3)  //o
  );
  Addition_TI l22_xor (
    .port_x0_0 (l3_xor_port_y_0 ), //i
    .port_x0_1 (l3_xor_port_y_1 ), //i
    .port_x0_2 (l3_xor_port_y_2 ), //i
    .port_x0_3 (l3_xor_port_y_3 ), //i
    .port_x1_0 (l12_xor_port_y_0), //i
    .port_x1_1 (l12_xor_port_y_1), //i
    .port_x1_2 (l12_xor_port_y_2), //i
    .port_x1_3 (l12_xor_port_y_3), //i
    .port_y_0  (l22_xor_port_y_0), //o
    .port_y_1  (l22_xor_port_y_1), //o
    .port_y_2  (l22_xor_port_y_2), //o
    .port_y_3  (l22_xor_port_y_3)  //o
  );
  Addition_TI l23_xor (
    .port_x0_0 (l18_xor_port_y_0), //i
    .port_x0_1 (l18_xor_port_y_1), //i
    .port_x0_2 (l18_xor_port_y_2), //i
    .port_x0_3 (l18_xor_port_y_3), //i
    .port_x1_0 (l2_xor_port_y_0 ), //i
    .port_x1_1 (l2_xor_port_y_1 ), //i
    .port_x1_2 (l2_xor_port_y_2 ), //i
    .port_x1_3 (l2_xor_port_y_3 ), //i
    .port_y_0  (l23_xor_port_y_0), //o
    .port_y_1  (l23_xor_port_y_1), //o
    .port_y_2  (l23_xor_port_y_2), //o
    .port_y_3  (l23_xor_port_y_3)  //o
  );
  Addition_TI l24_xor (
    .port_x0_0 (l15_xor_port_y_0), //i
    .port_x0_1 (l15_xor_port_y_1), //i
    .port_x0_2 (l15_xor_port_y_2), //i
    .port_x0_3 (l15_xor_port_y_3), //i
    .port_x1_0 (l9_xor_port_y_0 ), //i
    .port_x1_1 (l9_xor_port_y_1 ), //i
    .port_x1_2 (l9_xor_port_y_2 ), //i
    .port_x1_3 (l9_xor_port_y_3 ), //i
    .port_y_0  (l24_xor_port_y_0), //o
    .port_y_1  (l24_xor_port_y_1), //o
    .port_y_2  (l24_xor_port_y_2), //o
    .port_y_3  (l24_xor_port_y_3)  //o
  );
  Addition_TI l25_xor (
    .port_x0_0 (l6_xor_port_y_0 ), //i
    .port_x0_1 (l6_xor_port_y_1 ), //i
    .port_x0_2 (l6_xor_port_y_2 ), //i
    .port_x0_3 (l6_xor_port_y_3 ), //i
    .port_x1_0 (l10_xor_port_y_0), //i
    .port_x1_1 (l10_xor_port_y_1), //i
    .port_x1_2 (l10_xor_port_y_2), //i
    .port_x1_3 (l10_xor_port_y_3), //i
    .port_y_0  (l25_xor_port_y_0), //o
    .port_y_1  (l25_xor_port_y_1), //o
    .port_y_2  (l25_xor_port_y_2), //o
    .port_y_3  (l25_xor_port_y_3)  //o
  );
  Addition_TI l26_xor (
    .port_x0_0 (l7_xor_port_y_0 ), //i
    .port_x0_1 (l7_xor_port_y_1 ), //i
    .port_x0_2 (l7_xor_port_y_2 ), //i
    .port_x0_3 (l7_xor_port_y_3 ), //i
    .port_x1_0 (l9_xor_port_y_0 ), //i
    .port_x1_1 (l9_xor_port_y_1 ), //i
    .port_x1_2 (l9_xor_port_y_2 ), //i
    .port_x1_3 (l9_xor_port_y_3 ), //i
    .port_y_0  (l26_xor_port_y_0), //o
    .port_y_1  (l26_xor_port_y_1), //o
    .port_y_2  (l26_xor_port_y_2), //o
    .port_y_3  (l26_xor_port_y_3)  //o
  );
  Addition_TI l27_xor (
    .port_x0_0 (l8_xor_port_y_0 ), //i
    .port_x0_1 (l8_xor_port_y_1 ), //i
    .port_x0_2 (l8_xor_port_y_2 ), //i
    .port_x0_3 (l8_xor_port_y_3 ), //i
    .port_x1_0 (l10_xor_port_y_0), //i
    .port_x1_1 (l10_xor_port_y_1), //i
    .port_x1_2 (l10_xor_port_y_2), //i
    .port_x1_3 (l10_xor_port_y_3), //i
    .port_y_0  (l27_xor_port_y_0), //o
    .port_y_1  (l27_xor_port_y_1), //o
    .port_y_2  (l27_xor_port_y_2), //o
    .port_y_3  (l27_xor_port_y_3)  //o
  );
  Addition_TI l28_xor (
    .port_x0_0 (l11_xor_port_y_0), //i
    .port_x0_1 (l11_xor_port_y_1), //i
    .port_x0_2 (l11_xor_port_y_2), //i
    .port_x0_3 (l11_xor_port_y_3), //i
    .port_x1_0 (l14_xor_port_y_0), //i
    .port_x1_1 (l14_xor_port_y_1), //i
    .port_x1_2 (l14_xor_port_y_2), //i
    .port_x1_3 (l14_xor_port_y_3), //i
    .port_y_0  (l28_xor_port_y_0), //o
    .port_y_1  (l28_xor_port_y_1), //o
    .port_y_2  (l28_xor_port_y_2), //o
    .port_y_3  (l28_xor_port_y_3)  //o
  );
  Addition_TI l29_xor (
    .port_x0_0 (l11_xor_port_y_0), //i
    .port_x0_1 (l11_xor_port_y_1), //i
    .port_x0_2 (l11_xor_port_y_2), //i
    .port_x0_3 (l11_xor_port_y_3), //i
    .port_x1_0 (l17_xor_port_y_0), //i
    .port_x1_1 (l17_xor_port_y_1), //i
    .port_x1_2 (l17_xor_port_y_2), //i
    .port_x1_3 (l17_xor_port_y_3), //i
    .port_y_0  (l29_xor_port_y_0), //o
    .port_y_1  (l29_xor_port_y_1), //o
    .port_y_2  (l29_xor_port_y_2), //o
    .port_y_3  (l29_xor_port_y_3)  //o
  );
  Addition_TI s0 (
    .port_x0_0 (l6_xor_port_y_0 ), //i
    .port_x0_1 (l6_xor_port_y_1 ), //i
    .port_x0_2 (l6_xor_port_y_2 ), //i
    .port_x0_3 (l6_xor_port_y_3 ), //i
    .port_x1_0 (l24_xor_port_y_0), //i
    .port_x1_1 (l24_xor_port_y_1), //i
    .port_x1_2 (l24_xor_port_y_2), //i
    .port_x1_3 (l24_xor_port_y_3), //i
    .port_y_0  (s0_port_y_0     ), //o
    .port_y_1  (s0_port_y_1     ), //o
    .port_y_2  (s0_port_y_2     ), //o
    .port_y_3  (s0_port_y_3     )  //o
  );
  Addition_Inv_TI s1 (
    .port_x0_0 (l16_xor_port_y_0), //i
    .port_x0_1 (l16_xor_port_y_1), //i
    .port_x0_2 (l16_xor_port_y_2), //i
    .port_x0_3 (l16_xor_port_y_3), //i
    .port_x1_0 (l26_xor_port_y_0), //i
    .port_x1_1 (l26_xor_port_y_1), //i
    .port_x1_2 (l26_xor_port_y_2), //i
    .port_x1_3 (l26_xor_port_y_3), //i
    .port_y_0  (s1_port_y_0     ), //o
    .port_y_1  (s1_port_y_1     ), //o
    .port_y_2  (s1_port_y_2     ), //o
    .port_y_3  (s1_port_y_3     )  //o
  );
  Addition_Inv_TI s2 (
    .port_x0_0 (l19_xor_port_y_0), //i
    .port_x0_1 (l19_xor_port_y_1), //i
    .port_x0_2 (l19_xor_port_y_2), //i
    .port_x0_3 (l19_xor_port_y_3), //i
    .port_x1_0 (l28_xor_port_y_0), //i
    .port_x1_1 (l28_xor_port_y_1), //i
    .port_x1_2 (l28_xor_port_y_2), //i
    .port_x1_3 (l28_xor_port_y_3), //i
    .port_y_0  (s2_port_y_0     ), //o
    .port_y_1  (s2_port_y_1     ), //o
    .port_y_2  (s2_port_y_2     ), //o
    .port_y_3  (s2_port_y_3     )  //o
  );
  Addition_TI s3 (
    .port_x0_0 (l6_xor_port_y_0 ), //i
    .port_x0_1 (l6_xor_port_y_1 ), //i
    .port_x0_2 (l6_xor_port_y_2 ), //i
    .port_x0_3 (l6_xor_port_y_3 ), //i
    .port_x1_0 (l21_xor_port_y_0), //i
    .port_x1_1 (l21_xor_port_y_1), //i
    .port_x1_2 (l21_xor_port_y_2), //i
    .port_x1_3 (l21_xor_port_y_3), //i
    .port_y_0  (s3_port_y_0     ), //o
    .port_y_1  (s3_port_y_1     ), //o
    .port_y_2  (s3_port_y_2     ), //o
    .port_y_3  (s3_port_y_3     )  //o
  );
  Addition_TI s4 (
    .port_x0_0 (l20_xor_port_y_0), //i
    .port_x0_1 (l20_xor_port_y_1), //i
    .port_x0_2 (l20_xor_port_y_2), //i
    .port_x0_3 (l20_xor_port_y_3), //i
    .port_x1_0 (l22_xor_port_y_0), //i
    .port_x1_1 (l22_xor_port_y_1), //i
    .port_x1_2 (l22_xor_port_y_2), //i
    .port_x1_3 (l22_xor_port_y_3), //i
    .port_y_0  (s4_port_y_0     ), //o
    .port_y_1  (s4_port_y_1     ), //o
    .port_y_2  (s4_port_y_2     ), //o
    .port_y_3  (s4_port_y_3     )  //o
  );
  Addition_TI s5 (
    .port_x0_0 (l25_xor_port_y_0), //i
    .port_x0_1 (l25_xor_port_y_1), //i
    .port_x0_2 (l25_xor_port_y_2), //i
    .port_x0_3 (l25_xor_port_y_3), //i
    .port_x1_0 (l29_xor_port_y_0), //i
    .port_x1_1 (l29_xor_port_y_1), //i
    .port_x1_2 (l29_xor_port_y_2), //i
    .port_x1_3 (l29_xor_port_y_3), //i
    .port_y_0  (s5_port_y_0     ), //o
    .port_y_1  (s5_port_y_1     ), //o
    .port_y_2  (s5_port_y_2     ), //o
    .port_y_3  (s5_port_y_3     )  //o
  );
  Addition_Inv_TI s6 (
    .port_x0_0 (l13_xor_port_y_0), //i
    .port_x0_1 (l13_xor_port_y_1), //i
    .port_x0_2 (l13_xor_port_y_2), //i
    .port_x0_3 (l13_xor_port_y_3), //i
    .port_x1_0 (l27_xor_port_y_0), //i
    .port_x1_1 (l27_xor_port_y_1), //i
    .port_x1_2 (l27_xor_port_y_2), //i
    .port_x1_3 (l27_xor_port_y_3), //i
    .port_y_0  (s6_port_y_0     ), //o
    .port_y_1  (s6_port_y_1     ), //o
    .port_y_2  (s6_port_y_2     ), //o
    .port_y_3  (s6_port_y_3     )  //o
  );
  Addition_Inv_TI s7 (
    .port_x0_0 (l6_xor_port_y_0 ), //i
    .port_x0_1 (l6_xor_port_y_1 ), //i
    .port_x0_2 (l6_xor_port_y_2 ), //i
    .port_x0_3 (l6_xor_port_y_3 ), //i
    .port_x1_0 (l23_xor_port_y_0), //i
    .port_x1_1 (l23_xor_port_y_1), //i
    .port_x1_2 (l23_xor_port_y_2), //i
    .port_x1_3 (l23_xor_port_y_3), //i
    .port_y_0  (s7_port_y_0     ), //o
    .port_y_1  (s7_port_y_1     ), //o
    .port_y_2  (s7_port_y_2     ), //o
    .port_y_3  (s7_port_y_3     )  //o
  );
  assign in_x0_0 = port_i_0_7;
  assign in_x1_0 = port_i_0_6;
  assign in_x2_0 = port_i_0_5;
  assign in_x3_0 = port_i_0_4;
  assign in_x4_0 = port_i_0_3;
  assign in_x5_0 = port_i_0_2;
  assign in_x6_0 = port_i_0_1;
  assign in_x7_0 = port_i_0_0;
  assign in_x0_1 = port_i_1_7;
  assign in_x1_1 = port_i_1_6;
  assign in_x2_1 = port_i_1_5;
  assign in_x3_1 = port_i_1_4;
  assign in_x4_1 = port_i_1_3;
  assign in_x5_1 = port_i_1_2;
  assign in_x6_1 = port_i_1_1;
  assign in_x7_1 = port_i_1_0;
  assign in_x0_2 = port_i_2_7;
  assign in_x1_2 = port_i_2_6;
  assign in_x2_2 = port_i_2_5;
  assign in_x3_2 = port_i_2_4;
  assign in_x4_2 = port_i_2_3;
  assign in_x5_2 = port_i_2_2;
  assign in_x6_2 = port_i_2_1;
  assign in_x7_2 = port_i_2_0;
  assign in_x0_3 = port_i_3_7;
  assign in_x1_3 = port_i_3_6;
  assign in_x2_3 = port_i_3_5;
  assign in_x3_3 = port_i_3_4;
  assign in_x4_3 = port_i_3_3;
  assign in_x5_3 = port_i_3_2;
  assign in_x6_3 = port_i_3_1;
  assign in_x7_3 = port_i_3_0;
  assign out_y0_0 = s0_port_y_0;
  assign out_y0_1 = s0_port_y_1;
  assign out_y0_2 = s0_port_y_2;
  assign out_y0_3 = s0_port_y_3;
  assign out_y1_0 = s1_port_y_0;
  assign out_y1_1 = s1_port_y_1;
  assign out_y1_2 = s1_port_y_2;
  assign out_y1_3 = s1_port_y_3;
  assign out_y2_0 = s2_port_y_0;
  assign out_y2_1 = s2_port_y_1;
  assign out_y2_2 = s2_port_y_2;
  assign out_y2_3 = s2_port_y_3;
  assign out_y3_0 = s3_port_y_0;
  assign out_y3_1 = s3_port_y_1;
  assign out_y3_2 = s3_port_y_2;
  assign out_y3_3 = s3_port_y_3;
  assign out_y4_0 = s4_port_y_0;
  assign out_y4_1 = s4_port_y_1;
  assign out_y4_2 = s4_port_y_2;
  assign out_y4_3 = s4_port_y_3;
  assign out_y5_0 = s5_port_y_0;
  assign out_y5_1 = s5_port_y_1;
  assign out_y5_2 = s5_port_y_2;
  assign out_y5_3 = s5_port_y_3;
  assign out_y6_0 = s6_port_y_0;
  assign out_y6_1 = s6_port_y_1;
  assign out_y6_2 = s6_port_y_2;
  assign out_y6_3 = s6_port_y_3;
  assign out_y7_0 = s7_port_y_0;
  assign out_y7_1 = s7_port_y_1;
  assign out_y7_2 = s7_port_y_2;
  assign out_y7_3 = s7_port_y_3;
  assign port_o_0_7 = out_y0_0;
  assign port_o_0_6 = out_y1_0;
  assign port_o_0_5 = out_y2_0;
  assign port_o_0_4 = out_y3_0;
  assign port_o_0_3 = out_y4_0;
  assign port_o_0_2 = out_y5_0;
  assign port_o_0_1 = out_y6_0;
  assign port_o_0_0 = out_y7_0;
  assign port_o_1_7 = out_y0_1;
  assign port_o_1_6 = out_y1_1;
  assign port_o_1_5 = out_y2_1;
  assign port_o_1_4 = out_y3_1;
  assign port_o_1_3 = out_y4_1;
  assign port_o_1_2 = out_y5_1;
  assign port_o_1_1 = out_y6_1;
  assign port_o_1_0 = out_y7_1;
  assign port_o_2_7 = out_y0_2;
  assign port_o_2_6 = out_y1_2;
  assign port_o_2_5 = out_y2_2;
  assign port_o_2_4 = out_y3_2;
  assign port_o_2_3 = out_y4_2;
  assign port_o_2_2 = out_y5_2;
  assign port_o_2_1 = out_y6_2;
  assign port_o_2_0 = out_y7_2;
  assign port_o_3_7 = out_y0_3;
  assign port_o_3_6 = out_y1_3;
  assign port_o_3_5 = out_y2_3;
  assign port_o_3_4 = out_y3_3;
  assign port_o_3_3 = out_y4_3;
  assign port_o_3_2 = out_y5_3;
  assign port_o_3_1 = out_y6_3;
  assign port_o_3_0 = out_y7_3;
  always @(posedge clk) begin
    x7_0 <= in_x7_0;
    x7_1 <= in_x7_1;
    x7_2 <= in_x7_2;
    x7_3 <= in_x7_3;
    t1_0 <= t1_xor_port_y_0;
    t1_1 <= t1_xor_port_y_1;
    t1_2 <= t1_xor_port_y_2;
    t1_3 <= t1_xor_port_y_3;
    t2_0 <= t2_xor_port_y_0;
    t2_1 <= t2_xor_port_y_1;
    t2_2 <= t2_xor_port_y_2;
    t2_3 <= t2_xor_port_y_3;
    t3_0 <= t3_xor_port_y_0;
    t3_1 <= t3_xor_port_y_1;
    t3_2 <= t3_xor_port_y_2;
    t3_3 <= t3_xor_port_y_3;
    t4_0 <= t4_xor_port_y_0;
    t4_1 <= t4_xor_port_y_1;
    t4_2 <= t4_xor_port_y_2;
    t4_3 <= t4_xor_port_y_3;
    t6_0 <= t6_xor_port_y_0;
    t6_1 <= t6_xor_port_y_1;
    t6_2 <= t6_xor_port_y_2;
    t6_3 <= t6_xor_port_y_3;
    t7_0 <= t7_xor_port_y_0;
    t7_1 <= t7_xor_port_y_1;
    t7_2 <= t7_xor_port_y_2;
    t7_3 <= t7_xor_port_y_3;
    t8_0 <= t8_xor_port_y_0;
    t8_1 <= t8_xor_port_y_1;
    t8_2 <= t8_xor_port_y_2;
    t8_3 <= t8_xor_port_y_3;
    t9_0 <= t9_xor_port_y_0;
    t9_1 <= t9_xor_port_y_1;
    t9_2 <= t9_xor_port_y_2;
    t9_3 <= t9_xor_port_y_3;
    t10_0 <= t10_xor_port_y_0;
    t10_1 <= t10_xor_port_y_1;
    t10_2 <= t10_xor_port_y_2;
    t10_3 <= t10_xor_port_y_3;
    t13_0 <= t13_xor_port_y_0;
    t13_1 <= t13_xor_port_y_1;
    t13_2 <= t13_xor_port_y_2;
    t13_3 <= t13_xor_port_y_3;
    t14_0 <= t14_xor_port_y_0;
    t14_1 <= t14_xor_port_y_1;
    t14_2 <= t14_xor_port_y_2;
    t14_3 <= t14_xor_port_y_3;
    t15_0 <= t15_xor_port_y_0;
    t15_1 <= t15_xor_port_y_1;
    t15_2 <= t15_xor_port_y_2;
    t15_3 <= t15_xor_port_y_3;
    t16_0 <= t16_xor_port_y_0;
    t16_1 <= t16_xor_port_y_1;
    t16_2 <= t16_xor_port_y_2;
    t16_3 <= t16_xor_port_y_3;
    t17_0 <= t17_xor_port_y_0;
    t17_1 <= t17_xor_port_y_1;
    t17_2 <= t17_xor_port_y_2;
    t17_3 <= t17_xor_port_y_3;
    t19_0 <= t19_xor_port_y_0;
    t19_1 <= t19_xor_port_y_1;
    t19_2 <= t19_xor_port_y_2;
    t19_3 <= t19_xor_port_y_3;
    t20_0 <= t20_xor_port_y_0;
    t20_1 <= t20_xor_port_y_1;
    t20_2 <= t20_xor_port_y_2;
    t20_3 <= t20_xor_port_y_3;
    t22_0 <= t22_xor_port_y_0;
    t22_1 <= t22_xor_port_y_1;
    t22_2 <= t22_xor_port_y_2;
    t22_3 <= t22_xor_port_y_3;
    t23_0 <= t23_xor_port_y_0;
    t23_1 <= t23_xor_port_y_1;
    t23_2 <= t23_xor_port_y_2;
    t23_3 <= t23_xor_port_y_3;
    t24_0 <= t24_xor_port_y_0;
    t24_1 <= t24_xor_port_y_1;
    t24_2 <= t24_xor_port_y_2;
    t24_3 <= t24_xor_port_y_3;
    t25_0 <= t25_xor_port_y_0;
    t25_1 <= t25_xor_port_y_1;
    t25_2 <= t25_xor_port_y_2;
    t25_3 <= t25_xor_port_y_3;
    t26_0 <= t26_xor_port_y_0;
    t26_1 <= t26_xor_port_y_1;
    t26_2 <= t26_xor_port_y_2;
    t26_3 <= t26_xor_port_y_3;
    t27_0 <= t27_xor_port_y_0;
    t27_1 <= t27_xor_port_y_1;
    t27_2 <= t27_xor_port_y_2;
    t27_3 <= t27_xor_port_y_3;
    x7_1_0 <= x7_0;
    x7_1_1 <= x7_1;
    x7_1_2 <= x7_2;
    x7_1_3 <= x7_3;
    t1_1_0 <= t1_0;
    t1_1_1 <= t1_1;
    t1_1_2 <= t1_2;
    t1_1_3 <= t1_3;
    t2_1_0 <= t2_0;
    t2_1_1 <= t2_1;
    t2_1_2 <= t2_2;
    t2_1_3 <= t2_3;
    t3_1_0 <= t3_0;
    t3_1_1 <= t3_1;
    t3_1_2 <= t3_2;
    t3_1_3 <= t3_3;
    t4_1_0 <= t4_0;
    t4_1_1 <= t4_1;
    t4_1_2 <= t4_2;
    t4_1_3 <= t4_3;
    t6_1_0 <= t6_0;
    t6_1_1 <= t6_1;
    t6_1_2 <= t6_2;
    t6_1_3 <= t6_3;
    t8_1_0 <= t8_0;
    t8_1_1 <= t8_1;
    t8_1_2 <= t8_2;
    t8_1_3 <= t8_3;
    t9_1_0 <= t9_0;
    t9_1_1 <= t9_1;
    t9_1_2 <= t9_2;
    t9_1_3 <= t9_3;
    t10_1_0 <= t10_0;
    t10_1_1 <= t10_1;
    t10_1_2 <= t10_2;
    t10_1_3 <= t10_3;
    t13_1_0 <= t13_0;
    t13_1_1 <= t13_1;
    t13_1_2 <= t13_2;
    t13_1_3 <= t13_3;
    t15_1_0 <= t15_0;
    t15_1_1 <= t15_1;
    t15_1_2 <= t15_2;
    t15_1_3 <= t15_3;
    t16_1_0 <= t16_0;
    t16_1_1 <= t16_1;
    t16_1_2 <= t16_2;
    t16_1_3 <= t16_3;
    t17_1_0 <= t17_0;
    t17_1_1 <= t17_1;
    t17_1_2 <= t17_2;
    t17_1_3 <= t17_3;
    t19_1_0 <= t19_0;
    t19_1_1 <= t19_1;
    t19_1_2 <= t19_2;
    t19_1_3 <= t19_3;
    t20_1_0 <= t20_0;
    t20_1_1 <= t20_1;
    t20_1_2 <= t20_2;
    t20_1_3 <= t20_3;
    t22_1_0 <= t22_0;
    t22_1_1 <= t22_1;
    t22_1_2 <= t22_2;
    t22_1_3 <= t22_3;
    t23_1_0 <= t23_0;
    t23_1_1 <= t23_1;
    t23_1_2 <= t23_2;
    t23_1_3 <= t23_3;
    t27_1_0 <= t27_0;
    t27_1_1 <= t27_1;
    t27_1_2 <= t27_2;
    t27_1_3 <= t27_3;
    m21_0 <= m21_xor_port_y_0;
    m21_1 <= m21_xor_port_y_1;
    m21_2 <= m21_xor_port_y_2;
    m21_3 <= m21_xor_port_y_3;
    m23_0 <= m23_xor_port_y_0;
    m23_1 <= m23_xor_port_y_1;
    m23_2 <= m23_xor_port_y_2;
    m23_3 <= m23_xor_port_y_3;
    m24_0 <= m24_xor_port_y_0;
    m24_1 <= m24_xor_port_y_1;
    m24_2 <= m24_xor_port_y_2;
    m24_3 <= m24_xor_port_y_3;
    m27_0 <= m27_xor_port_y_0;
    m27_1 <= m27_xor_port_y_1;
    m27_2 <= m27_xor_port_y_2;
    m27_3 <= m27_xor_port_y_3;
    x7_2_0 <= x7_1_0;
    x7_2_1 <= x7_1_1;
    x7_2_2 <= x7_1_2;
    x7_2_3 <= x7_1_3;
    t1_2_0 <= t1_1_0;
    t1_2_1 <= t1_1_1;
    t1_2_2 <= t1_1_2;
    t1_2_3 <= t1_1_3;
    t2_2_0 <= t2_1_0;
    t2_2_1 <= t2_1_1;
    t2_2_2 <= t2_1_2;
    t2_2_3 <= t2_1_3;
    t3_2_0 <= t3_1_0;
    t3_2_1 <= t3_1_1;
    t3_2_2 <= t3_1_2;
    t3_2_3 <= t3_1_3;
    t4_2_0 <= t4_1_0;
    t4_2_1 <= t4_1_1;
    t4_2_2 <= t4_1_2;
    t4_2_3 <= t4_1_3;
    t6_2_0 <= t6_1_0;
    t6_2_1 <= t6_1_1;
    t6_2_2 <= t6_1_2;
    t6_2_3 <= t6_1_3;
    t8_2_0 <= t8_1_0;
    t8_2_1 <= t8_1_1;
    t8_2_2 <= t8_1_2;
    t8_2_3 <= t8_1_3;
    t9_2_0 <= t9_1_0;
    t9_2_1 <= t9_1_1;
    t9_2_2 <= t9_1_2;
    t9_2_3 <= t9_1_3;
    t10_2_0 <= t10_1_0;
    t10_2_1 <= t10_1_1;
    t10_2_2 <= t10_1_2;
    t10_2_3 <= t10_1_3;
    t13_2_0 <= t13_1_0;
    t13_2_1 <= t13_1_1;
    t13_2_2 <= t13_1_2;
    t13_2_3 <= t13_1_3;
    t15_2_0 <= t15_1_0;
    t15_2_1 <= t15_1_1;
    t15_2_2 <= t15_1_2;
    t15_2_3 <= t15_1_3;
    t16_2_0 <= t16_1_0;
    t16_2_1 <= t16_1_1;
    t16_2_2 <= t16_1_2;
    t16_2_3 <= t16_1_3;
    t17_2_0 <= t17_1_0;
    t17_2_1 <= t17_1_1;
    t17_2_2 <= t17_1_2;
    t17_2_3 <= t17_1_3;
    t19_2_0 <= t19_1_0;
    t19_2_1 <= t19_1_1;
    t19_2_2 <= t19_1_2;
    t19_2_3 <= t19_1_3;
    t20_2_0 <= t20_1_0;
    t20_2_1 <= t20_1_1;
    t20_2_2 <= t20_1_2;
    t20_2_3 <= t20_1_3;
    t22_2_0 <= t22_1_0;
    t22_2_1 <= t22_1_1;
    t22_2_2 <= t22_1_2;
    t22_2_3 <= t22_1_3;
    t23_2_0 <= t23_1_0;
    t23_2_1 <= t23_1_1;
    t23_2_2 <= t23_1_2;
    t23_2_3 <= t23_1_3;
    t27_2_0 <= t27_1_0;
    t27_2_1 <= t27_1_1;
    t27_2_2 <= t27_1_2;
    t27_2_3 <= t27_1_3;
    m21_1_0 <= m21_0;
    m21_1_1 <= m21_1;
    m21_1_2 <= m21_2;
    m21_1_3 <= m21_3;
    m23_1_0 <= m23_0;
    m23_1_1 <= m23_1;
    m23_1_2 <= m23_2;
    m23_1_3 <= m23_3;
    m33_0 <= m33_xor_port_y_0;
    m33_1 <= m33_xor_port_y_1;
    m33_2 <= m33_xor_port_y_2;
    m33_3 <= m33_xor_port_y_3;
    m36_0 <= m36_xor_port_y_0;
    m36_1 <= m36_xor_port_y_1;
    m36_2 <= m36_xor_port_y_2;
    m36_3 <= m36_xor_port_y_3;
  end


endmodule

module AES_KeyAddition (
  input      [0:0]    port_state_in_0_0_0,
  input      [0:0]    port_state_in_0_0_1,
  input      [0:0]    port_state_in_0_0_2,
  input      [0:0]    port_state_in_0_0_3,
  input      [0:0]    port_state_in_0_0_4,
  input      [0:0]    port_state_in_0_0_5,
  input      [0:0]    port_state_in_0_0_6,
  input      [0:0]    port_state_in_0_0_7,
  input      [0:0]    port_state_in_0_1_0,
  input      [0:0]    port_state_in_0_1_1,
  input      [0:0]    port_state_in_0_1_2,
  input      [0:0]    port_state_in_0_1_3,
  input      [0:0]    port_state_in_0_1_4,
  input      [0:0]    port_state_in_0_1_5,
  input      [0:0]    port_state_in_0_1_6,
  input      [0:0]    port_state_in_0_1_7,
  input      [0:0]    port_state_in_0_2_0,
  input      [0:0]    port_state_in_0_2_1,
  input      [0:0]    port_state_in_0_2_2,
  input      [0:0]    port_state_in_0_2_3,
  input      [0:0]    port_state_in_0_2_4,
  input      [0:0]    port_state_in_0_2_5,
  input      [0:0]    port_state_in_0_2_6,
  input      [0:0]    port_state_in_0_2_7,
  input      [0:0]    port_state_in_0_3_0,
  input      [0:0]    port_state_in_0_3_1,
  input      [0:0]    port_state_in_0_3_2,
  input      [0:0]    port_state_in_0_3_3,
  input      [0:0]    port_state_in_0_3_4,
  input      [0:0]    port_state_in_0_3_5,
  input      [0:0]    port_state_in_0_3_6,
  input      [0:0]    port_state_in_0_3_7,
  input      [0:0]    port_state_in_1_0_0,
  input      [0:0]    port_state_in_1_0_1,
  input      [0:0]    port_state_in_1_0_2,
  input      [0:0]    port_state_in_1_0_3,
  input      [0:0]    port_state_in_1_0_4,
  input      [0:0]    port_state_in_1_0_5,
  input      [0:0]    port_state_in_1_0_6,
  input      [0:0]    port_state_in_1_0_7,
  input      [0:0]    port_state_in_1_1_0,
  input      [0:0]    port_state_in_1_1_1,
  input      [0:0]    port_state_in_1_1_2,
  input      [0:0]    port_state_in_1_1_3,
  input      [0:0]    port_state_in_1_1_4,
  input      [0:0]    port_state_in_1_1_5,
  input      [0:0]    port_state_in_1_1_6,
  input      [0:0]    port_state_in_1_1_7,
  input      [0:0]    port_state_in_1_2_0,
  input      [0:0]    port_state_in_1_2_1,
  input      [0:0]    port_state_in_1_2_2,
  input      [0:0]    port_state_in_1_2_3,
  input      [0:0]    port_state_in_1_2_4,
  input      [0:0]    port_state_in_1_2_5,
  input      [0:0]    port_state_in_1_2_6,
  input      [0:0]    port_state_in_1_2_7,
  input      [0:0]    port_state_in_1_3_0,
  input      [0:0]    port_state_in_1_3_1,
  input      [0:0]    port_state_in_1_3_2,
  input      [0:0]    port_state_in_1_3_3,
  input      [0:0]    port_state_in_1_3_4,
  input      [0:0]    port_state_in_1_3_5,
  input      [0:0]    port_state_in_1_3_6,
  input      [0:0]    port_state_in_1_3_7,
  input      [0:0]    port_state_in_2_0_0,
  input      [0:0]    port_state_in_2_0_1,
  input      [0:0]    port_state_in_2_0_2,
  input      [0:0]    port_state_in_2_0_3,
  input      [0:0]    port_state_in_2_0_4,
  input      [0:0]    port_state_in_2_0_5,
  input      [0:0]    port_state_in_2_0_6,
  input      [0:0]    port_state_in_2_0_7,
  input      [0:0]    port_state_in_2_1_0,
  input      [0:0]    port_state_in_2_1_1,
  input      [0:0]    port_state_in_2_1_2,
  input      [0:0]    port_state_in_2_1_3,
  input      [0:0]    port_state_in_2_1_4,
  input      [0:0]    port_state_in_2_1_5,
  input      [0:0]    port_state_in_2_1_6,
  input      [0:0]    port_state_in_2_1_7,
  input      [0:0]    port_state_in_2_2_0,
  input      [0:0]    port_state_in_2_2_1,
  input      [0:0]    port_state_in_2_2_2,
  input      [0:0]    port_state_in_2_2_3,
  input      [0:0]    port_state_in_2_2_4,
  input      [0:0]    port_state_in_2_2_5,
  input      [0:0]    port_state_in_2_2_6,
  input      [0:0]    port_state_in_2_2_7,
  input      [0:0]    port_state_in_2_3_0,
  input      [0:0]    port_state_in_2_3_1,
  input      [0:0]    port_state_in_2_3_2,
  input      [0:0]    port_state_in_2_3_3,
  input      [0:0]    port_state_in_2_3_4,
  input      [0:0]    port_state_in_2_3_5,
  input      [0:0]    port_state_in_2_3_6,
  input      [0:0]    port_state_in_2_3_7,
  input      [0:0]    port_state_in_3_0_0,
  input      [0:0]    port_state_in_3_0_1,
  input      [0:0]    port_state_in_3_0_2,
  input      [0:0]    port_state_in_3_0_3,
  input      [0:0]    port_state_in_3_0_4,
  input      [0:0]    port_state_in_3_0_5,
  input      [0:0]    port_state_in_3_0_6,
  input      [0:0]    port_state_in_3_0_7,
  input      [0:0]    port_state_in_3_1_0,
  input      [0:0]    port_state_in_3_1_1,
  input      [0:0]    port_state_in_3_1_2,
  input      [0:0]    port_state_in_3_1_3,
  input      [0:0]    port_state_in_3_1_4,
  input      [0:0]    port_state_in_3_1_5,
  input      [0:0]    port_state_in_3_1_6,
  input      [0:0]    port_state_in_3_1_7,
  input      [0:0]    port_state_in_3_2_0,
  input      [0:0]    port_state_in_3_2_1,
  input      [0:0]    port_state_in_3_2_2,
  input      [0:0]    port_state_in_3_2_3,
  input      [0:0]    port_state_in_3_2_4,
  input      [0:0]    port_state_in_3_2_5,
  input      [0:0]    port_state_in_3_2_6,
  input      [0:0]    port_state_in_3_2_7,
  input      [0:0]    port_state_in_3_3_0,
  input      [0:0]    port_state_in_3_3_1,
  input      [0:0]    port_state_in_3_3_2,
  input      [0:0]    port_state_in_3_3_3,
  input      [0:0]    port_state_in_3_3_4,
  input      [0:0]    port_state_in_3_3_5,
  input      [0:0]    port_state_in_3_3_6,
  input      [0:0]    port_state_in_3_3_7,
  input      [0:0]    port_state_in_4_0_0,
  input      [0:0]    port_state_in_4_0_1,
  input      [0:0]    port_state_in_4_0_2,
  input      [0:0]    port_state_in_4_0_3,
  input      [0:0]    port_state_in_4_0_4,
  input      [0:0]    port_state_in_4_0_5,
  input      [0:0]    port_state_in_4_0_6,
  input      [0:0]    port_state_in_4_0_7,
  input      [0:0]    port_state_in_4_1_0,
  input      [0:0]    port_state_in_4_1_1,
  input      [0:0]    port_state_in_4_1_2,
  input      [0:0]    port_state_in_4_1_3,
  input      [0:0]    port_state_in_4_1_4,
  input      [0:0]    port_state_in_4_1_5,
  input      [0:0]    port_state_in_4_1_6,
  input      [0:0]    port_state_in_4_1_7,
  input      [0:0]    port_state_in_4_2_0,
  input      [0:0]    port_state_in_4_2_1,
  input      [0:0]    port_state_in_4_2_2,
  input      [0:0]    port_state_in_4_2_3,
  input      [0:0]    port_state_in_4_2_4,
  input      [0:0]    port_state_in_4_2_5,
  input      [0:0]    port_state_in_4_2_6,
  input      [0:0]    port_state_in_4_2_7,
  input      [0:0]    port_state_in_4_3_0,
  input      [0:0]    port_state_in_4_3_1,
  input      [0:0]    port_state_in_4_3_2,
  input      [0:0]    port_state_in_4_3_3,
  input      [0:0]    port_state_in_4_3_4,
  input      [0:0]    port_state_in_4_3_5,
  input      [0:0]    port_state_in_4_3_6,
  input      [0:0]    port_state_in_4_3_7,
  input      [0:0]    port_state_in_5_0_0,
  input      [0:0]    port_state_in_5_0_1,
  input      [0:0]    port_state_in_5_0_2,
  input      [0:0]    port_state_in_5_0_3,
  input      [0:0]    port_state_in_5_0_4,
  input      [0:0]    port_state_in_5_0_5,
  input      [0:0]    port_state_in_5_0_6,
  input      [0:0]    port_state_in_5_0_7,
  input      [0:0]    port_state_in_5_1_0,
  input      [0:0]    port_state_in_5_1_1,
  input      [0:0]    port_state_in_5_1_2,
  input      [0:0]    port_state_in_5_1_3,
  input      [0:0]    port_state_in_5_1_4,
  input      [0:0]    port_state_in_5_1_5,
  input      [0:0]    port_state_in_5_1_6,
  input      [0:0]    port_state_in_5_1_7,
  input      [0:0]    port_state_in_5_2_0,
  input      [0:0]    port_state_in_5_2_1,
  input      [0:0]    port_state_in_5_2_2,
  input      [0:0]    port_state_in_5_2_3,
  input      [0:0]    port_state_in_5_2_4,
  input      [0:0]    port_state_in_5_2_5,
  input      [0:0]    port_state_in_5_2_6,
  input      [0:0]    port_state_in_5_2_7,
  input      [0:0]    port_state_in_5_3_0,
  input      [0:0]    port_state_in_5_3_1,
  input      [0:0]    port_state_in_5_3_2,
  input      [0:0]    port_state_in_5_3_3,
  input      [0:0]    port_state_in_5_3_4,
  input      [0:0]    port_state_in_5_3_5,
  input      [0:0]    port_state_in_5_3_6,
  input      [0:0]    port_state_in_5_3_7,
  input      [0:0]    port_state_in_6_0_0,
  input      [0:0]    port_state_in_6_0_1,
  input      [0:0]    port_state_in_6_0_2,
  input      [0:0]    port_state_in_6_0_3,
  input      [0:0]    port_state_in_6_0_4,
  input      [0:0]    port_state_in_6_0_5,
  input      [0:0]    port_state_in_6_0_6,
  input      [0:0]    port_state_in_6_0_7,
  input      [0:0]    port_state_in_6_1_0,
  input      [0:0]    port_state_in_6_1_1,
  input      [0:0]    port_state_in_6_1_2,
  input      [0:0]    port_state_in_6_1_3,
  input      [0:0]    port_state_in_6_1_4,
  input      [0:0]    port_state_in_6_1_5,
  input      [0:0]    port_state_in_6_1_6,
  input      [0:0]    port_state_in_6_1_7,
  input      [0:0]    port_state_in_6_2_0,
  input      [0:0]    port_state_in_6_2_1,
  input      [0:0]    port_state_in_6_2_2,
  input      [0:0]    port_state_in_6_2_3,
  input      [0:0]    port_state_in_6_2_4,
  input      [0:0]    port_state_in_6_2_5,
  input      [0:0]    port_state_in_6_2_6,
  input      [0:0]    port_state_in_6_2_7,
  input      [0:0]    port_state_in_6_3_0,
  input      [0:0]    port_state_in_6_3_1,
  input      [0:0]    port_state_in_6_3_2,
  input      [0:0]    port_state_in_6_3_3,
  input      [0:0]    port_state_in_6_3_4,
  input      [0:0]    port_state_in_6_3_5,
  input      [0:0]    port_state_in_6_3_6,
  input      [0:0]    port_state_in_6_3_7,
  input      [0:0]    port_state_in_7_0_0,
  input      [0:0]    port_state_in_7_0_1,
  input      [0:0]    port_state_in_7_0_2,
  input      [0:0]    port_state_in_7_0_3,
  input      [0:0]    port_state_in_7_0_4,
  input      [0:0]    port_state_in_7_0_5,
  input      [0:0]    port_state_in_7_0_6,
  input      [0:0]    port_state_in_7_0_7,
  input      [0:0]    port_state_in_7_1_0,
  input      [0:0]    port_state_in_7_1_1,
  input      [0:0]    port_state_in_7_1_2,
  input      [0:0]    port_state_in_7_1_3,
  input      [0:0]    port_state_in_7_1_4,
  input      [0:0]    port_state_in_7_1_5,
  input      [0:0]    port_state_in_7_1_6,
  input      [0:0]    port_state_in_7_1_7,
  input      [0:0]    port_state_in_7_2_0,
  input      [0:0]    port_state_in_7_2_1,
  input      [0:0]    port_state_in_7_2_2,
  input      [0:0]    port_state_in_7_2_3,
  input      [0:0]    port_state_in_7_2_4,
  input      [0:0]    port_state_in_7_2_5,
  input      [0:0]    port_state_in_7_2_6,
  input      [0:0]    port_state_in_7_2_7,
  input      [0:0]    port_state_in_7_3_0,
  input      [0:0]    port_state_in_7_3_1,
  input      [0:0]    port_state_in_7_3_2,
  input      [0:0]    port_state_in_7_3_3,
  input      [0:0]    port_state_in_7_3_4,
  input      [0:0]    port_state_in_7_3_5,
  input      [0:0]    port_state_in_7_3_6,
  input      [0:0]    port_state_in_7_3_7,
  input      [0:0]    port_state_in_8_0_0,
  input      [0:0]    port_state_in_8_0_1,
  input      [0:0]    port_state_in_8_0_2,
  input      [0:0]    port_state_in_8_0_3,
  input      [0:0]    port_state_in_8_0_4,
  input      [0:0]    port_state_in_8_0_5,
  input      [0:0]    port_state_in_8_0_6,
  input      [0:0]    port_state_in_8_0_7,
  input      [0:0]    port_state_in_8_1_0,
  input      [0:0]    port_state_in_8_1_1,
  input      [0:0]    port_state_in_8_1_2,
  input      [0:0]    port_state_in_8_1_3,
  input      [0:0]    port_state_in_8_1_4,
  input      [0:0]    port_state_in_8_1_5,
  input      [0:0]    port_state_in_8_1_6,
  input      [0:0]    port_state_in_8_1_7,
  input      [0:0]    port_state_in_8_2_0,
  input      [0:0]    port_state_in_8_2_1,
  input      [0:0]    port_state_in_8_2_2,
  input      [0:0]    port_state_in_8_2_3,
  input      [0:0]    port_state_in_8_2_4,
  input      [0:0]    port_state_in_8_2_5,
  input      [0:0]    port_state_in_8_2_6,
  input      [0:0]    port_state_in_8_2_7,
  input      [0:0]    port_state_in_8_3_0,
  input      [0:0]    port_state_in_8_3_1,
  input      [0:0]    port_state_in_8_3_2,
  input      [0:0]    port_state_in_8_3_3,
  input      [0:0]    port_state_in_8_3_4,
  input      [0:0]    port_state_in_8_3_5,
  input      [0:0]    port_state_in_8_3_6,
  input      [0:0]    port_state_in_8_3_7,
  input      [0:0]    port_state_in_9_0_0,
  input      [0:0]    port_state_in_9_0_1,
  input      [0:0]    port_state_in_9_0_2,
  input      [0:0]    port_state_in_9_0_3,
  input      [0:0]    port_state_in_9_0_4,
  input      [0:0]    port_state_in_9_0_5,
  input      [0:0]    port_state_in_9_0_6,
  input      [0:0]    port_state_in_9_0_7,
  input      [0:0]    port_state_in_9_1_0,
  input      [0:0]    port_state_in_9_1_1,
  input      [0:0]    port_state_in_9_1_2,
  input      [0:0]    port_state_in_9_1_3,
  input      [0:0]    port_state_in_9_1_4,
  input      [0:0]    port_state_in_9_1_5,
  input      [0:0]    port_state_in_9_1_6,
  input      [0:0]    port_state_in_9_1_7,
  input      [0:0]    port_state_in_9_2_0,
  input      [0:0]    port_state_in_9_2_1,
  input      [0:0]    port_state_in_9_2_2,
  input      [0:0]    port_state_in_9_2_3,
  input      [0:0]    port_state_in_9_2_4,
  input      [0:0]    port_state_in_9_2_5,
  input      [0:0]    port_state_in_9_2_6,
  input      [0:0]    port_state_in_9_2_7,
  input      [0:0]    port_state_in_9_3_0,
  input      [0:0]    port_state_in_9_3_1,
  input      [0:0]    port_state_in_9_3_2,
  input      [0:0]    port_state_in_9_3_3,
  input      [0:0]    port_state_in_9_3_4,
  input      [0:0]    port_state_in_9_3_5,
  input      [0:0]    port_state_in_9_3_6,
  input      [0:0]    port_state_in_9_3_7,
  input      [0:0]    port_state_in_10_0_0,
  input      [0:0]    port_state_in_10_0_1,
  input      [0:0]    port_state_in_10_0_2,
  input      [0:0]    port_state_in_10_0_3,
  input      [0:0]    port_state_in_10_0_4,
  input      [0:0]    port_state_in_10_0_5,
  input      [0:0]    port_state_in_10_0_6,
  input      [0:0]    port_state_in_10_0_7,
  input      [0:0]    port_state_in_10_1_0,
  input      [0:0]    port_state_in_10_1_1,
  input      [0:0]    port_state_in_10_1_2,
  input      [0:0]    port_state_in_10_1_3,
  input      [0:0]    port_state_in_10_1_4,
  input      [0:0]    port_state_in_10_1_5,
  input      [0:0]    port_state_in_10_1_6,
  input      [0:0]    port_state_in_10_1_7,
  input      [0:0]    port_state_in_10_2_0,
  input      [0:0]    port_state_in_10_2_1,
  input      [0:0]    port_state_in_10_2_2,
  input      [0:0]    port_state_in_10_2_3,
  input      [0:0]    port_state_in_10_2_4,
  input      [0:0]    port_state_in_10_2_5,
  input      [0:0]    port_state_in_10_2_6,
  input      [0:0]    port_state_in_10_2_7,
  input      [0:0]    port_state_in_10_3_0,
  input      [0:0]    port_state_in_10_3_1,
  input      [0:0]    port_state_in_10_3_2,
  input      [0:0]    port_state_in_10_3_3,
  input      [0:0]    port_state_in_10_3_4,
  input      [0:0]    port_state_in_10_3_5,
  input      [0:0]    port_state_in_10_3_6,
  input      [0:0]    port_state_in_10_3_7,
  input      [0:0]    port_state_in_11_0_0,
  input      [0:0]    port_state_in_11_0_1,
  input      [0:0]    port_state_in_11_0_2,
  input      [0:0]    port_state_in_11_0_3,
  input      [0:0]    port_state_in_11_0_4,
  input      [0:0]    port_state_in_11_0_5,
  input      [0:0]    port_state_in_11_0_6,
  input      [0:0]    port_state_in_11_0_7,
  input      [0:0]    port_state_in_11_1_0,
  input      [0:0]    port_state_in_11_1_1,
  input      [0:0]    port_state_in_11_1_2,
  input      [0:0]    port_state_in_11_1_3,
  input      [0:0]    port_state_in_11_1_4,
  input      [0:0]    port_state_in_11_1_5,
  input      [0:0]    port_state_in_11_1_6,
  input      [0:0]    port_state_in_11_1_7,
  input      [0:0]    port_state_in_11_2_0,
  input      [0:0]    port_state_in_11_2_1,
  input      [0:0]    port_state_in_11_2_2,
  input      [0:0]    port_state_in_11_2_3,
  input      [0:0]    port_state_in_11_2_4,
  input      [0:0]    port_state_in_11_2_5,
  input      [0:0]    port_state_in_11_2_6,
  input      [0:0]    port_state_in_11_2_7,
  input      [0:0]    port_state_in_11_3_0,
  input      [0:0]    port_state_in_11_3_1,
  input      [0:0]    port_state_in_11_3_2,
  input      [0:0]    port_state_in_11_3_3,
  input      [0:0]    port_state_in_11_3_4,
  input      [0:0]    port_state_in_11_3_5,
  input      [0:0]    port_state_in_11_3_6,
  input      [0:0]    port_state_in_11_3_7,
  input      [0:0]    port_state_in_12_0_0,
  input      [0:0]    port_state_in_12_0_1,
  input      [0:0]    port_state_in_12_0_2,
  input      [0:0]    port_state_in_12_0_3,
  input      [0:0]    port_state_in_12_0_4,
  input      [0:0]    port_state_in_12_0_5,
  input      [0:0]    port_state_in_12_0_6,
  input      [0:0]    port_state_in_12_0_7,
  input      [0:0]    port_state_in_12_1_0,
  input      [0:0]    port_state_in_12_1_1,
  input      [0:0]    port_state_in_12_1_2,
  input      [0:0]    port_state_in_12_1_3,
  input      [0:0]    port_state_in_12_1_4,
  input      [0:0]    port_state_in_12_1_5,
  input      [0:0]    port_state_in_12_1_6,
  input      [0:0]    port_state_in_12_1_7,
  input      [0:0]    port_state_in_12_2_0,
  input      [0:0]    port_state_in_12_2_1,
  input      [0:0]    port_state_in_12_2_2,
  input      [0:0]    port_state_in_12_2_3,
  input      [0:0]    port_state_in_12_2_4,
  input      [0:0]    port_state_in_12_2_5,
  input      [0:0]    port_state_in_12_2_6,
  input      [0:0]    port_state_in_12_2_7,
  input      [0:0]    port_state_in_12_3_0,
  input      [0:0]    port_state_in_12_3_1,
  input      [0:0]    port_state_in_12_3_2,
  input      [0:0]    port_state_in_12_3_3,
  input      [0:0]    port_state_in_12_3_4,
  input      [0:0]    port_state_in_12_3_5,
  input      [0:0]    port_state_in_12_3_6,
  input      [0:0]    port_state_in_12_3_7,
  input      [0:0]    port_state_in_13_0_0,
  input      [0:0]    port_state_in_13_0_1,
  input      [0:0]    port_state_in_13_0_2,
  input      [0:0]    port_state_in_13_0_3,
  input      [0:0]    port_state_in_13_0_4,
  input      [0:0]    port_state_in_13_0_5,
  input      [0:0]    port_state_in_13_0_6,
  input      [0:0]    port_state_in_13_0_7,
  input      [0:0]    port_state_in_13_1_0,
  input      [0:0]    port_state_in_13_1_1,
  input      [0:0]    port_state_in_13_1_2,
  input      [0:0]    port_state_in_13_1_3,
  input      [0:0]    port_state_in_13_1_4,
  input      [0:0]    port_state_in_13_1_5,
  input      [0:0]    port_state_in_13_1_6,
  input      [0:0]    port_state_in_13_1_7,
  input      [0:0]    port_state_in_13_2_0,
  input      [0:0]    port_state_in_13_2_1,
  input      [0:0]    port_state_in_13_2_2,
  input      [0:0]    port_state_in_13_2_3,
  input      [0:0]    port_state_in_13_2_4,
  input      [0:0]    port_state_in_13_2_5,
  input      [0:0]    port_state_in_13_2_6,
  input      [0:0]    port_state_in_13_2_7,
  input      [0:0]    port_state_in_13_3_0,
  input      [0:0]    port_state_in_13_3_1,
  input      [0:0]    port_state_in_13_3_2,
  input      [0:0]    port_state_in_13_3_3,
  input      [0:0]    port_state_in_13_3_4,
  input      [0:0]    port_state_in_13_3_5,
  input      [0:0]    port_state_in_13_3_6,
  input      [0:0]    port_state_in_13_3_7,
  input      [0:0]    port_state_in_14_0_0,
  input      [0:0]    port_state_in_14_0_1,
  input      [0:0]    port_state_in_14_0_2,
  input      [0:0]    port_state_in_14_0_3,
  input      [0:0]    port_state_in_14_0_4,
  input      [0:0]    port_state_in_14_0_5,
  input      [0:0]    port_state_in_14_0_6,
  input      [0:0]    port_state_in_14_0_7,
  input      [0:0]    port_state_in_14_1_0,
  input      [0:0]    port_state_in_14_1_1,
  input      [0:0]    port_state_in_14_1_2,
  input      [0:0]    port_state_in_14_1_3,
  input      [0:0]    port_state_in_14_1_4,
  input      [0:0]    port_state_in_14_1_5,
  input      [0:0]    port_state_in_14_1_6,
  input      [0:0]    port_state_in_14_1_7,
  input      [0:0]    port_state_in_14_2_0,
  input      [0:0]    port_state_in_14_2_1,
  input      [0:0]    port_state_in_14_2_2,
  input      [0:0]    port_state_in_14_2_3,
  input      [0:0]    port_state_in_14_2_4,
  input      [0:0]    port_state_in_14_2_5,
  input      [0:0]    port_state_in_14_2_6,
  input      [0:0]    port_state_in_14_2_7,
  input      [0:0]    port_state_in_14_3_0,
  input      [0:0]    port_state_in_14_3_1,
  input      [0:0]    port_state_in_14_3_2,
  input      [0:0]    port_state_in_14_3_3,
  input      [0:0]    port_state_in_14_3_4,
  input      [0:0]    port_state_in_14_3_5,
  input      [0:0]    port_state_in_14_3_6,
  input      [0:0]    port_state_in_14_3_7,
  input      [0:0]    port_state_in_15_0_0,
  input      [0:0]    port_state_in_15_0_1,
  input      [0:0]    port_state_in_15_0_2,
  input      [0:0]    port_state_in_15_0_3,
  input      [0:0]    port_state_in_15_0_4,
  input      [0:0]    port_state_in_15_0_5,
  input      [0:0]    port_state_in_15_0_6,
  input      [0:0]    port_state_in_15_0_7,
  input      [0:0]    port_state_in_15_1_0,
  input      [0:0]    port_state_in_15_1_1,
  input      [0:0]    port_state_in_15_1_2,
  input      [0:0]    port_state_in_15_1_3,
  input      [0:0]    port_state_in_15_1_4,
  input      [0:0]    port_state_in_15_1_5,
  input      [0:0]    port_state_in_15_1_6,
  input      [0:0]    port_state_in_15_1_7,
  input      [0:0]    port_state_in_15_2_0,
  input      [0:0]    port_state_in_15_2_1,
  input      [0:0]    port_state_in_15_2_2,
  input      [0:0]    port_state_in_15_2_3,
  input      [0:0]    port_state_in_15_2_4,
  input      [0:0]    port_state_in_15_2_5,
  input      [0:0]    port_state_in_15_2_6,
  input      [0:0]    port_state_in_15_2_7,
  input      [0:0]    port_state_in_15_3_0,
  input      [0:0]    port_state_in_15_3_1,
  input      [0:0]    port_state_in_15_3_2,
  input      [0:0]    port_state_in_15_3_3,
  input      [0:0]    port_state_in_15_3_4,
  input      [0:0]    port_state_in_15_3_5,
  input      [0:0]    port_state_in_15_3_6,
  input      [0:0]    port_state_in_15_3_7,
  input      [0:0]    port_key_0_0_0,
  input      [0:0]    port_key_0_0_1,
  input      [0:0]    port_key_0_0_2,
  input      [0:0]    port_key_0_0_3,
  input      [0:0]    port_key_0_0_4,
  input      [0:0]    port_key_0_0_5,
  input      [0:0]    port_key_0_0_6,
  input      [0:0]    port_key_0_0_7,
  input      [0:0]    port_key_0_1_0,
  input      [0:0]    port_key_0_1_1,
  input      [0:0]    port_key_0_1_2,
  input      [0:0]    port_key_0_1_3,
  input      [0:0]    port_key_0_1_4,
  input      [0:0]    port_key_0_1_5,
  input      [0:0]    port_key_0_1_6,
  input      [0:0]    port_key_0_1_7,
  input      [0:0]    port_key_0_2_0,
  input      [0:0]    port_key_0_2_1,
  input      [0:0]    port_key_0_2_2,
  input      [0:0]    port_key_0_2_3,
  input      [0:0]    port_key_0_2_4,
  input      [0:0]    port_key_0_2_5,
  input      [0:0]    port_key_0_2_6,
  input      [0:0]    port_key_0_2_7,
  input      [0:0]    port_key_0_3_0,
  input      [0:0]    port_key_0_3_1,
  input      [0:0]    port_key_0_3_2,
  input      [0:0]    port_key_0_3_3,
  input      [0:0]    port_key_0_3_4,
  input      [0:0]    port_key_0_3_5,
  input      [0:0]    port_key_0_3_6,
  input      [0:0]    port_key_0_3_7,
  input      [0:0]    port_key_1_0_0,
  input      [0:0]    port_key_1_0_1,
  input      [0:0]    port_key_1_0_2,
  input      [0:0]    port_key_1_0_3,
  input      [0:0]    port_key_1_0_4,
  input      [0:0]    port_key_1_0_5,
  input      [0:0]    port_key_1_0_6,
  input      [0:0]    port_key_1_0_7,
  input      [0:0]    port_key_1_1_0,
  input      [0:0]    port_key_1_1_1,
  input      [0:0]    port_key_1_1_2,
  input      [0:0]    port_key_1_1_3,
  input      [0:0]    port_key_1_1_4,
  input      [0:0]    port_key_1_1_5,
  input      [0:0]    port_key_1_1_6,
  input      [0:0]    port_key_1_1_7,
  input      [0:0]    port_key_1_2_0,
  input      [0:0]    port_key_1_2_1,
  input      [0:0]    port_key_1_2_2,
  input      [0:0]    port_key_1_2_3,
  input      [0:0]    port_key_1_2_4,
  input      [0:0]    port_key_1_2_5,
  input      [0:0]    port_key_1_2_6,
  input      [0:0]    port_key_1_2_7,
  input      [0:0]    port_key_1_3_0,
  input      [0:0]    port_key_1_3_1,
  input      [0:0]    port_key_1_3_2,
  input      [0:0]    port_key_1_3_3,
  input      [0:0]    port_key_1_3_4,
  input      [0:0]    port_key_1_3_5,
  input      [0:0]    port_key_1_3_6,
  input      [0:0]    port_key_1_3_7,
  input      [0:0]    port_key_2_0_0,
  input      [0:0]    port_key_2_0_1,
  input      [0:0]    port_key_2_0_2,
  input      [0:0]    port_key_2_0_3,
  input      [0:0]    port_key_2_0_4,
  input      [0:0]    port_key_2_0_5,
  input      [0:0]    port_key_2_0_6,
  input      [0:0]    port_key_2_0_7,
  input      [0:0]    port_key_2_1_0,
  input      [0:0]    port_key_2_1_1,
  input      [0:0]    port_key_2_1_2,
  input      [0:0]    port_key_2_1_3,
  input      [0:0]    port_key_2_1_4,
  input      [0:0]    port_key_2_1_5,
  input      [0:0]    port_key_2_1_6,
  input      [0:0]    port_key_2_1_7,
  input      [0:0]    port_key_2_2_0,
  input      [0:0]    port_key_2_2_1,
  input      [0:0]    port_key_2_2_2,
  input      [0:0]    port_key_2_2_3,
  input      [0:0]    port_key_2_2_4,
  input      [0:0]    port_key_2_2_5,
  input      [0:0]    port_key_2_2_6,
  input      [0:0]    port_key_2_2_7,
  input      [0:0]    port_key_2_3_0,
  input      [0:0]    port_key_2_3_1,
  input      [0:0]    port_key_2_3_2,
  input      [0:0]    port_key_2_3_3,
  input      [0:0]    port_key_2_3_4,
  input      [0:0]    port_key_2_3_5,
  input      [0:0]    port_key_2_3_6,
  input      [0:0]    port_key_2_3_7,
  input      [0:0]    port_key_3_0_0,
  input      [0:0]    port_key_3_0_1,
  input      [0:0]    port_key_3_0_2,
  input      [0:0]    port_key_3_0_3,
  input      [0:0]    port_key_3_0_4,
  input      [0:0]    port_key_3_0_5,
  input      [0:0]    port_key_3_0_6,
  input      [0:0]    port_key_3_0_7,
  input      [0:0]    port_key_3_1_0,
  input      [0:0]    port_key_3_1_1,
  input      [0:0]    port_key_3_1_2,
  input      [0:0]    port_key_3_1_3,
  input      [0:0]    port_key_3_1_4,
  input      [0:0]    port_key_3_1_5,
  input      [0:0]    port_key_3_1_6,
  input      [0:0]    port_key_3_1_7,
  input      [0:0]    port_key_3_2_0,
  input      [0:0]    port_key_3_2_1,
  input      [0:0]    port_key_3_2_2,
  input      [0:0]    port_key_3_2_3,
  input      [0:0]    port_key_3_2_4,
  input      [0:0]    port_key_3_2_5,
  input      [0:0]    port_key_3_2_6,
  input      [0:0]    port_key_3_2_7,
  input      [0:0]    port_key_3_3_0,
  input      [0:0]    port_key_3_3_1,
  input      [0:0]    port_key_3_3_2,
  input      [0:0]    port_key_3_3_3,
  input      [0:0]    port_key_3_3_4,
  input      [0:0]    port_key_3_3_5,
  input      [0:0]    port_key_3_3_6,
  input      [0:0]    port_key_3_3_7,
  input      [0:0]    port_key_4_0_0,
  input      [0:0]    port_key_4_0_1,
  input      [0:0]    port_key_4_0_2,
  input      [0:0]    port_key_4_0_3,
  input      [0:0]    port_key_4_0_4,
  input      [0:0]    port_key_4_0_5,
  input      [0:0]    port_key_4_0_6,
  input      [0:0]    port_key_4_0_7,
  input      [0:0]    port_key_4_1_0,
  input      [0:0]    port_key_4_1_1,
  input      [0:0]    port_key_4_1_2,
  input      [0:0]    port_key_4_1_3,
  input      [0:0]    port_key_4_1_4,
  input      [0:0]    port_key_4_1_5,
  input      [0:0]    port_key_4_1_6,
  input      [0:0]    port_key_4_1_7,
  input      [0:0]    port_key_4_2_0,
  input      [0:0]    port_key_4_2_1,
  input      [0:0]    port_key_4_2_2,
  input      [0:0]    port_key_4_2_3,
  input      [0:0]    port_key_4_2_4,
  input      [0:0]    port_key_4_2_5,
  input      [0:0]    port_key_4_2_6,
  input      [0:0]    port_key_4_2_7,
  input      [0:0]    port_key_4_3_0,
  input      [0:0]    port_key_4_3_1,
  input      [0:0]    port_key_4_3_2,
  input      [0:0]    port_key_4_3_3,
  input      [0:0]    port_key_4_3_4,
  input      [0:0]    port_key_4_3_5,
  input      [0:0]    port_key_4_3_6,
  input      [0:0]    port_key_4_3_7,
  input      [0:0]    port_key_5_0_0,
  input      [0:0]    port_key_5_0_1,
  input      [0:0]    port_key_5_0_2,
  input      [0:0]    port_key_5_0_3,
  input      [0:0]    port_key_5_0_4,
  input      [0:0]    port_key_5_0_5,
  input      [0:0]    port_key_5_0_6,
  input      [0:0]    port_key_5_0_7,
  input      [0:0]    port_key_5_1_0,
  input      [0:0]    port_key_5_1_1,
  input      [0:0]    port_key_5_1_2,
  input      [0:0]    port_key_5_1_3,
  input      [0:0]    port_key_5_1_4,
  input      [0:0]    port_key_5_1_5,
  input      [0:0]    port_key_5_1_6,
  input      [0:0]    port_key_5_1_7,
  input      [0:0]    port_key_5_2_0,
  input      [0:0]    port_key_5_2_1,
  input      [0:0]    port_key_5_2_2,
  input      [0:0]    port_key_5_2_3,
  input      [0:0]    port_key_5_2_4,
  input      [0:0]    port_key_5_2_5,
  input      [0:0]    port_key_5_2_6,
  input      [0:0]    port_key_5_2_7,
  input      [0:0]    port_key_5_3_0,
  input      [0:0]    port_key_5_3_1,
  input      [0:0]    port_key_5_3_2,
  input      [0:0]    port_key_5_3_3,
  input      [0:0]    port_key_5_3_4,
  input      [0:0]    port_key_5_3_5,
  input      [0:0]    port_key_5_3_6,
  input      [0:0]    port_key_5_3_7,
  input      [0:0]    port_key_6_0_0,
  input      [0:0]    port_key_6_0_1,
  input      [0:0]    port_key_6_0_2,
  input      [0:0]    port_key_6_0_3,
  input      [0:0]    port_key_6_0_4,
  input      [0:0]    port_key_6_0_5,
  input      [0:0]    port_key_6_0_6,
  input      [0:0]    port_key_6_0_7,
  input      [0:0]    port_key_6_1_0,
  input      [0:0]    port_key_6_1_1,
  input      [0:0]    port_key_6_1_2,
  input      [0:0]    port_key_6_1_3,
  input      [0:0]    port_key_6_1_4,
  input      [0:0]    port_key_6_1_5,
  input      [0:0]    port_key_6_1_6,
  input      [0:0]    port_key_6_1_7,
  input      [0:0]    port_key_6_2_0,
  input      [0:0]    port_key_6_2_1,
  input      [0:0]    port_key_6_2_2,
  input      [0:0]    port_key_6_2_3,
  input      [0:0]    port_key_6_2_4,
  input      [0:0]    port_key_6_2_5,
  input      [0:0]    port_key_6_2_6,
  input      [0:0]    port_key_6_2_7,
  input      [0:0]    port_key_6_3_0,
  input      [0:0]    port_key_6_3_1,
  input      [0:0]    port_key_6_3_2,
  input      [0:0]    port_key_6_3_3,
  input      [0:0]    port_key_6_3_4,
  input      [0:0]    port_key_6_3_5,
  input      [0:0]    port_key_6_3_6,
  input      [0:0]    port_key_6_3_7,
  input      [0:0]    port_key_7_0_0,
  input      [0:0]    port_key_7_0_1,
  input      [0:0]    port_key_7_0_2,
  input      [0:0]    port_key_7_0_3,
  input      [0:0]    port_key_7_0_4,
  input      [0:0]    port_key_7_0_5,
  input      [0:0]    port_key_7_0_6,
  input      [0:0]    port_key_7_0_7,
  input      [0:0]    port_key_7_1_0,
  input      [0:0]    port_key_7_1_1,
  input      [0:0]    port_key_7_1_2,
  input      [0:0]    port_key_7_1_3,
  input      [0:0]    port_key_7_1_4,
  input      [0:0]    port_key_7_1_5,
  input      [0:0]    port_key_7_1_6,
  input      [0:0]    port_key_7_1_7,
  input      [0:0]    port_key_7_2_0,
  input      [0:0]    port_key_7_2_1,
  input      [0:0]    port_key_7_2_2,
  input      [0:0]    port_key_7_2_3,
  input      [0:0]    port_key_7_2_4,
  input      [0:0]    port_key_7_2_5,
  input      [0:0]    port_key_7_2_6,
  input      [0:0]    port_key_7_2_7,
  input      [0:0]    port_key_7_3_0,
  input      [0:0]    port_key_7_3_1,
  input      [0:0]    port_key_7_3_2,
  input      [0:0]    port_key_7_3_3,
  input      [0:0]    port_key_7_3_4,
  input      [0:0]    port_key_7_3_5,
  input      [0:0]    port_key_7_3_6,
  input      [0:0]    port_key_7_3_7,
  input      [0:0]    port_key_8_0_0,
  input      [0:0]    port_key_8_0_1,
  input      [0:0]    port_key_8_0_2,
  input      [0:0]    port_key_8_0_3,
  input      [0:0]    port_key_8_0_4,
  input      [0:0]    port_key_8_0_5,
  input      [0:0]    port_key_8_0_6,
  input      [0:0]    port_key_8_0_7,
  input      [0:0]    port_key_8_1_0,
  input      [0:0]    port_key_8_1_1,
  input      [0:0]    port_key_8_1_2,
  input      [0:0]    port_key_8_1_3,
  input      [0:0]    port_key_8_1_4,
  input      [0:0]    port_key_8_1_5,
  input      [0:0]    port_key_8_1_6,
  input      [0:0]    port_key_8_1_7,
  input      [0:0]    port_key_8_2_0,
  input      [0:0]    port_key_8_2_1,
  input      [0:0]    port_key_8_2_2,
  input      [0:0]    port_key_8_2_3,
  input      [0:0]    port_key_8_2_4,
  input      [0:0]    port_key_8_2_5,
  input      [0:0]    port_key_8_2_6,
  input      [0:0]    port_key_8_2_7,
  input      [0:0]    port_key_8_3_0,
  input      [0:0]    port_key_8_3_1,
  input      [0:0]    port_key_8_3_2,
  input      [0:0]    port_key_8_3_3,
  input      [0:0]    port_key_8_3_4,
  input      [0:0]    port_key_8_3_5,
  input      [0:0]    port_key_8_3_6,
  input      [0:0]    port_key_8_3_7,
  input      [0:0]    port_key_9_0_0,
  input      [0:0]    port_key_9_0_1,
  input      [0:0]    port_key_9_0_2,
  input      [0:0]    port_key_9_0_3,
  input      [0:0]    port_key_9_0_4,
  input      [0:0]    port_key_9_0_5,
  input      [0:0]    port_key_9_0_6,
  input      [0:0]    port_key_9_0_7,
  input      [0:0]    port_key_9_1_0,
  input      [0:0]    port_key_9_1_1,
  input      [0:0]    port_key_9_1_2,
  input      [0:0]    port_key_9_1_3,
  input      [0:0]    port_key_9_1_4,
  input      [0:0]    port_key_9_1_5,
  input      [0:0]    port_key_9_1_6,
  input      [0:0]    port_key_9_1_7,
  input      [0:0]    port_key_9_2_0,
  input      [0:0]    port_key_9_2_1,
  input      [0:0]    port_key_9_2_2,
  input      [0:0]    port_key_9_2_3,
  input      [0:0]    port_key_9_2_4,
  input      [0:0]    port_key_9_2_5,
  input      [0:0]    port_key_9_2_6,
  input      [0:0]    port_key_9_2_7,
  input      [0:0]    port_key_9_3_0,
  input      [0:0]    port_key_9_3_1,
  input      [0:0]    port_key_9_3_2,
  input      [0:0]    port_key_9_3_3,
  input      [0:0]    port_key_9_3_4,
  input      [0:0]    port_key_9_3_5,
  input      [0:0]    port_key_9_3_6,
  input      [0:0]    port_key_9_3_7,
  input      [0:0]    port_key_10_0_0,
  input      [0:0]    port_key_10_0_1,
  input      [0:0]    port_key_10_0_2,
  input      [0:0]    port_key_10_0_3,
  input      [0:0]    port_key_10_0_4,
  input      [0:0]    port_key_10_0_5,
  input      [0:0]    port_key_10_0_6,
  input      [0:0]    port_key_10_0_7,
  input      [0:0]    port_key_10_1_0,
  input      [0:0]    port_key_10_1_1,
  input      [0:0]    port_key_10_1_2,
  input      [0:0]    port_key_10_1_3,
  input      [0:0]    port_key_10_1_4,
  input      [0:0]    port_key_10_1_5,
  input      [0:0]    port_key_10_1_6,
  input      [0:0]    port_key_10_1_7,
  input      [0:0]    port_key_10_2_0,
  input      [0:0]    port_key_10_2_1,
  input      [0:0]    port_key_10_2_2,
  input      [0:0]    port_key_10_2_3,
  input      [0:0]    port_key_10_2_4,
  input      [0:0]    port_key_10_2_5,
  input      [0:0]    port_key_10_2_6,
  input      [0:0]    port_key_10_2_7,
  input      [0:0]    port_key_10_3_0,
  input      [0:0]    port_key_10_3_1,
  input      [0:0]    port_key_10_3_2,
  input      [0:0]    port_key_10_3_3,
  input      [0:0]    port_key_10_3_4,
  input      [0:0]    port_key_10_3_5,
  input      [0:0]    port_key_10_3_6,
  input      [0:0]    port_key_10_3_7,
  input      [0:0]    port_key_11_0_0,
  input      [0:0]    port_key_11_0_1,
  input      [0:0]    port_key_11_0_2,
  input      [0:0]    port_key_11_0_3,
  input      [0:0]    port_key_11_0_4,
  input      [0:0]    port_key_11_0_5,
  input      [0:0]    port_key_11_0_6,
  input      [0:0]    port_key_11_0_7,
  input      [0:0]    port_key_11_1_0,
  input      [0:0]    port_key_11_1_1,
  input      [0:0]    port_key_11_1_2,
  input      [0:0]    port_key_11_1_3,
  input      [0:0]    port_key_11_1_4,
  input      [0:0]    port_key_11_1_5,
  input      [0:0]    port_key_11_1_6,
  input      [0:0]    port_key_11_1_7,
  input      [0:0]    port_key_11_2_0,
  input      [0:0]    port_key_11_2_1,
  input      [0:0]    port_key_11_2_2,
  input      [0:0]    port_key_11_2_3,
  input      [0:0]    port_key_11_2_4,
  input      [0:0]    port_key_11_2_5,
  input      [0:0]    port_key_11_2_6,
  input      [0:0]    port_key_11_2_7,
  input      [0:0]    port_key_11_3_0,
  input      [0:0]    port_key_11_3_1,
  input      [0:0]    port_key_11_3_2,
  input      [0:0]    port_key_11_3_3,
  input      [0:0]    port_key_11_3_4,
  input      [0:0]    port_key_11_3_5,
  input      [0:0]    port_key_11_3_6,
  input      [0:0]    port_key_11_3_7,
  input      [0:0]    port_key_12_0_0,
  input      [0:0]    port_key_12_0_1,
  input      [0:0]    port_key_12_0_2,
  input      [0:0]    port_key_12_0_3,
  input      [0:0]    port_key_12_0_4,
  input      [0:0]    port_key_12_0_5,
  input      [0:0]    port_key_12_0_6,
  input      [0:0]    port_key_12_0_7,
  input      [0:0]    port_key_12_1_0,
  input      [0:0]    port_key_12_1_1,
  input      [0:0]    port_key_12_1_2,
  input      [0:0]    port_key_12_1_3,
  input      [0:0]    port_key_12_1_4,
  input      [0:0]    port_key_12_1_5,
  input      [0:0]    port_key_12_1_6,
  input      [0:0]    port_key_12_1_7,
  input      [0:0]    port_key_12_2_0,
  input      [0:0]    port_key_12_2_1,
  input      [0:0]    port_key_12_2_2,
  input      [0:0]    port_key_12_2_3,
  input      [0:0]    port_key_12_2_4,
  input      [0:0]    port_key_12_2_5,
  input      [0:0]    port_key_12_2_6,
  input      [0:0]    port_key_12_2_7,
  input      [0:0]    port_key_12_3_0,
  input      [0:0]    port_key_12_3_1,
  input      [0:0]    port_key_12_3_2,
  input      [0:0]    port_key_12_3_3,
  input      [0:0]    port_key_12_3_4,
  input      [0:0]    port_key_12_3_5,
  input      [0:0]    port_key_12_3_6,
  input      [0:0]    port_key_12_3_7,
  input      [0:0]    port_key_13_0_0,
  input      [0:0]    port_key_13_0_1,
  input      [0:0]    port_key_13_0_2,
  input      [0:0]    port_key_13_0_3,
  input      [0:0]    port_key_13_0_4,
  input      [0:0]    port_key_13_0_5,
  input      [0:0]    port_key_13_0_6,
  input      [0:0]    port_key_13_0_7,
  input      [0:0]    port_key_13_1_0,
  input      [0:0]    port_key_13_1_1,
  input      [0:0]    port_key_13_1_2,
  input      [0:0]    port_key_13_1_3,
  input      [0:0]    port_key_13_1_4,
  input      [0:0]    port_key_13_1_5,
  input      [0:0]    port_key_13_1_6,
  input      [0:0]    port_key_13_1_7,
  input      [0:0]    port_key_13_2_0,
  input      [0:0]    port_key_13_2_1,
  input      [0:0]    port_key_13_2_2,
  input      [0:0]    port_key_13_2_3,
  input      [0:0]    port_key_13_2_4,
  input      [0:0]    port_key_13_2_5,
  input      [0:0]    port_key_13_2_6,
  input      [0:0]    port_key_13_2_7,
  input      [0:0]    port_key_13_3_0,
  input      [0:0]    port_key_13_3_1,
  input      [0:0]    port_key_13_3_2,
  input      [0:0]    port_key_13_3_3,
  input      [0:0]    port_key_13_3_4,
  input      [0:0]    port_key_13_3_5,
  input      [0:0]    port_key_13_3_6,
  input      [0:0]    port_key_13_3_7,
  input      [0:0]    port_key_14_0_0,
  input      [0:0]    port_key_14_0_1,
  input      [0:0]    port_key_14_0_2,
  input      [0:0]    port_key_14_0_3,
  input      [0:0]    port_key_14_0_4,
  input      [0:0]    port_key_14_0_5,
  input      [0:0]    port_key_14_0_6,
  input      [0:0]    port_key_14_0_7,
  input      [0:0]    port_key_14_1_0,
  input      [0:0]    port_key_14_1_1,
  input      [0:0]    port_key_14_1_2,
  input      [0:0]    port_key_14_1_3,
  input      [0:0]    port_key_14_1_4,
  input      [0:0]    port_key_14_1_5,
  input      [0:0]    port_key_14_1_6,
  input      [0:0]    port_key_14_1_7,
  input      [0:0]    port_key_14_2_0,
  input      [0:0]    port_key_14_2_1,
  input      [0:0]    port_key_14_2_2,
  input      [0:0]    port_key_14_2_3,
  input      [0:0]    port_key_14_2_4,
  input      [0:0]    port_key_14_2_5,
  input      [0:0]    port_key_14_2_6,
  input      [0:0]    port_key_14_2_7,
  input      [0:0]    port_key_14_3_0,
  input      [0:0]    port_key_14_3_1,
  input      [0:0]    port_key_14_3_2,
  input      [0:0]    port_key_14_3_3,
  input      [0:0]    port_key_14_3_4,
  input      [0:0]    port_key_14_3_5,
  input      [0:0]    port_key_14_3_6,
  input      [0:0]    port_key_14_3_7,
  input      [0:0]    port_key_15_0_0,
  input      [0:0]    port_key_15_0_1,
  input      [0:0]    port_key_15_0_2,
  input      [0:0]    port_key_15_0_3,
  input      [0:0]    port_key_15_0_4,
  input      [0:0]    port_key_15_0_5,
  input      [0:0]    port_key_15_0_6,
  input      [0:0]    port_key_15_0_7,
  input      [0:0]    port_key_15_1_0,
  input      [0:0]    port_key_15_1_1,
  input      [0:0]    port_key_15_1_2,
  input      [0:0]    port_key_15_1_3,
  input      [0:0]    port_key_15_1_4,
  input      [0:0]    port_key_15_1_5,
  input      [0:0]    port_key_15_1_6,
  input      [0:0]    port_key_15_1_7,
  input      [0:0]    port_key_15_2_0,
  input      [0:0]    port_key_15_2_1,
  input      [0:0]    port_key_15_2_2,
  input      [0:0]    port_key_15_2_3,
  input      [0:0]    port_key_15_2_4,
  input      [0:0]    port_key_15_2_5,
  input      [0:0]    port_key_15_2_6,
  input      [0:0]    port_key_15_2_7,
  input      [0:0]    port_key_15_3_0,
  input      [0:0]    port_key_15_3_1,
  input      [0:0]    port_key_15_3_2,
  input      [0:0]    port_key_15_3_3,
  input      [0:0]    port_key_15_3_4,
  input      [0:0]    port_key_15_3_5,
  input      [0:0]    port_key_15_3_6,
  input      [0:0]    port_key_15_3_7,
  output     [0:0]    port_state_out_0_0_0,
  output     [0:0]    port_state_out_0_0_1,
  output     [0:0]    port_state_out_0_0_2,
  output     [0:0]    port_state_out_0_0_3,
  output     [0:0]    port_state_out_0_0_4,
  output     [0:0]    port_state_out_0_0_5,
  output     [0:0]    port_state_out_0_0_6,
  output     [0:0]    port_state_out_0_0_7,
  output     [0:0]    port_state_out_0_1_0,
  output     [0:0]    port_state_out_0_1_1,
  output     [0:0]    port_state_out_0_1_2,
  output     [0:0]    port_state_out_0_1_3,
  output     [0:0]    port_state_out_0_1_4,
  output     [0:0]    port_state_out_0_1_5,
  output     [0:0]    port_state_out_0_1_6,
  output     [0:0]    port_state_out_0_1_7,
  output     [0:0]    port_state_out_0_2_0,
  output     [0:0]    port_state_out_0_2_1,
  output     [0:0]    port_state_out_0_2_2,
  output     [0:0]    port_state_out_0_2_3,
  output     [0:0]    port_state_out_0_2_4,
  output     [0:0]    port_state_out_0_2_5,
  output     [0:0]    port_state_out_0_2_6,
  output     [0:0]    port_state_out_0_2_7,
  output     [0:0]    port_state_out_0_3_0,
  output     [0:0]    port_state_out_0_3_1,
  output     [0:0]    port_state_out_0_3_2,
  output     [0:0]    port_state_out_0_3_3,
  output     [0:0]    port_state_out_0_3_4,
  output     [0:0]    port_state_out_0_3_5,
  output     [0:0]    port_state_out_0_3_6,
  output     [0:0]    port_state_out_0_3_7,
  output     [0:0]    port_state_out_1_0_0,
  output     [0:0]    port_state_out_1_0_1,
  output     [0:0]    port_state_out_1_0_2,
  output     [0:0]    port_state_out_1_0_3,
  output     [0:0]    port_state_out_1_0_4,
  output     [0:0]    port_state_out_1_0_5,
  output     [0:0]    port_state_out_1_0_6,
  output     [0:0]    port_state_out_1_0_7,
  output     [0:0]    port_state_out_1_1_0,
  output     [0:0]    port_state_out_1_1_1,
  output     [0:0]    port_state_out_1_1_2,
  output     [0:0]    port_state_out_1_1_3,
  output     [0:0]    port_state_out_1_1_4,
  output     [0:0]    port_state_out_1_1_5,
  output     [0:0]    port_state_out_1_1_6,
  output     [0:0]    port_state_out_1_1_7,
  output     [0:0]    port_state_out_1_2_0,
  output     [0:0]    port_state_out_1_2_1,
  output     [0:0]    port_state_out_1_2_2,
  output     [0:0]    port_state_out_1_2_3,
  output     [0:0]    port_state_out_1_2_4,
  output     [0:0]    port_state_out_1_2_5,
  output     [0:0]    port_state_out_1_2_6,
  output     [0:0]    port_state_out_1_2_7,
  output     [0:0]    port_state_out_1_3_0,
  output     [0:0]    port_state_out_1_3_1,
  output     [0:0]    port_state_out_1_3_2,
  output     [0:0]    port_state_out_1_3_3,
  output     [0:0]    port_state_out_1_3_4,
  output     [0:0]    port_state_out_1_3_5,
  output     [0:0]    port_state_out_1_3_6,
  output     [0:0]    port_state_out_1_3_7,
  output     [0:0]    port_state_out_2_0_0,
  output     [0:0]    port_state_out_2_0_1,
  output     [0:0]    port_state_out_2_0_2,
  output     [0:0]    port_state_out_2_0_3,
  output     [0:0]    port_state_out_2_0_4,
  output     [0:0]    port_state_out_2_0_5,
  output     [0:0]    port_state_out_2_0_6,
  output     [0:0]    port_state_out_2_0_7,
  output     [0:0]    port_state_out_2_1_0,
  output     [0:0]    port_state_out_2_1_1,
  output     [0:0]    port_state_out_2_1_2,
  output     [0:0]    port_state_out_2_1_3,
  output     [0:0]    port_state_out_2_1_4,
  output     [0:0]    port_state_out_2_1_5,
  output     [0:0]    port_state_out_2_1_6,
  output     [0:0]    port_state_out_2_1_7,
  output     [0:0]    port_state_out_2_2_0,
  output     [0:0]    port_state_out_2_2_1,
  output     [0:0]    port_state_out_2_2_2,
  output     [0:0]    port_state_out_2_2_3,
  output     [0:0]    port_state_out_2_2_4,
  output     [0:0]    port_state_out_2_2_5,
  output     [0:0]    port_state_out_2_2_6,
  output     [0:0]    port_state_out_2_2_7,
  output     [0:0]    port_state_out_2_3_0,
  output     [0:0]    port_state_out_2_3_1,
  output     [0:0]    port_state_out_2_3_2,
  output     [0:0]    port_state_out_2_3_3,
  output     [0:0]    port_state_out_2_3_4,
  output     [0:0]    port_state_out_2_3_5,
  output     [0:0]    port_state_out_2_3_6,
  output     [0:0]    port_state_out_2_3_7,
  output     [0:0]    port_state_out_3_0_0,
  output     [0:0]    port_state_out_3_0_1,
  output     [0:0]    port_state_out_3_0_2,
  output     [0:0]    port_state_out_3_0_3,
  output     [0:0]    port_state_out_3_0_4,
  output     [0:0]    port_state_out_3_0_5,
  output     [0:0]    port_state_out_3_0_6,
  output     [0:0]    port_state_out_3_0_7,
  output     [0:0]    port_state_out_3_1_0,
  output     [0:0]    port_state_out_3_1_1,
  output     [0:0]    port_state_out_3_1_2,
  output     [0:0]    port_state_out_3_1_3,
  output     [0:0]    port_state_out_3_1_4,
  output     [0:0]    port_state_out_3_1_5,
  output     [0:0]    port_state_out_3_1_6,
  output     [0:0]    port_state_out_3_1_7,
  output     [0:0]    port_state_out_3_2_0,
  output     [0:0]    port_state_out_3_2_1,
  output     [0:0]    port_state_out_3_2_2,
  output     [0:0]    port_state_out_3_2_3,
  output     [0:0]    port_state_out_3_2_4,
  output     [0:0]    port_state_out_3_2_5,
  output     [0:0]    port_state_out_3_2_6,
  output     [0:0]    port_state_out_3_2_7,
  output     [0:0]    port_state_out_3_3_0,
  output     [0:0]    port_state_out_3_3_1,
  output     [0:0]    port_state_out_3_3_2,
  output     [0:0]    port_state_out_3_3_3,
  output     [0:0]    port_state_out_3_3_4,
  output     [0:0]    port_state_out_3_3_5,
  output     [0:0]    port_state_out_3_3_6,
  output     [0:0]    port_state_out_3_3_7,
  output     [0:0]    port_state_out_4_0_0,
  output     [0:0]    port_state_out_4_0_1,
  output     [0:0]    port_state_out_4_0_2,
  output     [0:0]    port_state_out_4_0_3,
  output     [0:0]    port_state_out_4_0_4,
  output     [0:0]    port_state_out_4_0_5,
  output     [0:0]    port_state_out_4_0_6,
  output     [0:0]    port_state_out_4_0_7,
  output     [0:0]    port_state_out_4_1_0,
  output     [0:0]    port_state_out_4_1_1,
  output     [0:0]    port_state_out_4_1_2,
  output     [0:0]    port_state_out_4_1_3,
  output     [0:0]    port_state_out_4_1_4,
  output     [0:0]    port_state_out_4_1_5,
  output     [0:0]    port_state_out_4_1_6,
  output     [0:0]    port_state_out_4_1_7,
  output     [0:0]    port_state_out_4_2_0,
  output     [0:0]    port_state_out_4_2_1,
  output     [0:0]    port_state_out_4_2_2,
  output     [0:0]    port_state_out_4_2_3,
  output     [0:0]    port_state_out_4_2_4,
  output     [0:0]    port_state_out_4_2_5,
  output     [0:0]    port_state_out_4_2_6,
  output     [0:0]    port_state_out_4_2_7,
  output     [0:0]    port_state_out_4_3_0,
  output     [0:0]    port_state_out_4_3_1,
  output     [0:0]    port_state_out_4_3_2,
  output     [0:0]    port_state_out_4_3_3,
  output     [0:0]    port_state_out_4_3_4,
  output     [0:0]    port_state_out_4_3_5,
  output     [0:0]    port_state_out_4_3_6,
  output     [0:0]    port_state_out_4_3_7,
  output     [0:0]    port_state_out_5_0_0,
  output     [0:0]    port_state_out_5_0_1,
  output     [0:0]    port_state_out_5_0_2,
  output     [0:0]    port_state_out_5_0_3,
  output     [0:0]    port_state_out_5_0_4,
  output     [0:0]    port_state_out_5_0_5,
  output     [0:0]    port_state_out_5_0_6,
  output     [0:0]    port_state_out_5_0_7,
  output     [0:0]    port_state_out_5_1_0,
  output     [0:0]    port_state_out_5_1_1,
  output     [0:0]    port_state_out_5_1_2,
  output     [0:0]    port_state_out_5_1_3,
  output     [0:0]    port_state_out_5_1_4,
  output     [0:0]    port_state_out_5_1_5,
  output     [0:0]    port_state_out_5_1_6,
  output     [0:0]    port_state_out_5_1_7,
  output     [0:0]    port_state_out_5_2_0,
  output     [0:0]    port_state_out_5_2_1,
  output     [0:0]    port_state_out_5_2_2,
  output     [0:0]    port_state_out_5_2_3,
  output     [0:0]    port_state_out_5_2_4,
  output     [0:0]    port_state_out_5_2_5,
  output     [0:0]    port_state_out_5_2_6,
  output     [0:0]    port_state_out_5_2_7,
  output     [0:0]    port_state_out_5_3_0,
  output     [0:0]    port_state_out_5_3_1,
  output     [0:0]    port_state_out_5_3_2,
  output     [0:0]    port_state_out_5_3_3,
  output     [0:0]    port_state_out_5_3_4,
  output     [0:0]    port_state_out_5_3_5,
  output     [0:0]    port_state_out_5_3_6,
  output     [0:0]    port_state_out_5_3_7,
  output     [0:0]    port_state_out_6_0_0,
  output     [0:0]    port_state_out_6_0_1,
  output     [0:0]    port_state_out_6_0_2,
  output     [0:0]    port_state_out_6_0_3,
  output     [0:0]    port_state_out_6_0_4,
  output     [0:0]    port_state_out_6_0_5,
  output     [0:0]    port_state_out_6_0_6,
  output     [0:0]    port_state_out_6_0_7,
  output     [0:0]    port_state_out_6_1_0,
  output     [0:0]    port_state_out_6_1_1,
  output     [0:0]    port_state_out_6_1_2,
  output     [0:0]    port_state_out_6_1_3,
  output     [0:0]    port_state_out_6_1_4,
  output     [0:0]    port_state_out_6_1_5,
  output     [0:0]    port_state_out_6_1_6,
  output     [0:0]    port_state_out_6_1_7,
  output     [0:0]    port_state_out_6_2_0,
  output     [0:0]    port_state_out_6_2_1,
  output     [0:0]    port_state_out_6_2_2,
  output     [0:0]    port_state_out_6_2_3,
  output     [0:0]    port_state_out_6_2_4,
  output     [0:0]    port_state_out_6_2_5,
  output     [0:0]    port_state_out_6_2_6,
  output     [0:0]    port_state_out_6_2_7,
  output     [0:0]    port_state_out_6_3_0,
  output     [0:0]    port_state_out_6_3_1,
  output     [0:0]    port_state_out_6_3_2,
  output     [0:0]    port_state_out_6_3_3,
  output     [0:0]    port_state_out_6_3_4,
  output     [0:0]    port_state_out_6_3_5,
  output     [0:0]    port_state_out_6_3_6,
  output     [0:0]    port_state_out_6_3_7,
  output     [0:0]    port_state_out_7_0_0,
  output     [0:0]    port_state_out_7_0_1,
  output     [0:0]    port_state_out_7_0_2,
  output     [0:0]    port_state_out_7_0_3,
  output     [0:0]    port_state_out_7_0_4,
  output     [0:0]    port_state_out_7_0_5,
  output     [0:0]    port_state_out_7_0_6,
  output     [0:0]    port_state_out_7_0_7,
  output     [0:0]    port_state_out_7_1_0,
  output     [0:0]    port_state_out_7_1_1,
  output     [0:0]    port_state_out_7_1_2,
  output     [0:0]    port_state_out_7_1_3,
  output     [0:0]    port_state_out_7_1_4,
  output     [0:0]    port_state_out_7_1_5,
  output     [0:0]    port_state_out_7_1_6,
  output     [0:0]    port_state_out_7_1_7,
  output     [0:0]    port_state_out_7_2_0,
  output     [0:0]    port_state_out_7_2_1,
  output     [0:0]    port_state_out_7_2_2,
  output     [0:0]    port_state_out_7_2_3,
  output     [0:0]    port_state_out_7_2_4,
  output     [0:0]    port_state_out_7_2_5,
  output     [0:0]    port_state_out_7_2_6,
  output     [0:0]    port_state_out_7_2_7,
  output     [0:0]    port_state_out_7_3_0,
  output     [0:0]    port_state_out_7_3_1,
  output     [0:0]    port_state_out_7_3_2,
  output     [0:0]    port_state_out_7_3_3,
  output     [0:0]    port_state_out_7_3_4,
  output     [0:0]    port_state_out_7_3_5,
  output     [0:0]    port_state_out_7_3_6,
  output     [0:0]    port_state_out_7_3_7,
  output     [0:0]    port_state_out_8_0_0,
  output     [0:0]    port_state_out_8_0_1,
  output     [0:0]    port_state_out_8_0_2,
  output     [0:0]    port_state_out_8_0_3,
  output     [0:0]    port_state_out_8_0_4,
  output     [0:0]    port_state_out_8_0_5,
  output     [0:0]    port_state_out_8_0_6,
  output     [0:0]    port_state_out_8_0_7,
  output     [0:0]    port_state_out_8_1_0,
  output     [0:0]    port_state_out_8_1_1,
  output     [0:0]    port_state_out_8_1_2,
  output     [0:0]    port_state_out_8_1_3,
  output     [0:0]    port_state_out_8_1_4,
  output     [0:0]    port_state_out_8_1_5,
  output     [0:0]    port_state_out_8_1_6,
  output     [0:0]    port_state_out_8_1_7,
  output     [0:0]    port_state_out_8_2_0,
  output     [0:0]    port_state_out_8_2_1,
  output     [0:0]    port_state_out_8_2_2,
  output     [0:0]    port_state_out_8_2_3,
  output     [0:0]    port_state_out_8_2_4,
  output     [0:0]    port_state_out_8_2_5,
  output     [0:0]    port_state_out_8_2_6,
  output     [0:0]    port_state_out_8_2_7,
  output     [0:0]    port_state_out_8_3_0,
  output     [0:0]    port_state_out_8_3_1,
  output     [0:0]    port_state_out_8_3_2,
  output     [0:0]    port_state_out_8_3_3,
  output     [0:0]    port_state_out_8_3_4,
  output     [0:0]    port_state_out_8_3_5,
  output     [0:0]    port_state_out_8_3_6,
  output     [0:0]    port_state_out_8_3_7,
  output     [0:0]    port_state_out_9_0_0,
  output     [0:0]    port_state_out_9_0_1,
  output     [0:0]    port_state_out_9_0_2,
  output     [0:0]    port_state_out_9_0_3,
  output     [0:0]    port_state_out_9_0_4,
  output     [0:0]    port_state_out_9_0_5,
  output     [0:0]    port_state_out_9_0_6,
  output     [0:0]    port_state_out_9_0_7,
  output     [0:0]    port_state_out_9_1_0,
  output     [0:0]    port_state_out_9_1_1,
  output     [0:0]    port_state_out_9_1_2,
  output     [0:0]    port_state_out_9_1_3,
  output     [0:0]    port_state_out_9_1_4,
  output     [0:0]    port_state_out_9_1_5,
  output     [0:0]    port_state_out_9_1_6,
  output     [0:0]    port_state_out_9_1_7,
  output     [0:0]    port_state_out_9_2_0,
  output     [0:0]    port_state_out_9_2_1,
  output     [0:0]    port_state_out_9_2_2,
  output     [0:0]    port_state_out_9_2_3,
  output     [0:0]    port_state_out_9_2_4,
  output     [0:0]    port_state_out_9_2_5,
  output     [0:0]    port_state_out_9_2_6,
  output     [0:0]    port_state_out_9_2_7,
  output     [0:0]    port_state_out_9_3_0,
  output     [0:0]    port_state_out_9_3_1,
  output     [0:0]    port_state_out_9_3_2,
  output     [0:0]    port_state_out_9_3_3,
  output     [0:0]    port_state_out_9_3_4,
  output     [0:0]    port_state_out_9_3_5,
  output     [0:0]    port_state_out_9_3_6,
  output     [0:0]    port_state_out_9_3_7,
  output     [0:0]    port_state_out_10_0_0,
  output     [0:0]    port_state_out_10_0_1,
  output     [0:0]    port_state_out_10_0_2,
  output     [0:0]    port_state_out_10_0_3,
  output     [0:0]    port_state_out_10_0_4,
  output     [0:0]    port_state_out_10_0_5,
  output     [0:0]    port_state_out_10_0_6,
  output     [0:0]    port_state_out_10_0_7,
  output     [0:0]    port_state_out_10_1_0,
  output     [0:0]    port_state_out_10_1_1,
  output     [0:0]    port_state_out_10_1_2,
  output     [0:0]    port_state_out_10_1_3,
  output     [0:0]    port_state_out_10_1_4,
  output     [0:0]    port_state_out_10_1_5,
  output     [0:0]    port_state_out_10_1_6,
  output     [0:0]    port_state_out_10_1_7,
  output     [0:0]    port_state_out_10_2_0,
  output     [0:0]    port_state_out_10_2_1,
  output     [0:0]    port_state_out_10_2_2,
  output     [0:0]    port_state_out_10_2_3,
  output     [0:0]    port_state_out_10_2_4,
  output     [0:0]    port_state_out_10_2_5,
  output     [0:0]    port_state_out_10_2_6,
  output     [0:0]    port_state_out_10_2_7,
  output     [0:0]    port_state_out_10_3_0,
  output     [0:0]    port_state_out_10_3_1,
  output     [0:0]    port_state_out_10_3_2,
  output     [0:0]    port_state_out_10_3_3,
  output     [0:0]    port_state_out_10_3_4,
  output     [0:0]    port_state_out_10_3_5,
  output     [0:0]    port_state_out_10_3_6,
  output     [0:0]    port_state_out_10_3_7,
  output     [0:0]    port_state_out_11_0_0,
  output     [0:0]    port_state_out_11_0_1,
  output     [0:0]    port_state_out_11_0_2,
  output     [0:0]    port_state_out_11_0_3,
  output     [0:0]    port_state_out_11_0_4,
  output     [0:0]    port_state_out_11_0_5,
  output     [0:0]    port_state_out_11_0_6,
  output     [0:0]    port_state_out_11_0_7,
  output     [0:0]    port_state_out_11_1_0,
  output     [0:0]    port_state_out_11_1_1,
  output     [0:0]    port_state_out_11_1_2,
  output     [0:0]    port_state_out_11_1_3,
  output     [0:0]    port_state_out_11_1_4,
  output     [0:0]    port_state_out_11_1_5,
  output     [0:0]    port_state_out_11_1_6,
  output     [0:0]    port_state_out_11_1_7,
  output     [0:0]    port_state_out_11_2_0,
  output     [0:0]    port_state_out_11_2_1,
  output     [0:0]    port_state_out_11_2_2,
  output     [0:0]    port_state_out_11_2_3,
  output     [0:0]    port_state_out_11_2_4,
  output     [0:0]    port_state_out_11_2_5,
  output     [0:0]    port_state_out_11_2_6,
  output     [0:0]    port_state_out_11_2_7,
  output     [0:0]    port_state_out_11_3_0,
  output     [0:0]    port_state_out_11_3_1,
  output     [0:0]    port_state_out_11_3_2,
  output     [0:0]    port_state_out_11_3_3,
  output     [0:0]    port_state_out_11_3_4,
  output     [0:0]    port_state_out_11_3_5,
  output     [0:0]    port_state_out_11_3_6,
  output     [0:0]    port_state_out_11_3_7,
  output     [0:0]    port_state_out_12_0_0,
  output     [0:0]    port_state_out_12_0_1,
  output     [0:0]    port_state_out_12_0_2,
  output     [0:0]    port_state_out_12_0_3,
  output     [0:0]    port_state_out_12_0_4,
  output     [0:0]    port_state_out_12_0_5,
  output     [0:0]    port_state_out_12_0_6,
  output     [0:0]    port_state_out_12_0_7,
  output     [0:0]    port_state_out_12_1_0,
  output     [0:0]    port_state_out_12_1_1,
  output     [0:0]    port_state_out_12_1_2,
  output     [0:0]    port_state_out_12_1_3,
  output     [0:0]    port_state_out_12_1_4,
  output     [0:0]    port_state_out_12_1_5,
  output     [0:0]    port_state_out_12_1_6,
  output     [0:0]    port_state_out_12_1_7,
  output     [0:0]    port_state_out_12_2_0,
  output     [0:0]    port_state_out_12_2_1,
  output     [0:0]    port_state_out_12_2_2,
  output     [0:0]    port_state_out_12_2_3,
  output     [0:0]    port_state_out_12_2_4,
  output     [0:0]    port_state_out_12_2_5,
  output     [0:0]    port_state_out_12_2_6,
  output     [0:0]    port_state_out_12_2_7,
  output     [0:0]    port_state_out_12_3_0,
  output     [0:0]    port_state_out_12_3_1,
  output     [0:0]    port_state_out_12_3_2,
  output     [0:0]    port_state_out_12_3_3,
  output     [0:0]    port_state_out_12_3_4,
  output     [0:0]    port_state_out_12_3_5,
  output     [0:0]    port_state_out_12_3_6,
  output     [0:0]    port_state_out_12_3_7,
  output     [0:0]    port_state_out_13_0_0,
  output     [0:0]    port_state_out_13_0_1,
  output     [0:0]    port_state_out_13_0_2,
  output     [0:0]    port_state_out_13_0_3,
  output     [0:0]    port_state_out_13_0_4,
  output     [0:0]    port_state_out_13_0_5,
  output     [0:0]    port_state_out_13_0_6,
  output     [0:0]    port_state_out_13_0_7,
  output     [0:0]    port_state_out_13_1_0,
  output     [0:0]    port_state_out_13_1_1,
  output     [0:0]    port_state_out_13_1_2,
  output     [0:0]    port_state_out_13_1_3,
  output     [0:0]    port_state_out_13_1_4,
  output     [0:0]    port_state_out_13_1_5,
  output     [0:0]    port_state_out_13_1_6,
  output     [0:0]    port_state_out_13_1_7,
  output     [0:0]    port_state_out_13_2_0,
  output     [0:0]    port_state_out_13_2_1,
  output     [0:0]    port_state_out_13_2_2,
  output     [0:0]    port_state_out_13_2_3,
  output     [0:0]    port_state_out_13_2_4,
  output     [0:0]    port_state_out_13_2_5,
  output     [0:0]    port_state_out_13_2_6,
  output     [0:0]    port_state_out_13_2_7,
  output     [0:0]    port_state_out_13_3_0,
  output     [0:0]    port_state_out_13_3_1,
  output     [0:0]    port_state_out_13_3_2,
  output     [0:0]    port_state_out_13_3_3,
  output     [0:0]    port_state_out_13_3_4,
  output     [0:0]    port_state_out_13_3_5,
  output     [0:0]    port_state_out_13_3_6,
  output     [0:0]    port_state_out_13_3_7,
  output     [0:0]    port_state_out_14_0_0,
  output     [0:0]    port_state_out_14_0_1,
  output     [0:0]    port_state_out_14_0_2,
  output     [0:0]    port_state_out_14_0_3,
  output     [0:0]    port_state_out_14_0_4,
  output     [0:0]    port_state_out_14_0_5,
  output     [0:0]    port_state_out_14_0_6,
  output     [0:0]    port_state_out_14_0_7,
  output     [0:0]    port_state_out_14_1_0,
  output     [0:0]    port_state_out_14_1_1,
  output     [0:0]    port_state_out_14_1_2,
  output     [0:0]    port_state_out_14_1_3,
  output     [0:0]    port_state_out_14_1_4,
  output     [0:0]    port_state_out_14_1_5,
  output     [0:0]    port_state_out_14_1_6,
  output     [0:0]    port_state_out_14_1_7,
  output     [0:0]    port_state_out_14_2_0,
  output     [0:0]    port_state_out_14_2_1,
  output     [0:0]    port_state_out_14_2_2,
  output     [0:0]    port_state_out_14_2_3,
  output     [0:0]    port_state_out_14_2_4,
  output     [0:0]    port_state_out_14_2_5,
  output     [0:0]    port_state_out_14_2_6,
  output     [0:0]    port_state_out_14_2_7,
  output     [0:0]    port_state_out_14_3_0,
  output     [0:0]    port_state_out_14_3_1,
  output     [0:0]    port_state_out_14_3_2,
  output     [0:0]    port_state_out_14_3_3,
  output     [0:0]    port_state_out_14_3_4,
  output     [0:0]    port_state_out_14_3_5,
  output     [0:0]    port_state_out_14_3_6,
  output     [0:0]    port_state_out_14_3_7,
  output     [0:0]    port_state_out_15_0_0,
  output     [0:0]    port_state_out_15_0_1,
  output     [0:0]    port_state_out_15_0_2,
  output     [0:0]    port_state_out_15_0_3,
  output     [0:0]    port_state_out_15_0_4,
  output     [0:0]    port_state_out_15_0_5,
  output     [0:0]    port_state_out_15_0_6,
  output     [0:0]    port_state_out_15_0_7,
  output     [0:0]    port_state_out_15_1_0,
  output     [0:0]    port_state_out_15_1_1,
  output     [0:0]    port_state_out_15_1_2,
  output     [0:0]    port_state_out_15_1_3,
  output     [0:0]    port_state_out_15_1_4,
  output     [0:0]    port_state_out_15_1_5,
  output     [0:0]    port_state_out_15_1_6,
  output     [0:0]    port_state_out_15_1_7,
  output     [0:0]    port_state_out_15_2_0,
  output     [0:0]    port_state_out_15_2_1,
  output     [0:0]    port_state_out_15_2_2,
  output     [0:0]    port_state_out_15_2_3,
  output     [0:0]    port_state_out_15_2_4,
  output     [0:0]    port_state_out_15_2_5,
  output     [0:0]    port_state_out_15_2_6,
  output     [0:0]    port_state_out_15_2_7,
  output     [0:0]    port_state_out_15_3_0,
  output     [0:0]    port_state_out_15_3_1,
  output     [0:0]    port_state_out_15_3_2,
  output     [0:0]    port_state_out_15_3_3,
  output     [0:0]    port_state_out_15_3_4,
  output     [0:0]    port_state_out_15_3_5,
  output     [0:0]    port_state_out_15_3_6,
  output     [0:0]    port_state_out_15_3_7
);


  assign port_state_out_0_0_0 = (port_state_in_0_0_0 ^ port_key_0_0_0);
  assign port_state_out_0_0_1 = (port_state_in_0_0_1 ^ port_key_0_0_1);
  assign port_state_out_0_0_2 = (port_state_in_0_0_2 ^ port_key_0_0_2);
  assign port_state_out_0_0_3 = (port_state_in_0_0_3 ^ port_key_0_0_3);
  assign port_state_out_0_0_4 = (port_state_in_0_0_4 ^ port_key_0_0_4);
  assign port_state_out_0_0_5 = (port_state_in_0_0_5 ^ port_key_0_0_5);
  assign port_state_out_0_0_6 = (port_state_in_0_0_6 ^ port_key_0_0_6);
  assign port_state_out_0_0_7 = (port_state_in_0_0_7 ^ port_key_0_0_7);
  assign port_state_out_0_1_0 = (port_state_in_0_1_0 ^ port_key_0_1_0);
  assign port_state_out_0_1_1 = (port_state_in_0_1_1 ^ port_key_0_1_1);
  assign port_state_out_0_1_2 = (port_state_in_0_1_2 ^ port_key_0_1_2);
  assign port_state_out_0_1_3 = (port_state_in_0_1_3 ^ port_key_0_1_3);
  assign port_state_out_0_1_4 = (port_state_in_0_1_4 ^ port_key_0_1_4);
  assign port_state_out_0_1_5 = (port_state_in_0_1_5 ^ port_key_0_1_5);
  assign port_state_out_0_1_6 = (port_state_in_0_1_6 ^ port_key_0_1_6);
  assign port_state_out_0_1_7 = (port_state_in_0_1_7 ^ port_key_0_1_7);
  assign port_state_out_0_2_0 = (port_state_in_0_2_0 ^ port_key_0_2_0);
  assign port_state_out_0_2_1 = (port_state_in_0_2_1 ^ port_key_0_2_1);
  assign port_state_out_0_2_2 = (port_state_in_0_2_2 ^ port_key_0_2_2);
  assign port_state_out_0_2_3 = (port_state_in_0_2_3 ^ port_key_0_2_3);
  assign port_state_out_0_2_4 = (port_state_in_0_2_4 ^ port_key_0_2_4);
  assign port_state_out_0_2_5 = (port_state_in_0_2_5 ^ port_key_0_2_5);
  assign port_state_out_0_2_6 = (port_state_in_0_2_6 ^ port_key_0_2_6);
  assign port_state_out_0_2_7 = (port_state_in_0_2_7 ^ port_key_0_2_7);
  assign port_state_out_0_3_0 = (port_state_in_0_3_0 ^ port_key_0_3_0);
  assign port_state_out_0_3_1 = (port_state_in_0_3_1 ^ port_key_0_3_1);
  assign port_state_out_0_3_2 = (port_state_in_0_3_2 ^ port_key_0_3_2);
  assign port_state_out_0_3_3 = (port_state_in_0_3_3 ^ port_key_0_3_3);
  assign port_state_out_0_3_4 = (port_state_in_0_3_4 ^ port_key_0_3_4);
  assign port_state_out_0_3_5 = (port_state_in_0_3_5 ^ port_key_0_3_5);
  assign port_state_out_0_3_6 = (port_state_in_0_3_6 ^ port_key_0_3_6);
  assign port_state_out_0_3_7 = (port_state_in_0_3_7 ^ port_key_0_3_7);
  assign port_state_out_1_0_0 = (port_state_in_1_0_0 ^ port_key_1_0_0);
  assign port_state_out_1_0_1 = (port_state_in_1_0_1 ^ port_key_1_0_1);
  assign port_state_out_1_0_2 = (port_state_in_1_0_2 ^ port_key_1_0_2);
  assign port_state_out_1_0_3 = (port_state_in_1_0_3 ^ port_key_1_0_3);
  assign port_state_out_1_0_4 = (port_state_in_1_0_4 ^ port_key_1_0_4);
  assign port_state_out_1_0_5 = (port_state_in_1_0_5 ^ port_key_1_0_5);
  assign port_state_out_1_0_6 = (port_state_in_1_0_6 ^ port_key_1_0_6);
  assign port_state_out_1_0_7 = (port_state_in_1_0_7 ^ port_key_1_0_7);
  assign port_state_out_1_1_0 = (port_state_in_1_1_0 ^ port_key_1_1_0);
  assign port_state_out_1_1_1 = (port_state_in_1_1_1 ^ port_key_1_1_1);
  assign port_state_out_1_1_2 = (port_state_in_1_1_2 ^ port_key_1_1_2);
  assign port_state_out_1_1_3 = (port_state_in_1_1_3 ^ port_key_1_1_3);
  assign port_state_out_1_1_4 = (port_state_in_1_1_4 ^ port_key_1_1_4);
  assign port_state_out_1_1_5 = (port_state_in_1_1_5 ^ port_key_1_1_5);
  assign port_state_out_1_1_6 = (port_state_in_1_1_6 ^ port_key_1_1_6);
  assign port_state_out_1_1_7 = (port_state_in_1_1_7 ^ port_key_1_1_7);
  assign port_state_out_1_2_0 = (port_state_in_1_2_0 ^ port_key_1_2_0);
  assign port_state_out_1_2_1 = (port_state_in_1_2_1 ^ port_key_1_2_1);
  assign port_state_out_1_2_2 = (port_state_in_1_2_2 ^ port_key_1_2_2);
  assign port_state_out_1_2_3 = (port_state_in_1_2_3 ^ port_key_1_2_3);
  assign port_state_out_1_2_4 = (port_state_in_1_2_4 ^ port_key_1_2_4);
  assign port_state_out_1_2_5 = (port_state_in_1_2_5 ^ port_key_1_2_5);
  assign port_state_out_1_2_6 = (port_state_in_1_2_6 ^ port_key_1_2_6);
  assign port_state_out_1_2_7 = (port_state_in_1_2_7 ^ port_key_1_2_7);
  assign port_state_out_1_3_0 = (port_state_in_1_3_0 ^ port_key_1_3_0);
  assign port_state_out_1_3_1 = (port_state_in_1_3_1 ^ port_key_1_3_1);
  assign port_state_out_1_3_2 = (port_state_in_1_3_2 ^ port_key_1_3_2);
  assign port_state_out_1_3_3 = (port_state_in_1_3_3 ^ port_key_1_3_3);
  assign port_state_out_1_3_4 = (port_state_in_1_3_4 ^ port_key_1_3_4);
  assign port_state_out_1_3_5 = (port_state_in_1_3_5 ^ port_key_1_3_5);
  assign port_state_out_1_3_6 = (port_state_in_1_3_6 ^ port_key_1_3_6);
  assign port_state_out_1_3_7 = (port_state_in_1_3_7 ^ port_key_1_3_7);
  assign port_state_out_2_0_0 = (port_state_in_2_0_0 ^ port_key_2_0_0);
  assign port_state_out_2_0_1 = (port_state_in_2_0_1 ^ port_key_2_0_1);
  assign port_state_out_2_0_2 = (port_state_in_2_0_2 ^ port_key_2_0_2);
  assign port_state_out_2_0_3 = (port_state_in_2_0_3 ^ port_key_2_0_3);
  assign port_state_out_2_0_4 = (port_state_in_2_0_4 ^ port_key_2_0_4);
  assign port_state_out_2_0_5 = (port_state_in_2_0_5 ^ port_key_2_0_5);
  assign port_state_out_2_0_6 = (port_state_in_2_0_6 ^ port_key_2_0_6);
  assign port_state_out_2_0_7 = (port_state_in_2_0_7 ^ port_key_2_0_7);
  assign port_state_out_2_1_0 = (port_state_in_2_1_0 ^ port_key_2_1_0);
  assign port_state_out_2_1_1 = (port_state_in_2_1_1 ^ port_key_2_1_1);
  assign port_state_out_2_1_2 = (port_state_in_2_1_2 ^ port_key_2_1_2);
  assign port_state_out_2_1_3 = (port_state_in_2_1_3 ^ port_key_2_1_3);
  assign port_state_out_2_1_4 = (port_state_in_2_1_4 ^ port_key_2_1_4);
  assign port_state_out_2_1_5 = (port_state_in_2_1_5 ^ port_key_2_1_5);
  assign port_state_out_2_1_6 = (port_state_in_2_1_6 ^ port_key_2_1_6);
  assign port_state_out_2_1_7 = (port_state_in_2_1_7 ^ port_key_2_1_7);
  assign port_state_out_2_2_0 = (port_state_in_2_2_0 ^ port_key_2_2_0);
  assign port_state_out_2_2_1 = (port_state_in_2_2_1 ^ port_key_2_2_1);
  assign port_state_out_2_2_2 = (port_state_in_2_2_2 ^ port_key_2_2_2);
  assign port_state_out_2_2_3 = (port_state_in_2_2_3 ^ port_key_2_2_3);
  assign port_state_out_2_2_4 = (port_state_in_2_2_4 ^ port_key_2_2_4);
  assign port_state_out_2_2_5 = (port_state_in_2_2_5 ^ port_key_2_2_5);
  assign port_state_out_2_2_6 = (port_state_in_2_2_6 ^ port_key_2_2_6);
  assign port_state_out_2_2_7 = (port_state_in_2_2_7 ^ port_key_2_2_7);
  assign port_state_out_2_3_0 = (port_state_in_2_3_0 ^ port_key_2_3_0);
  assign port_state_out_2_3_1 = (port_state_in_2_3_1 ^ port_key_2_3_1);
  assign port_state_out_2_3_2 = (port_state_in_2_3_2 ^ port_key_2_3_2);
  assign port_state_out_2_3_3 = (port_state_in_2_3_3 ^ port_key_2_3_3);
  assign port_state_out_2_3_4 = (port_state_in_2_3_4 ^ port_key_2_3_4);
  assign port_state_out_2_3_5 = (port_state_in_2_3_5 ^ port_key_2_3_5);
  assign port_state_out_2_3_6 = (port_state_in_2_3_6 ^ port_key_2_3_6);
  assign port_state_out_2_3_7 = (port_state_in_2_3_7 ^ port_key_2_3_7);
  assign port_state_out_3_0_0 = (port_state_in_3_0_0 ^ port_key_3_0_0);
  assign port_state_out_3_0_1 = (port_state_in_3_0_1 ^ port_key_3_0_1);
  assign port_state_out_3_0_2 = (port_state_in_3_0_2 ^ port_key_3_0_2);
  assign port_state_out_3_0_3 = (port_state_in_3_0_3 ^ port_key_3_0_3);
  assign port_state_out_3_0_4 = (port_state_in_3_0_4 ^ port_key_3_0_4);
  assign port_state_out_3_0_5 = (port_state_in_3_0_5 ^ port_key_3_0_5);
  assign port_state_out_3_0_6 = (port_state_in_3_0_6 ^ port_key_3_0_6);
  assign port_state_out_3_0_7 = (port_state_in_3_0_7 ^ port_key_3_0_7);
  assign port_state_out_3_1_0 = (port_state_in_3_1_0 ^ port_key_3_1_0);
  assign port_state_out_3_1_1 = (port_state_in_3_1_1 ^ port_key_3_1_1);
  assign port_state_out_3_1_2 = (port_state_in_3_1_2 ^ port_key_3_1_2);
  assign port_state_out_3_1_3 = (port_state_in_3_1_3 ^ port_key_3_1_3);
  assign port_state_out_3_1_4 = (port_state_in_3_1_4 ^ port_key_3_1_4);
  assign port_state_out_3_1_5 = (port_state_in_3_1_5 ^ port_key_3_1_5);
  assign port_state_out_3_1_6 = (port_state_in_3_1_6 ^ port_key_3_1_6);
  assign port_state_out_3_1_7 = (port_state_in_3_1_7 ^ port_key_3_1_7);
  assign port_state_out_3_2_0 = (port_state_in_3_2_0 ^ port_key_3_2_0);
  assign port_state_out_3_2_1 = (port_state_in_3_2_1 ^ port_key_3_2_1);
  assign port_state_out_3_2_2 = (port_state_in_3_2_2 ^ port_key_3_2_2);
  assign port_state_out_3_2_3 = (port_state_in_3_2_3 ^ port_key_3_2_3);
  assign port_state_out_3_2_4 = (port_state_in_3_2_4 ^ port_key_3_2_4);
  assign port_state_out_3_2_5 = (port_state_in_3_2_5 ^ port_key_3_2_5);
  assign port_state_out_3_2_6 = (port_state_in_3_2_6 ^ port_key_3_2_6);
  assign port_state_out_3_2_7 = (port_state_in_3_2_7 ^ port_key_3_2_7);
  assign port_state_out_3_3_0 = (port_state_in_3_3_0 ^ port_key_3_3_0);
  assign port_state_out_3_3_1 = (port_state_in_3_3_1 ^ port_key_3_3_1);
  assign port_state_out_3_3_2 = (port_state_in_3_3_2 ^ port_key_3_3_2);
  assign port_state_out_3_3_3 = (port_state_in_3_3_3 ^ port_key_3_3_3);
  assign port_state_out_3_3_4 = (port_state_in_3_3_4 ^ port_key_3_3_4);
  assign port_state_out_3_3_5 = (port_state_in_3_3_5 ^ port_key_3_3_5);
  assign port_state_out_3_3_6 = (port_state_in_3_3_6 ^ port_key_3_3_6);
  assign port_state_out_3_3_7 = (port_state_in_3_3_7 ^ port_key_3_3_7);
  assign port_state_out_4_0_0 = (port_state_in_4_0_0 ^ port_key_4_0_0);
  assign port_state_out_4_0_1 = (port_state_in_4_0_1 ^ port_key_4_0_1);
  assign port_state_out_4_0_2 = (port_state_in_4_0_2 ^ port_key_4_0_2);
  assign port_state_out_4_0_3 = (port_state_in_4_0_3 ^ port_key_4_0_3);
  assign port_state_out_4_0_4 = (port_state_in_4_0_4 ^ port_key_4_0_4);
  assign port_state_out_4_0_5 = (port_state_in_4_0_5 ^ port_key_4_0_5);
  assign port_state_out_4_0_6 = (port_state_in_4_0_6 ^ port_key_4_0_6);
  assign port_state_out_4_0_7 = (port_state_in_4_0_7 ^ port_key_4_0_7);
  assign port_state_out_4_1_0 = (port_state_in_4_1_0 ^ port_key_4_1_0);
  assign port_state_out_4_1_1 = (port_state_in_4_1_1 ^ port_key_4_1_1);
  assign port_state_out_4_1_2 = (port_state_in_4_1_2 ^ port_key_4_1_2);
  assign port_state_out_4_1_3 = (port_state_in_4_1_3 ^ port_key_4_1_3);
  assign port_state_out_4_1_4 = (port_state_in_4_1_4 ^ port_key_4_1_4);
  assign port_state_out_4_1_5 = (port_state_in_4_1_5 ^ port_key_4_1_5);
  assign port_state_out_4_1_6 = (port_state_in_4_1_6 ^ port_key_4_1_6);
  assign port_state_out_4_1_7 = (port_state_in_4_1_7 ^ port_key_4_1_7);
  assign port_state_out_4_2_0 = (port_state_in_4_2_0 ^ port_key_4_2_0);
  assign port_state_out_4_2_1 = (port_state_in_4_2_1 ^ port_key_4_2_1);
  assign port_state_out_4_2_2 = (port_state_in_4_2_2 ^ port_key_4_2_2);
  assign port_state_out_4_2_3 = (port_state_in_4_2_3 ^ port_key_4_2_3);
  assign port_state_out_4_2_4 = (port_state_in_4_2_4 ^ port_key_4_2_4);
  assign port_state_out_4_2_5 = (port_state_in_4_2_5 ^ port_key_4_2_5);
  assign port_state_out_4_2_6 = (port_state_in_4_2_6 ^ port_key_4_2_6);
  assign port_state_out_4_2_7 = (port_state_in_4_2_7 ^ port_key_4_2_7);
  assign port_state_out_4_3_0 = (port_state_in_4_3_0 ^ port_key_4_3_0);
  assign port_state_out_4_3_1 = (port_state_in_4_3_1 ^ port_key_4_3_1);
  assign port_state_out_4_3_2 = (port_state_in_4_3_2 ^ port_key_4_3_2);
  assign port_state_out_4_3_3 = (port_state_in_4_3_3 ^ port_key_4_3_3);
  assign port_state_out_4_3_4 = (port_state_in_4_3_4 ^ port_key_4_3_4);
  assign port_state_out_4_3_5 = (port_state_in_4_3_5 ^ port_key_4_3_5);
  assign port_state_out_4_3_6 = (port_state_in_4_3_6 ^ port_key_4_3_6);
  assign port_state_out_4_3_7 = (port_state_in_4_3_7 ^ port_key_4_3_7);
  assign port_state_out_5_0_0 = (port_state_in_5_0_0 ^ port_key_5_0_0);
  assign port_state_out_5_0_1 = (port_state_in_5_0_1 ^ port_key_5_0_1);
  assign port_state_out_5_0_2 = (port_state_in_5_0_2 ^ port_key_5_0_2);
  assign port_state_out_5_0_3 = (port_state_in_5_0_3 ^ port_key_5_0_3);
  assign port_state_out_5_0_4 = (port_state_in_5_0_4 ^ port_key_5_0_4);
  assign port_state_out_5_0_5 = (port_state_in_5_0_5 ^ port_key_5_0_5);
  assign port_state_out_5_0_6 = (port_state_in_5_0_6 ^ port_key_5_0_6);
  assign port_state_out_5_0_7 = (port_state_in_5_0_7 ^ port_key_5_0_7);
  assign port_state_out_5_1_0 = (port_state_in_5_1_0 ^ port_key_5_1_0);
  assign port_state_out_5_1_1 = (port_state_in_5_1_1 ^ port_key_5_1_1);
  assign port_state_out_5_1_2 = (port_state_in_5_1_2 ^ port_key_5_1_2);
  assign port_state_out_5_1_3 = (port_state_in_5_1_3 ^ port_key_5_1_3);
  assign port_state_out_5_1_4 = (port_state_in_5_1_4 ^ port_key_5_1_4);
  assign port_state_out_5_1_5 = (port_state_in_5_1_5 ^ port_key_5_1_5);
  assign port_state_out_5_1_6 = (port_state_in_5_1_6 ^ port_key_5_1_6);
  assign port_state_out_5_1_7 = (port_state_in_5_1_7 ^ port_key_5_1_7);
  assign port_state_out_5_2_0 = (port_state_in_5_2_0 ^ port_key_5_2_0);
  assign port_state_out_5_2_1 = (port_state_in_5_2_1 ^ port_key_5_2_1);
  assign port_state_out_5_2_2 = (port_state_in_5_2_2 ^ port_key_5_2_2);
  assign port_state_out_5_2_3 = (port_state_in_5_2_3 ^ port_key_5_2_3);
  assign port_state_out_5_2_4 = (port_state_in_5_2_4 ^ port_key_5_2_4);
  assign port_state_out_5_2_5 = (port_state_in_5_2_5 ^ port_key_5_2_5);
  assign port_state_out_5_2_6 = (port_state_in_5_2_6 ^ port_key_5_2_6);
  assign port_state_out_5_2_7 = (port_state_in_5_2_7 ^ port_key_5_2_7);
  assign port_state_out_5_3_0 = (port_state_in_5_3_0 ^ port_key_5_3_0);
  assign port_state_out_5_3_1 = (port_state_in_5_3_1 ^ port_key_5_3_1);
  assign port_state_out_5_3_2 = (port_state_in_5_3_2 ^ port_key_5_3_2);
  assign port_state_out_5_3_3 = (port_state_in_5_3_3 ^ port_key_5_3_3);
  assign port_state_out_5_3_4 = (port_state_in_5_3_4 ^ port_key_5_3_4);
  assign port_state_out_5_3_5 = (port_state_in_5_3_5 ^ port_key_5_3_5);
  assign port_state_out_5_3_6 = (port_state_in_5_3_6 ^ port_key_5_3_6);
  assign port_state_out_5_3_7 = (port_state_in_5_3_7 ^ port_key_5_3_7);
  assign port_state_out_6_0_0 = (port_state_in_6_0_0 ^ port_key_6_0_0);
  assign port_state_out_6_0_1 = (port_state_in_6_0_1 ^ port_key_6_0_1);
  assign port_state_out_6_0_2 = (port_state_in_6_0_2 ^ port_key_6_0_2);
  assign port_state_out_6_0_3 = (port_state_in_6_0_3 ^ port_key_6_0_3);
  assign port_state_out_6_0_4 = (port_state_in_6_0_4 ^ port_key_6_0_4);
  assign port_state_out_6_0_5 = (port_state_in_6_0_5 ^ port_key_6_0_5);
  assign port_state_out_6_0_6 = (port_state_in_6_0_6 ^ port_key_6_0_6);
  assign port_state_out_6_0_7 = (port_state_in_6_0_7 ^ port_key_6_0_7);
  assign port_state_out_6_1_0 = (port_state_in_6_1_0 ^ port_key_6_1_0);
  assign port_state_out_6_1_1 = (port_state_in_6_1_1 ^ port_key_6_1_1);
  assign port_state_out_6_1_2 = (port_state_in_6_1_2 ^ port_key_6_1_2);
  assign port_state_out_6_1_3 = (port_state_in_6_1_3 ^ port_key_6_1_3);
  assign port_state_out_6_1_4 = (port_state_in_6_1_4 ^ port_key_6_1_4);
  assign port_state_out_6_1_5 = (port_state_in_6_1_5 ^ port_key_6_1_5);
  assign port_state_out_6_1_6 = (port_state_in_6_1_6 ^ port_key_6_1_6);
  assign port_state_out_6_1_7 = (port_state_in_6_1_7 ^ port_key_6_1_7);
  assign port_state_out_6_2_0 = (port_state_in_6_2_0 ^ port_key_6_2_0);
  assign port_state_out_6_2_1 = (port_state_in_6_2_1 ^ port_key_6_2_1);
  assign port_state_out_6_2_2 = (port_state_in_6_2_2 ^ port_key_6_2_2);
  assign port_state_out_6_2_3 = (port_state_in_6_2_3 ^ port_key_6_2_3);
  assign port_state_out_6_2_4 = (port_state_in_6_2_4 ^ port_key_6_2_4);
  assign port_state_out_6_2_5 = (port_state_in_6_2_5 ^ port_key_6_2_5);
  assign port_state_out_6_2_6 = (port_state_in_6_2_6 ^ port_key_6_2_6);
  assign port_state_out_6_2_7 = (port_state_in_6_2_7 ^ port_key_6_2_7);
  assign port_state_out_6_3_0 = (port_state_in_6_3_0 ^ port_key_6_3_0);
  assign port_state_out_6_3_1 = (port_state_in_6_3_1 ^ port_key_6_3_1);
  assign port_state_out_6_3_2 = (port_state_in_6_3_2 ^ port_key_6_3_2);
  assign port_state_out_6_3_3 = (port_state_in_6_3_3 ^ port_key_6_3_3);
  assign port_state_out_6_3_4 = (port_state_in_6_3_4 ^ port_key_6_3_4);
  assign port_state_out_6_3_5 = (port_state_in_6_3_5 ^ port_key_6_3_5);
  assign port_state_out_6_3_6 = (port_state_in_6_3_6 ^ port_key_6_3_6);
  assign port_state_out_6_3_7 = (port_state_in_6_3_7 ^ port_key_6_3_7);
  assign port_state_out_7_0_0 = (port_state_in_7_0_0 ^ port_key_7_0_0);
  assign port_state_out_7_0_1 = (port_state_in_7_0_1 ^ port_key_7_0_1);
  assign port_state_out_7_0_2 = (port_state_in_7_0_2 ^ port_key_7_0_2);
  assign port_state_out_7_0_3 = (port_state_in_7_0_3 ^ port_key_7_0_3);
  assign port_state_out_7_0_4 = (port_state_in_7_0_4 ^ port_key_7_0_4);
  assign port_state_out_7_0_5 = (port_state_in_7_0_5 ^ port_key_7_0_5);
  assign port_state_out_7_0_6 = (port_state_in_7_0_6 ^ port_key_7_0_6);
  assign port_state_out_7_0_7 = (port_state_in_7_0_7 ^ port_key_7_0_7);
  assign port_state_out_7_1_0 = (port_state_in_7_1_0 ^ port_key_7_1_0);
  assign port_state_out_7_1_1 = (port_state_in_7_1_1 ^ port_key_7_1_1);
  assign port_state_out_7_1_2 = (port_state_in_7_1_2 ^ port_key_7_1_2);
  assign port_state_out_7_1_3 = (port_state_in_7_1_3 ^ port_key_7_1_3);
  assign port_state_out_7_1_4 = (port_state_in_7_1_4 ^ port_key_7_1_4);
  assign port_state_out_7_1_5 = (port_state_in_7_1_5 ^ port_key_7_1_5);
  assign port_state_out_7_1_6 = (port_state_in_7_1_6 ^ port_key_7_1_6);
  assign port_state_out_7_1_7 = (port_state_in_7_1_7 ^ port_key_7_1_7);
  assign port_state_out_7_2_0 = (port_state_in_7_2_0 ^ port_key_7_2_0);
  assign port_state_out_7_2_1 = (port_state_in_7_2_1 ^ port_key_7_2_1);
  assign port_state_out_7_2_2 = (port_state_in_7_2_2 ^ port_key_7_2_2);
  assign port_state_out_7_2_3 = (port_state_in_7_2_3 ^ port_key_7_2_3);
  assign port_state_out_7_2_4 = (port_state_in_7_2_4 ^ port_key_7_2_4);
  assign port_state_out_7_2_5 = (port_state_in_7_2_5 ^ port_key_7_2_5);
  assign port_state_out_7_2_6 = (port_state_in_7_2_6 ^ port_key_7_2_6);
  assign port_state_out_7_2_7 = (port_state_in_7_2_7 ^ port_key_7_2_7);
  assign port_state_out_7_3_0 = (port_state_in_7_3_0 ^ port_key_7_3_0);
  assign port_state_out_7_3_1 = (port_state_in_7_3_1 ^ port_key_7_3_1);
  assign port_state_out_7_3_2 = (port_state_in_7_3_2 ^ port_key_7_3_2);
  assign port_state_out_7_3_3 = (port_state_in_7_3_3 ^ port_key_7_3_3);
  assign port_state_out_7_3_4 = (port_state_in_7_3_4 ^ port_key_7_3_4);
  assign port_state_out_7_3_5 = (port_state_in_7_3_5 ^ port_key_7_3_5);
  assign port_state_out_7_3_6 = (port_state_in_7_3_6 ^ port_key_7_3_6);
  assign port_state_out_7_3_7 = (port_state_in_7_3_7 ^ port_key_7_3_7);
  assign port_state_out_8_0_0 = (port_state_in_8_0_0 ^ port_key_8_0_0);
  assign port_state_out_8_0_1 = (port_state_in_8_0_1 ^ port_key_8_0_1);
  assign port_state_out_8_0_2 = (port_state_in_8_0_2 ^ port_key_8_0_2);
  assign port_state_out_8_0_3 = (port_state_in_8_0_3 ^ port_key_8_0_3);
  assign port_state_out_8_0_4 = (port_state_in_8_0_4 ^ port_key_8_0_4);
  assign port_state_out_8_0_5 = (port_state_in_8_0_5 ^ port_key_8_0_5);
  assign port_state_out_8_0_6 = (port_state_in_8_0_6 ^ port_key_8_0_6);
  assign port_state_out_8_0_7 = (port_state_in_8_0_7 ^ port_key_8_0_7);
  assign port_state_out_8_1_0 = (port_state_in_8_1_0 ^ port_key_8_1_0);
  assign port_state_out_8_1_1 = (port_state_in_8_1_1 ^ port_key_8_1_1);
  assign port_state_out_8_1_2 = (port_state_in_8_1_2 ^ port_key_8_1_2);
  assign port_state_out_8_1_3 = (port_state_in_8_1_3 ^ port_key_8_1_3);
  assign port_state_out_8_1_4 = (port_state_in_8_1_4 ^ port_key_8_1_4);
  assign port_state_out_8_1_5 = (port_state_in_8_1_5 ^ port_key_8_1_5);
  assign port_state_out_8_1_6 = (port_state_in_8_1_6 ^ port_key_8_1_6);
  assign port_state_out_8_1_7 = (port_state_in_8_1_7 ^ port_key_8_1_7);
  assign port_state_out_8_2_0 = (port_state_in_8_2_0 ^ port_key_8_2_0);
  assign port_state_out_8_2_1 = (port_state_in_8_2_1 ^ port_key_8_2_1);
  assign port_state_out_8_2_2 = (port_state_in_8_2_2 ^ port_key_8_2_2);
  assign port_state_out_8_2_3 = (port_state_in_8_2_3 ^ port_key_8_2_3);
  assign port_state_out_8_2_4 = (port_state_in_8_2_4 ^ port_key_8_2_4);
  assign port_state_out_8_2_5 = (port_state_in_8_2_5 ^ port_key_8_2_5);
  assign port_state_out_8_2_6 = (port_state_in_8_2_6 ^ port_key_8_2_6);
  assign port_state_out_8_2_7 = (port_state_in_8_2_7 ^ port_key_8_2_7);
  assign port_state_out_8_3_0 = (port_state_in_8_3_0 ^ port_key_8_3_0);
  assign port_state_out_8_3_1 = (port_state_in_8_3_1 ^ port_key_8_3_1);
  assign port_state_out_8_3_2 = (port_state_in_8_3_2 ^ port_key_8_3_2);
  assign port_state_out_8_3_3 = (port_state_in_8_3_3 ^ port_key_8_3_3);
  assign port_state_out_8_3_4 = (port_state_in_8_3_4 ^ port_key_8_3_4);
  assign port_state_out_8_3_5 = (port_state_in_8_3_5 ^ port_key_8_3_5);
  assign port_state_out_8_3_6 = (port_state_in_8_3_6 ^ port_key_8_3_6);
  assign port_state_out_8_3_7 = (port_state_in_8_3_7 ^ port_key_8_3_7);
  assign port_state_out_9_0_0 = (port_state_in_9_0_0 ^ port_key_9_0_0);
  assign port_state_out_9_0_1 = (port_state_in_9_0_1 ^ port_key_9_0_1);
  assign port_state_out_9_0_2 = (port_state_in_9_0_2 ^ port_key_9_0_2);
  assign port_state_out_9_0_3 = (port_state_in_9_0_3 ^ port_key_9_0_3);
  assign port_state_out_9_0_4 = (port_state_in_9_0_4 ^ port_key_9_0_4);
  assign port_state_out_9_0_5 = (port_state_in_9_0_5 ^ port_key_9_0_5);
  assign port_state_out_9_0_6 = (port_state_in_9_0_6 ^ port_key_9_0_6);
  assign port_state_out_9_0_7 = (port_state_in_9_0_7 ^ port_key_9_0_7);
  assign port_state_out_9_1_0 = (port_state_in_9_1_0 ^ port_key_9_1_0);
  assign port_state_out_9_1_1 = (port_state_in_9_1_1 ^ port_key_9_1_1);
  assign port_state_out_9_1_2 = (port_state_in_9_1_2 ^ port_key_9_1_2);
  assign port_state_out_9_1_3 = (port_state_in_9_1_3 ^ port_key_9_1_3);
  assign port_state_out_9_1_4 = (port_state_in_9_1_4 ^ port_key_9_1_4);
  assign port_state_out_9_1_5 = (port_state_in_9_1_5 ^ port_key_9_1_5);
  assign port_state_out_9_1_6 = (port_state_in_9_1_6 ^ port_key_9_1_6);
  assign port_state_out_9_1_7 = (port_state_in_9_1_7 ^ port_key_9_1_7);
  assign port_state_out_9_2_0 = (port_state_in_9_2_0 ^ port_key_9_2_0);
  assign port_state_out_9_2_1 = (port_state_in_9_2_1 ^ port_key_9_2_1);
  assign port_state_out_9_2_2 = (port_state_in_9_2_2 ^ port_key_9_2_2);
  assign port_state_out_9_2_3 = (port_state_in_9_2_3 ^ port_key_9_2_3);
  assign port_state_out_9_2_4 = (port_state_in_9_2_4 ^ port_key_9_2_4);
  assign port_state_out_9_2_5 = (port_state_in_9_2_5 ^ port_key_9_2_5);
  assign port_state_out_9_2_6 = (port_state_in_9_2_6 ^ port_key_9_2_6);
  assign port_state_out_9_2_7 = (port_state_in_9_2_7 ^ port_key_9_2_7);
  assign port_state_out_9_3_0 = (port_state_in_9_3_0 ^ port_key_9_3_0);
  assign port_state_out_9_3_1 = (port_state_in_9_3_1 ^ port_key_9_3_1);
  assign port_state_out_9_3_2 = (port_state_in_9_3_2 ^ port_key_9_3_2);
  assign port_state_out_9_3_3 = (port_state_in_9_3_3 ^ port_key_9_3_3);
  assign port_state_out_9_3_4 = (port_state_in_9_3_4 ^ port_key_9_3_4);
  assign port_state_out_9_3_5 = (port_state_in_9_3_5 ^ port_key_9_3_5);
  assign port_state_out_9_3_6 = (port_state_in_9_3_6 ^ port_key_9_3_6);
  assign port_state_out_9_3_7 = (port_state_in_9_3_7 ^ port_key_9_3_7);
  assign port_state_out_10_0_0 = (port_state_in_10_0_0 ^ port_key_10_0_0);
  assign port_state_out_10_0_1 = (port_state_in_10_0_1 ^ port_key_10_0_1);
  assign port_state_out_10_0_2 = (port_state_in_10_0_2 ^ port_key_10_0_2);
  assign port_state_out_10_0_3 = (port_state_in_10_0_3 ^ port_key_10_0_3);
  assign port_state_out_10_0_4 = (port_state_in_10_0_4 ^ port_key_10_0_4);
  assign port_state_out_10_0_5 = (port_state_in_10_0_5 ^ port_key_10_0_5);
  assign port_state_out_10_0_6 = (port_state_in_10_0_6 ^ port_key_10_0_6);
  assign port_state_out_10_0_7 = (port_state_in_10_0_7 ^ port_key_10_0_7);
  assign port_state_out_10_1_0 = (port_state_in_10_1_0 ^ port_key_10_1_0);
  assign port_state_out_10_1_1 = (port_state_in_10_1_1 ^ port_key_10_1_1);
  assign port_state_out_10_1_2 = (port_state_in_10_1_2 ^ port_key_10_1_2);
  assign port_state_out_10_1_3 = (port_state_in_10_1_3 ^ port_key_10_1_3);
  assign port_state_out_10_1_4 = (port_state_in_10_1_4 ^ port_key_10_1_4);
  assign port_state_out_10_1_5 = (port_state_in_10_1_5 ^ port_key_10_1_5);
  assign port_state_out_10_1_6 = (port_state_in_10_1_6 ^ port_key_10_1_6);
  assign port_state_out_10_1_7 = (port_state_in_10_1_7 ^ port_key_10_1_7);
  assign port_state_out_10_2_0 = (port_state_in_10_2_0 ^ port_key_10_2_0);
  assign port_state_out_10_2_1 = (port_state_in_10_2_1 ^ port_key_10_2_1);
  assign port_state_out_10_2_2 = (port_state_in_10_2_2 ^ port_key_10_2_2);
  assign port_state_out_10_2_3 = (port_state_in_10_2_3 ^ port_key_10_2_3);
  assign port_state_out_10_2_4 = (port_state_in_10_2_4 ^ port_key_10_2_4);
  assign port_state_out_10_2_5 = (port_state_in_10_2_5 ^ port_key_10_2_5);
  assign port_state_out_10_2_6 = (port_state_in_10_2_6 ^ port_key_10_2_6);
  assign port_state_out_10_2_7 = (port_state_in_10_2_7 ^ port_key_10_2_7);
  assign port_state_out_10_3_0 = (port_state_in_10_3_0 ^ port_key_10_3_0);
  assign port_state_out_10_3_1 = (port_state_in_10_3_1 ^ port_key_10_3_1);
  assign port_state_out_10_3_2 = (port_state_in_10_3_2 ^ port_key_10_3_2);
  assign port_state_out_10_3_3 = (port_state_in_10_3_3 ^ port_key_10_3_3);
  assign port_state_out_10_3_4 = (port_state_in_10_3_4 ^ port_key_10_3_4);
  assign port_state_out_10_3_5 = (port_state_in_10_3_5 ^ port_key_10_3_5);
  assign port_state_out_10_3_6 = (port_state_in_10_3_6 ^ port_key_10_3_6);
  assign port_state_out_10_3_7 = (port_state_in_10_3_7 ^ port_key_10_3_7);
  assign port_state_out_11_0_0 = (port_state_in_11_0_0 ^ port_key_11_0_0);
  assign port_state_out_11_0_1 = (port_state_in_11_0_1 ^ port_key_11_0_1);
  assign port_state_out_11_0_2 = (port_state_in_11_0_2 ^ port_key_11_0_2);
  assign port_state_out_11_0_3 = (port_state_in_11_0_3 ^ port_key_11_0_3);
  assign port_state_out_11_0_4 = (port_state_in_11_0_4 ^ port_key_11_0_4);
  assign port_state_out_11_0_5 = (port_state_in_11_0_5 ^ port_key_11_0_5);
  assign port_state_out_11_0_6 = (port_state_in_11_0_6 ^ port_key_11_0_6);
  assign port_state_out_11_0_7 = (port_state_in_11_0_7 ^ port_key_11_0_7);
  assign port_state_out_11_1_0 = (port_state_in_11_1_0 ^ port_key_11_1_0);
  assign port_state_out_11_1_1 = (port_state_in_11_1_1 ^ port_key_11_1_1);
  assign port_state_out_11_1_2 = (port_state_in_11_1_2 ^ port_key_11_1_2);
  assign port_state_out_11_1_3 = (port_state_in_11_1_3 ^ port_key_11_1_3);
  assign port_state_out_11_1_4 = (port_state_in_11_1_4 ^ port_key_11_1_4);
  assign port_state_out_11_1_5 = (port_state_in_11_1_5 ^ port_key_11_1_5);
  assign port_state_out_11_1_6 = (port_state_in_11_1_6 ^ port_key_11_1_6);
  assign port_state_out_11_1_7 = (port_state_in_11_1_7 ^ port_key_11_1_7);
  assign port_state_out_11_2_0 = (port_state_in_11_2_0 ^ port_key_11_2_0);
  assign port_state_out_11_2_1 = (port_state_in_11_2_1 ^ port_key_11_2_1);
  assign port_state_out_11_2_2 = (port_state_in_11_2_2 ^ port_key_11_2_2);
  assign port_state_out_11_2_3 = (port_state_in_11_2_3 ^ port_key_11_2_3);
  assign port_state_out_11_2_4 = (port_state_in_11_2_4 ^ port_key_11_2_4);
  assign port_state_out_11_2_5 = (port_state_in_11_2_5 ^ port_key_11_2_5);
  assign port_state_out_11_2_6 = (port_state_in_11_2_6 ^ port_key_11_2_6);
  assign port_state_out_11_2_7 = (port_state_in_11_2_7 ^ port_key_11_2_7);
  assign port_state_out_11_3_0 = (port_state_in_11_3_0 ^ port_key_11_3_0);
  assign port_state_out_11_3_1 = (port_state_in_11_3_1 ^ port_key_11_3_1);
  assign port_state_out_11_3_2 = (port_state_in_11_3_2 ^ port_key_11_3_2);
  assign port_state_out_11_3_3 = (port_state_in_11_3_3 ^ port_key_11_3_3);
  assign port_state_out_11_3_4 = (port_state_in_11_3_4 ^ port_key_11_3_4);
  assign port_state_out_11_3_5 = (port_state_in_11_3_5 ^ port_key_11_3_5);
  assign port_state_out_11_3_6 = (port_state_in_11_3_6 ^ port_key_11_3_6);
  assign port_state_out_11_3_7 = (port_state_in_11_3_7 ^ port_key_11_3_7);
  assign port_state_out_12_0_0 = (port_state_in_12_0_0 ^ port_key_12_0_0);
  assign port_state_out_12_0_1 = (port_state_in_12_0_1 ^ port_key_12_0_1);
  assign port_state_out_12_0_2 = (port_state_in_12_0_2 ^ port_key_12_0_2);
  assign port_state_out_12_0_3 = (port_state_in_12_0_3 ^ port_key_12_0_3);
  assign port_state_out_12_0_4 = (port_state_in_12_0_4 ^ port_key_12_0_4);
  assign port_state_out_12_0_5 = (port_state_in_12_0_5 ^ port_key_12_0_5);
  assign port_state_out_12_0_6 = (port_state_in_12_0_6 ^ port_key_12_0_6);
  assign port_state_out_12_0_7 = (port_state_in_12_0_7 ^ port_key_12_0_7);
  assign port_state_out_12_1_0 = (port_state_in_12_1_0 ^ port_key_12_1_0);
  assign port_state_out_12_1_1 = (port_state_in_12_1_1 ^ port_key_12_1_1);
  assign port_state_out_12_1_2 = (port_state_in_12_1_2 ^ port_key_12_1_2);
  assign port_state_out_12_1_3 = (port_state_in_12_1_3 ^ port_key_12_1_3);
  assign port_state_out_12_1_4 = (port_state_in_12_1_4 ^ port_key_12_1_4);
  assign port_state_out_12_1_5 = (port_state_in_12_1_5 ^ port_key_12_1_5);
  assign port_state_out_12_1_6 = (port_state_in_12_1_6 ^ port_key_12_1_6);
  assign port_state_out_12_1_7 = (port_state_in_12_1_7 ^ port_key_12_1_7);
  assign port_state_out_12_2_0 = (port_state_in_12_2_0 ^ port_key_12_2_0);
  assign port_state_out_12_2_1 = (port_state_in_12_2_1 ^ port_key_12_2_1);
  assign port_state_out_12_2_2 = (port_state_in_12_2_2 ^ port_key_12_2_2);
  assign port_state_out_12_2_3 = (port_state_in_12_2_3 ^ port_key_12_2_3);
  assign port_state_out_12_2_4 = (port_state_in_12_2_4 ^ port_key_12_2_4);
  assign port_state_out_12_2_5 = (port_state_in_12_2_5 ^ port_key_12_2_5);
  assign port_state_out_12_2_6 = (port_state_in_12_2_6 ^ port_key_12_2_6);
  assign port_state_out_12_2_7 = (port_state_in_12_2_7 ^ port_key_12_2_7);
  assign port_state_out_12_3_0 = (port_state_in_12_3_0 ^ port_key_12_3_0);
  assign port_state_out_12_3_1 = (port_state_in_12_3_1 ^ port_key_12_3_1);
  assign port_state_out_12_3_2 = (port_state_in_12_3_2 ^ port_key_12_3_2);
  assign port_state_out_12_3_3 = (port_state_in_12_3_3 ^ port_key_12_3_3);
  assign port_state_out_12_3_4 = (port_state_in_12_3_4 ^ port_key_12_3_4);
  assign port_state_out_12_3_5 = (port_state_in_12_3_5 ^ port_key_12_3_5);
  assign port_state_out_12_3_6 = (port_state_in_12_3_6 ^ port_key_12_3_6);
  assign port_state_out_12_3_7 = (port_state_in_12_3_7 ^ port_key_12_3_7);
  assign port_state_out_13_0_0 = (port_state_in_13_0_0 ^ port_key_13_0_0);
  assign port_state_out_13_0_1 = (port_state_in_13_0_1 ^ port_key_13_0_1);
  assign port_state_out_13_0_2 = (port_state_in_13_0_2 ^ port_key_13_0_2);
  assign port_state_out_13_0_3 = (port_state_in_13_0_3 ^ port_key_13_0_3);
  assign port_state_out_13_0_4 = (port_state_in_13_0_4 ^ port_key_13_0_4);
  assign port_state_out_13_0_5 = (port_state_in_13_0_5 ^ port_key_13_0_5);
  assign port_state_out_13_0_6 = (port_state_in_13_0_6 ^ port_key_13_0_6);
  assign port_state_out_13_0_7 = (port_state_in_13_0_7 ^ port_key_13_0_7);
  assign port_state_out_13_1_0 = (port_state_in_13_1_0 ^ port_key_13_1_0);
  assign port_state_out_13_1_1 = (port_state_in_13_1_1 ^ port_key_13_1_1);
  assign port_state_out_13_1_2 = (port_state_in_13_1_2 ^ port_key_13_1_2);
  assign port_state_out_13_1_3 = (port_state_in_13_1_3 ^ port_key_13_1_3);
  assign port_state_out_13_1_4 = (port_state_in_13_1_4 ^ port_key_13_1_4);
  assign port_state_out_13_1_5 = (port_state_in_13_1_5 ^ port_key_13_1_5);
  assign port_state_out_13_1_6 = (port_state_in_13_1_6 ^ port_key_13_1_6);
  assign port_state_out_13_1_7 = (port_state_in_13_1_7 ^ port_key_13_1_7);
  assign port_state_out_13_2_0 = (port_state_in_13_2_0 ^ port_key_13_2_0);
  assign port_state_out_13_2_1 = (port_state_in_13_2_1 ^ port_key_13_2_1);
  assign port_state_out_13_2_2 = (port_state_in_13_2_2 ^ port_key_13_2_2);
  assign port_state_out_13_2_3 = (port_state_in_13_2_3 ^ port_key_13_2_3);
  assign port_state_out_13_2_4 = (port_state_in_13_2_4 ^ port_key_13_2_4);
  assign port_state_out_13_2_5 = (port_state_in_13_2_5 ^ port_key_13_2_5);
  assign port_state_out_13_2_6 = (port_state_in_13_2_6 ^ port_key_13_2_6);
  assign port_state_out_13_2_7 = (port_state_in_13_2_7 ^ port_key_13_2_7);
  assign port_state_out_13_3_0 = (port_state_in_13_3_0 ^ port_key_13_3_0);
  assign port_state_out_13_3_1 = (port_state_in_13_3_1 ^ port_key_13_3_1);
  assign port_state_out_13_3_2 = (port_state_in_13_3_2 ^ port_key_13_3_2);
  assign port_state_out_13_3_3 = (port_state_in_13_3_3 ^ port_key_13_3_3);
  assign port_state_out_13_3_4 = (port_state_in_13_3_4 ^ port_key_13_3_4);
  assign port_state_out_13_3_5 = (port_state_in_13_3_5 ^ port_key_13_3_5);
  assign port_state_out_13_3_6 = (port_state_in_13_3_6 ^ port_key_13_3_6);
  assign port_state_out_13_3_7 = (port_state_in_13_3_7 ^ port_key_13_3_7);
  assign port_state_out_14_0_0 = (port_state_in_14_0_0 ^ port_key_14_0_0);
  assign port_state_out_14_0_1 = (port_state_in_14_0_1 ^ port_key_14_0_1);
  assign port_state_out_14_0_2 = (port_state_in_14_0_2 ^ port_key_14_0_2);
  assign port_state_out_14_0_3 = (port_state_in_14_0_3 ^ port_key_14_0_3);
  assign port_state_out_14_0_4 = (port_state_in_14_0_4 ^ port_key_14_0_4);
  assign port_state_out_14_0_5 = (port_state_in_14_0_5 ^ port_key_14_0_5);
  assign port_state_out_14_0_6 = (port_state_in_14_0_6 ^ port_key_14_0_6);
  assign port_state_out_14_0_7 = (port_state_in_14_0_7 ^ port_key_14_0_7);
  assign port_state_out_14_1_0 = (port_state_in_14_1_0 ^ port_key_14_1_0);
  assign port_state_out_14_1_1 = (port_state_in_14_1_1 ^ port_key_14_1_1);
  assign port_state_out_14_1_2 = (port_state_in_14_1_2 ^ port_key_14_1_2);
  assign port_state_out_14_1_3 = (port_state_in_14_1_3 ^ port_key_14_1_3);
  assign port_state_out_14_1_4 = (port_state_in_14_1_4 ^ port_key_14_1_4);
  assign port_state_out_14_1_5 = (port_state_in_14_1_5 ^ port_key_14_1_5);
  assign port_state_out_14_1_6 = (port_state_in_14_1_6 ^ port_key_14_1_6);
  assign port_state_out_14_1_7 = (port_state_in_14_1_7 ^ port_key_14_1_7);
  assign port_state_out_14_2_0 = (port_state_in_14_2_0 ^ port_key_14_2_0);
  assign port_state_out_14_2_1 = (port_state_in_14_2_1 ^ port_key_14_2_1);
  assign port_state_out_14_2_2 = (port_state_in_14_2_2 ^ port_key_14_2_2);
  assign port_state_out_14_2_3 = (port_state_in_14_2_3 ^ port_key_14_2_3);
  assign port_state_out_14_2_4 = (port_state_in_14_2_4 ^ port_key_14_2_4);
  assign port_state_out_14_2_5 = (port_state_in_14_2_5 ^ port_key_14_2_5);
  assign port_state_out_14_2_6 = (port_state_in_14_2_6 ^ port_key_14_2_6);
  assign port_state_out_14_2_7 = (port_state_in_14_2_7 ^ port_key_14_2_7);
  assign port_state_out_14_3_0 = (port_state_in_14_3_0 ^ port_key_14_3_0);
  assign port_state_out_14_3_1 = (port_state_in_14_3_1 ^ port_key_14_3_1);
  assign port_state_out_14_3_2 = (port_state_in_14_3_2 ^ port_key_14_3_2);
  assign port_state_out_14_3_3 = (port_state_in_14_3_3 ^ port_key_14_3_3);
  assign port_state_out_14_3_4 = (port_state_in_14_3_4 ^ port_key_14_3_4);
  assign port_state_out_14_3_5 = (port_state_in_14_3_5 ^ port_key_14_3_5);
  assign port_state_out_14_3_6 = (port_state_in_14_3_6 ^ port_key_14_3_6);
  assign port_state_out_14_3_7 = (port_state_in_14_3_7 ^ port_key_14_3_7);
  assign port_state_out_15_0_0 = (port_state_in_15_0_0 ^ port_key_15_0_0);
  assign port_state_out_15_0_1 = (port_state_in_15_0_1 ^ port_key_15_0_1);
  assign port_state_out_15_0_2 = (port_state_in_15_0_2 ^ port_key_15_0_2);
  assign port_state_out_15_0_3 = (port_state_in_15_0_3 ^ port_key_15_0_3);
  assign port_state_out_15_0_4 = (port_state_in_15_0_4 ^ port_key_15_0_4);
  assign port_state_out_15_0_5 = (port_state_in_15_0_5 ^ port_key_15_0_5);
  assign port_state_out_15_0_6 = (port_state_in_15_0_6 ^ port_key_15_0_6);
  assign port_state_out_15_0_7 = (port_state_in_15_0_7 ^ port_key_15_0_7);
  assign port_state_out_15_1_0 = (port_state_in_15_1_0 ^ port_key_15_1_0);
  assign port_state_out_15_1_1 = (port_state_in_15_1_1 ^ port_key_15_1_1);
  assign port_state_out_15_1_2 = (port_state_in_15_1_2 ^ port_key_15_1_2);
  assign port_state_out_15_1_3 = (port_state_in_15_1_3 ^ port_key_15_1_3);
  assign port_state_out_15_1_4 = (port_state_in_15_1_4 ^ port_key_15_1_4);
  assign port_state_out_15_1_5 = (port_state_in_15_1_5 ^ port_key_15_1_5);
  assign port_state_out_15_1_6 = (port_state_in_15_1_6 ^ port_key_15_1_6);
  assign port_state_out_15_1_7 = (port_state_in_15_1_7 ^ port_key_15_1_7);
  assign port_state_out_15_2_0 = (port_state_in_15_2_0 ^ port_key_15_2_0);
  assign port_state_out_15_2_1 = (port_state_in_15_2_1 ^ port_key_15_2_1);
  assign port_state_out_15_2_2 = (port_state_in_15_2_2 ^ port_key_15_2_2);
  assign port_state_out_15_2_3 = (port_state_in_15_2_3 ^ port_key_15_2_3);
  assign port_state_out_15_2_4 = (port_state_in_15_2_4 ^ port_key_15_2_4);
  assign port_state_out_15_2_5 = (port_state_in_15_2_5 ^ port_key_15_2_5);
  assign port_state_out_15_2_6 = (port_state_in_15_2_6 ^ port_key_15_2_6);
  assign port_state_out_15_2_7 = (port_state_in_15_2_7 ^ port_key_15_2_7);
  assign port_state_out_15_3_0 = (port_state_in_15_3_0 ^ port_key_15_3_0);
  assign port_state_out_15_3_1 = (port_state_in_15_3_1 ^ port_key_15_3_1);
  assign port_state_out_15_3_2 = (port_state_in_15_3_2 ^ port_key_15_3_2);
  assign port_state_out_15_3_3 = (port_state_in_15_3_3 ^ port_key_15_3_3);
  assign port_state_out_15_3_4 = (port_state_in_15_3_4 ^ port_key_15_3_4);
  assign port_state_out_15_3_5 = (port_state_in_15_3_5 ^ port_key_15_3_5);
  assign port_state_out_15_3_6 = (port_state_in_15_3_6 ^ port_key_15_3_6);
  assign port_state_out_15_3_7 = (port_state_in_15_3_7 ^ port_key_15_3_7);

endmodule

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

module Mul3 (
  input      [0:0]    port_byte_in_0,
  input      [0:0]    port_byte_in_1,
  input      [0:0]    port_byte_in_2,
  input      [0:0]    port_byte_in_3,
  input      [0:0]    port_byte_in_4,
  input      [0:0]    port_byte_in_5,
  input      [0:0]    port_byte_in_6,
  input      [0:0]    port_byte_in_7,
  output     [0:0]    port_byte_out_0,
  output     [0:0]    port_byte_out_1,
  output     [0:0]    port_byte_out_2,
  output     [0:0]    port_byte_out_3,
  output     [0:0]    port_byte_out_4,
  output     [0:0]    port_byte_out_5,
  output     [0:0]    port_byte_out_6,
  output     [0:0]    port_byte_out_7
);


  assign port_byte_out_7 = (port_byte_in_7 ^ port_byte_in_6);
  assign port_byte_out_6 = (port_byte_in_6 ^ port_byte_in_5);
  assign port_byte_out_5 = (port_byte_in_5 ^ port_byte_in_4);
  assign port_byte_out_4 = ((port_byte_in_7 ^ port_byte_in_4) ^ port_byte_in_3);
  assign port_byte_out_3 = ((port_byte_in_7 ^ port_byte_in_3) ^ port_byte_in_2);
  assign port_byte_out_2 = (port_byte_in_2 ^ port_byte_in_1);
  assign port_byte_out_1 = ((port_byte_in_7 ^ port_byte_in_1) ^ port_byte_in_0);
  assign port_byte_out_0 = (port_byte_in_7 ^ port_byte_in_0);

endmodule

module Mul2 (
  input      [0:0]    port_byte_in_0,
  input      [0:0]    port_byte_in_1,
  input      [0:0]    port_byte_in_2,
  input      [0:0]    port_byte_in_3,
  input      [0:0]    port_byte_in_4,
  input      [0:0]    port_byte_in_5,
  input      [0:0]    port_byte_in_6,
  input      [0:0]    port_byte_in_7,
  output     [0:0]    port_byte_out_0,
  output     [0:0]    port_byte_out_1,
  output     [0:0]    port_byte_out_2,
  output     [0:0]    port_byte_out_3,
  output     [0:0]    port_byte_out_4,
  output     [0:0]    port_byte_out_5,
  output     [0:0]    port_byte_out_6,
  output     [0:0]    port_byte_out_7
);


  assign port_byte_out_7 = port_byte_in_6;
  assign port_byte_out_6 = port_byte_in_5;
  assign port_byte_out_5 = port_byte_in_4;
  assign port_byte_out_4 = (port_byte_in_7 ^ port_byte_in_3);
  assign port_byte_out_3 = (port_byte_in_7 ^ port_byte_in_2);
  assign port_byte_out_2 = port_byte_in_1;
  assign port_byte_out_1 = (port_byte_in_7 ^ port_byte_in_0);
  assign port_byte_out_0 = port_byte_in_7;

endmodule

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

module Addition_Inv_TI (
  input      [0:0]    port_x0_0,
  input      [0:0]    port_x0_1,
  input      [0:0]    port_x0_2,
  input      [0:0]    port_x0_3,
  input      [0:0]    port_x1_0,
  input      [0:0]    port_x1_1,
  input      [0:0]    port_x1_2,
  input      [0:0]    port_x1_3,
  output     [0:0]    port_y_0,
  output     [0:0]    port_y_1,
  output     [0:0]    port_y_2,
  output     [0:0]    port_y_3
);


  assign port_y_0[0] = (! (port_x0_0[0] ^ port_x1_0[0]));
  assign port_y_1[0] = (port_x0_1[0] ^ port_x1_1[0]);
  assign port_y_2[0] = (port_x0_2[0] ^ port_x1_2[0]);
  assign port_y_3[0] = (port_x0_3[0] ^ port_x1_3[0]);

endmodule

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

module Multiplication_TI_noReg (
  input      [0:0]    port_x0_0,
  input      [0:0]    port_x0_1,
  input      [0:0]    port_x0_2,
  input      [0:0]    port_x0_3,
  input      [0:0]    port_x1_0,
  input      [0:0]    port_x1_1,
  input      [0:0]    port_x1_2,
  input      [0:0]    port_x1_3,
  output     [0:0]    port_y_0,
  output     [0:0]    port_y_1,
  output     [0:0]    port_y_2,
  output     [0:0]    port_y_3
);

  wire       [0:0]    _zz_port_y_0;
  wire       [0:0]    _zz_port_y_1;
  wire       [0:0]    _zz_port_y_2;
  wire       [0:0]    _zz_port_y_3;

  assign _zz_port_y_0[0] = (((((port_x0_1[0] ^ port_x0_2[0]) ^ port_x0_3[0]) && (port_x1_1[0] ^ port_x1_2[0])) ^ port_x1_3[0]) ^ port_x1_2[0]);
  assign _zz_port_y_1[0] = ((((port_x0_0[0] ^ port_x0_2[0]) && (port_x1_0[0] ^ port_x1_3[0])) ^ (port_x0_0[0] && port_x1_2[0])) ^ port_x0_3[0]);
  assign _zz_port_y_2[0] = ((((port_x0_1[0] ^ port_x0_3[0]) && (port_x1_0[0] ^ port_x1_3[0])) ^ port_x0_3[0]) ^ port_x1_3[0]);
  assign _zz_port_y_3[0] = ((port_x0_0[0] && port_x1_1[0]) ^ port_x1_2[0]);
  assign port_y_0 = _zz_port_y_0;
  assign port_y_1 = _zz_port_y_1;
  assign port_y_2 = _zz_port_y_2;
  assign port_y_3 = _zz_port_y_3;

endmodule

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

module Multiplication_TI (
  input      [0:0]    port_x0_0,
  input      [0:0]    port_x0_1,
  input      [0:0]    port_x0_2,
  input      [0:0]    port_x0_3,
  input      [0:0]    port_x1_0,
  input      [0:0]    port_x1_1,
  input      [0:0]    port_x1_2,
  input      [0:0]    port_x1_3,
  output     [0:0]    port_y_0,
  output     [0:0]    port_y_1,
  output     [0:0]    port_y_2,
  output     [0:0]    port_y_3,
  input               clk,
  input               reset
);

  wire       [0:0]    _zz_port_y_0;
  wire       [0:0]    _zz_port_y_1;
  wire       [0:0]    _zz_port_y_2;
  wire       [0:0]    _zz_port_y_3;
  reg        [0:0]    _zz_port_y_0_1;
  reg        [0:0]    _zz_port_y_1_1;
  reg        [0:0]    _zz_port_y_2_1;
  reg        [0:0]    _zz_port_y_3_1;

  assign _zz_port_y_0[0] = (((((port_x0_1[0] ^ port_x0_2[0]) ^ port_x0_3[0]) && (port_x1_1[0] ^ port_x1_2[0])) ^ port_x1_3[0]) ^ port_x1_2[0]);
  assign _zz_port_y_1[0] = ((((port_x0_0[0] ^ port_x0_2[0]) && (port_x1_0[0] ^ port_x1_3[0])) ^ (port_x0_0[0] && port_x1_2[0])) ^ port_x0_3[0]);
  assign _zz_port_y_2[0] = ((((port_x0_1[0] ^ port_x0_3[0]) && (port_x1_0[0] ^ port_x1_3[0])) ^ port_x0_3[0]) ^ port_x1_3[0]);
  assign _zz_port_y_3[0] = ((port_x0_0[0] && port_x1_1[0]) ^ port_x1_2[0]);
  assign port_y_0 = _zz_port_y_0_1;
  assign port_y_1 = _zz_port_y_1_1;
  assign port_y_2 = _zz_port_y_2_1;
  assign port_y_3 = _zz_port_y_3_1;
  always @(posedge clk) begin
    _zz_port_y_0_1 <= _zz_port_y_0;
    _zz_port_y_1_1 <= _zz_port_y_1;
    _zz_port_y_2_1 <= _zz_port_y_2;
    _zz_port_y_3_1 <= _zz_port_y_3;
  end


endmodule

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

module Addition_TI (
  input      [0:0]    port_x0_0,
  input      [0:0]    port_x0_1,
  input      [0:0]    port_x0_2,
  input      [0:0]    port_x0_3,
  input      [0:0]    port_x1_0,
  input      [0:0]    port_x1_1,
  input      [0:0]    port_x1_2,
  input      [0:0]    port_x1_3,
  output     [0:0]    port_y_0,
  output     [0:0]    port_y_1,
  output     [0:0]    port_y_2,
  output     [0:0]    port_y_3
);


  assign port_y_0[0] = (port_x0_0[0] ^ port_x1_0[0]);
  assign port_y_1[0] = (port_x0_1[0] ^ port_x1_1[0]);
  assign port_y_2[0] = (port_x0_2[0] ^ port_x1_2[0]);
  assign port_y_3[0] = (port_x0_3[0] ^ port_x1_3[0]);

endmodule
