// Generator : SpinalHDL v1.7.3    git head : aeaeece704fe43c766e0d36a93f2ecbb8a9f2003
// Component : AES_Round
// Git hash  : db593c14fe8e83f0a4a5d43cf13325e631d65148

`timescale 1ns/1ps

module Round_AES_CMS_d1 (
  input      [0:0]    port_state_in_0_0_0,
  input      [0:0]    port_state_in_0_0_1,
  input      [0:0]    port_state_in_0_0_2,
  input      [0:0]    port_state_in_0_0_3,
  input      [0:0]    port_state_in_0_0_4,
  input      [0:0]    port_state_in_0_0_5,
  input      [0:0]    port_state_in_0_0_6,
  input      [0:0]    port_state_in_0_0_7,
  input      [0:0]    port_state_in_0_1_0,
  input      [0:0]    port_state_in_0_1_1,
  input      [0:0]    port_state_in_0_1_2,
  input      [0:0]    port_state_in_0_1_3,
  input      [0:0]    port_state_in_0_1_4,
  input      [0:0]    port_state_in_0_1_5,
  input      [0:0]    port_state_in_0_1_6,
  input      [0:0]    port_state_in_0_1_7,
  input      [0:0]    port_state_in_1_0_0,
  input      [0:0]    port_state_in_1_0_1,
  input      [0:0]    port_state_in_1_0_2,
  input      [0:0]    port_state_in_1_0_3,
  input      [0:0]    port_state_in_1_0_4,
  input      [0:0]    port_state_in_1_0_5,
  input      [0:0]    port_state_in_1_0_6,
  input      [0:0]    port_state_in_1_0_7,
  input      [0:0]    port_state_in_1_1_0,
  input      [0:0]    port_state_in_1_1_1,
  input      [0:0]    port_state_in_1_1_2,
  input      [0:0]    port_state_in_1_1_3,
  input      [0:0]    port_state_in_1_1_4,
  input      [0:0]    port_state_in_1_1_5,
  input      [0:0]    port_state_in_1_1_6,
  input      [0:0]    port_state_in_1_1_7,
  input      [0:0]    port_state_in_2_0_0,
  input      [0:0]    port_state_in_2_0_1,
  input      [0:0]    port_state_in_2_0_2,
  input      [0:0]    port_state_in_2_0_3,
  input      [0:0]    port_state_in_2_0_4,
  input      [0:0]    port_state_in_2_0_5,
  input      [0:0]    port_state_in_2_0_6,
  input      [0:0]    port_state_in_2_0_7,
  input      [0:0]    port_state_in_2_1_0,
  input      [0:0]    port_state_in_2_1_1,
  input      [0:0]    port_state_in_2_1_2,
  input      [0:0]    port_state_in_2_1_3,
  input      [0:0]    port_state_in_2_1_4,
  input      [0:0]    port_state_in_2_1_5,
  input      [0:0]    port_state_in_2_1_6,
  input      [0:0]    port_state_in_2_1_7,
  input      [0:0]    port_state_in_3_0_0,
  input      [0:0]    port_state_in_3_0_1,
  input      [0:0]    port_state_in_3_0_2,
  input      [0:0]    port_state_in_3_0_3,
  input      [0:0]    port_state_in_3_0_4,
  input      [0:0]    port_state_in_3_0_5,
  input      [0:0]    port_state_in_3_0_6,
  input      [0:0]    port_state_in_3_0_7,
  input      [0:0]    port_state_in_3_1_0,
  input      [0:0]    port_state_in_3_1_1,
  input      [0:0]    port_state_in_3_1_2,
  input      [0:0]    port_state_in_3_1_3,
  input      [0:0]    port_state_in_3_1_4,
  input      [0:0]    port_state_in_3_1_5,
  input      [0:0]    port_state_in_3_1_6,
  input      [0:0]    port_state_in_3_1_7,
  input      [0:0]    port_state_in_4_0_0,
  input      [0:0]    port_state_in_4_0_1,
  input      [0:0]    port_state_in_4_0_2,
  input      [0:0]    port_state_in_4_0_3,
  input      [0:0]    port_state_in_4_0_4,
  input      [0:0]    port_state_in_4_0_5,
  input      [0:0]    port_state_in_4_0_6,
  input      [0:0]    port_state_in_4_0_7,
  input      [0:0]    port_state_in_4_1_0,
  input      [0:0]    port_state_in_4_1_1,
  input      [0:0]    port_state_in_4_1_2,
  input      [0:0]    port_state_in_4_1_3,
  input      [0:0]    port_state_in_4_1_4,
  input      [0:0]    port_state_in_4_1_5,
  input      [0:0]    port_state_in_4_1_6,
  input      [0:0]    port_state_in_4_1_7,
  input      [0:0]    port_state_in_5_0_0,
  input      [0:0]    port_state_in_5_0_1,
  input      [0:0]    port_state_in_5_0_2,
  input      [0:0]    port_state_in_5_0_3,
  input      [0:0]    port_state_in_5_0_4,
  input      [0:0]    port_state_in_5_0_5,
  input      [0:0]    port_state_in_5_0_6,
  input      [0:0]    port_state_in_5_0_7,
  input      [0:0]    port_state_in_5_1_0,
  input      [0:0]    port_state_in_5_1_1,
  input      [0:0]    port_state_in_5_1_2,
  input      [0:0]    port_state_in_5_1_3,
  input      [0:0]    port_state_in_5_1_4,
  input      [0:0]    port_state_in_5_1_5,
  input      [0:0]    port_state_in_5_1_6,
  input      [0:0]    port_state_in_5_1_7,
  input      [0:0]    port_state_in_6_0_0,
  input      [0:0]    port_state_in_6_0_1,
  input      [0:0]    port_state_in_6_0_2,
  input      [0:0]    port_state_in_6_0_3,
  input      [0:0]    port_state_in_6_0_4,
  input      [0:0]    port_state_in_6_0_5,
  input      [0:0]    port_state_in_6_0_6,
  input      [0:0]    port_state_in_6_0_7,
  input      [0:0]    port_state_in_6_1_0,
  input      [0:0]    port_state_in_6_1_1,
  input      [0:0]    port_state_in_6_1_2,
  input      [0:0]    port_state_in_6_1_3,
  input      [0:0]    port_state_in_6_1_4,
  input      [0:0]    port_state_in_6_1_5,
  input      [0:0]    port_state_in_6_1_6,
  input      [0:0]    port_state_in_6_1_7,
  input      [0:0]    port_state_in_7_0_0,
  input      [0:0]    port_state_in_7_0_1,
  input      [0:0]    port_state_in_7_0_2,
  input      [0:0]    port_state_in_7_0_3,
  input      [0:0]    port_state_in_7_0_4,
  input      [0:0]    port_state_in_7_0_5,
  input      [0:0]    port_state_in_7_0_6,
  input      [0:0]    port_state_in_7_0_7,
  input      [0:0]    port_state_in_7_1_0,
  input      [0:0]    port_state_in_7_1_1,
  input      [0:0]    port_state_in_7_1_2,
  input      [0:0]    port_state_in_7_1_3,
  input      [0:0]    port_state_in_7_1_4,
  input      [0:0]    port_state_in_7_1_5,
  input      [0:0]    port_state_in_7_1_6,
  input      [0:0]    port_state_in_7_1_7,
  input      [0:0]    port_state_in_8_0_0,
  input      [0:0]    port_state_in_8_0_1,
  input      [0:0]    port_state_in_8_0_2,
  input      [0:0]    port_state_in_8_0_3,
  input      [0:0]    port_state_in_8_0_4,
  input      [0:0]    port_state_in_8_0_5,
  input      [0:0]    port_state_in_8_0_6,
  input      [0:0]    port_state_in_8_0_7,
  input      [0:0]    port_state_in_8_1_0,
  input      [0:0]    port_state_in_8_1_1,
  input      [0:0]    port_state_in_8_1_2,
  input      [0:0]    port_state_in_8_1_3,
  input      [0:0]    port_state_in_8_1_4,
  input      [0:0]    port_state_in_8_1_5,
  input      [0:0]    port_state_in_8_1_6,
  input      [0:0]    port_state_in_8_1_7,
  input      [0:0]    port_state_in_9_0_0,
  input      [0:0]    port_state_in_9_0_1,
  input      [0:0]    port_state_in_9_0_2,
  input      [0:0]    port_state_in_9_0_3,
  input      [0:0]    port_state_in_9_0_4,
  input      [0:0]    port_state_in_9_0_5,
  input      [0:0]    port_state_in_9_0_6,
  input      [0:0]    port_state_in_9_0_7,
  input      [0:0]    port_state_in_9_1_0,
  input      [0:0]    port_state_in_9_1_1,
  input      [0:0]    port_state_in_9_1_2,
  input      [0:0]    port_state_in_9_1_3,
  input      [0:0]    port_state_in_9_1_4,
  input      [0:0]    port_state_in_9_1_5,
  input      [0:0]    port_state_in_9_1_6,
  input      [0:0]    port_state_in_9_1_7,
  input      [0:0]    port_state_in_10_0_0,
  input      [0:0]    port_state_in_10_0_1,
  input      [0:0]    port_state_in_10_0_2,
  input      [0:0]    port_state_in_10_0_3,
  input      [0:0]    port_state_in_10_0_4,
  input      [0:0]    port_state_in_10_0_5,
  input      [0:0]    port_state_in_10_0_6,
  input      [0:0]    port_state_in_10_0_7,
  input      [0:0]    port_state_in_10_1_0,
  input      [0:0]    port_state_in_10_1_1,
  input      [0:0]    port_state_in_10_1_2,
  input      [0:0]    port_state_in_10_1_3,
  input      [0:0]    port_state_in_10_1_4,
  input      [0:0]    port_state_in_10_1_5,
  input      [0:0]    port_state_in_10_1_6,
  input      [0:0]    port_state_in_10_1_7,
  input      [0:0]    port_state_in_11_0_0,
  input      [0:0]    port_state_in_11_0_1,
  input      [0:0]    port_state_in_11_0_2,
  input      [0:0]    port_state_in_11_0_3,
  input      [0:0]    port_state_in_11_0_4,
  input      [0:0]    port_state_in_11_0_5,
  input      [0:0]    port_state_in_11_0_6,
  input      [0:0]    port_state_in_11_0_7,
  input      [0:0]    port_state_in_11_1_0,
  input      [0:0]    port_state_in_11_1_1,
  input      [0:0]    port_state_in_11_1_2,
  input      [0:0]    port_state_in_11_1_3,
  input      [0:0]    port_state_in_11_1_4,
  input      [0:0]    port_state_in_11_1_5,
  input      [0:0]    port_state_in_11_1_6,
  input      [0:0]    port_state_in_11_1_7,
  input      [0:0]    port_state_in_12_0_0,
  input      [0:0]    port_state_in_12_0_1,
  input      [0:0]    port_state_in_12_0_2,
  input      [0:0]    port_state_in_12_0_3,
  input      [0:0]    port_state_in_12_0_4,
  input      [0:0]    port_state_in_12_0_5,
  input      [0:0]    port_state_in_12_0_6,
  input      [0:0]    port_state_in_12_0_7,
  input      [0:0]    port_state_in_12_1_0,
  input      [0:0]    port_state_in_12_1_1,
  input      [0:0]    port_state_in_12_1_2,
  input      [0:0]    port_state_in_12_1_3,
  input      [0:0]    port_state_in_12_1_4,
  input      [0:0]    port_state_in_12_1_5,
  input      [0:0]    port_state_in_12_1_6,
  input      [0:0]    port_state_in_12_1_7,
  input      [0:0]    port_state_in_13_0_0,
  input      [0:0]    port_state_in_13_0_1,
  input      [0:0]    port_state_in_13_0_2,
  input      [0:0]    port_state_in_13_0_3,
  input      [0:0]    port_state_in_13_0_4,
  input      [0:0]    port_state_in_13_0_5,
  input      [0:0]    port_state_in_13_0_6,
  input      [0:0]    port_state_in_13_0_7,
  input      [0:0]    port_state_in_13_1_0,
  input      [0:0]    port_state_in_13_1_1,
  input      [0:0]    port_state_in_13_1_2,
  input      [0:0]    port_state_in_13_1_3,
  input      [0:0]    port_state_in_13_1_4,
  input      [0:0]    port_state_in_13_1_5,
  input      [0:0]    port_state_in_13_1_6,
  input      [0:0]    port_state_in_13_1_7,
  input      [0:0]    port_state_in_14_0_0,
  input      [0:0]    port_state_in_14_0_1,
  input      [0:0]    port_state_in_14_0_2,
  input      [0:0]    port_state_in_14_0_3,
  input      [0:0]    port_state_in_14_0_4,
  input      [0:0]    port_state_in_14_0_5,
  input      [0:0]    port_state_in_14_0_6,
  input      [0:0]    port_state_in_14_0_7,
  input      [0:0]    port_state_in_14_1_0,
  input      [0:0]    port_state_in_14_1_1,
  input      [0:0]    port_state_in_14_1_2,
  input      [0:0]    port_state_in_14_1_3,
  input      [0:0]    port_state_in_14_1_4,
  input      [0:0]    port_state_in_14_1_5,
  input      [0:0]    port_state_in_14_1_6,
  input      [0:0]    port_state_in_14_1_7,
  input      [0:0]    port_state_in_15_0_0,
  input      [0:0]    port_state_in_15_0_1,
  input      [0:0]    port_state_in_15_0_2,
  input      [0:0]    port_state_in_15_0_3,
  input      [0:0]    port_state_in_15_0_4,
  input      [0:0]    port_state_in_15_0_5,
  input      [0:0]    port_state_in_15_0_6,
  input      [0:0]    port_state_in_15_0_7,
  input      [0:0]    port_state_in_15_1_0,
  input      [0:0]    port_state_in_15_1_1,
  input      [0:0]    port_state_in_15_1_2,
  input      [0:0]    port_state_in_15_1_3,
  input      [0:0]    port_state_in_15_1_4,
  input      [0:0]    port_state_in_15_1_5,
  input      [0:0]    port_state_in_15_1_6,
  input      [0:0]    port_state_in_15_1_7,
  input      [0:0]    port_key_0_0_0,
  input      [0:0]    port_key_0_0_1,
  input      [0:0]    port_key_0_0_2,
  input      [0:0]    port_key_0_0_3,
  input      [0:0]    port_key_0_0_4,
  input      [0:0]    port_key_0_0_5,
  input      [0:0]    port_key_0_0_6,
  input      [0:0]    port_key_0_0_7,
  input      [0:0]    port_key_0_1_0,
  input      [0:0]    port_key_0_1_1,
  input      [0:0]    port_key_0_1_2,
  input      [0:0]    port_key_0_1_3,
  input      [0:0]    port_key_0_1_4,
  input      [0:0]    port_key_0_1_5,
  input      [0:0]    port_key_0_1_6,
  input      [0:0]    port_key_0_1_7,
  input      [0:0]    port_key_1_0_0,
  input      [0:0]    port_key_1_0_1,
  input      [0:0]    port_key_1_0_2,
  input      [0:0]    port_key_1_0_3,
  input      [0:0]    port_key_1_0_4,
  input      [0:0]    port_key_1_0_5,
  input      [0:0]    port_key_1_0_6,
  input      [0:0]    port_key_1_0_7,
  input      [0:0]    port_key_1_1_0,
  input      [0:0]    port_key_1_1_1,
  input      [0:0]    port_key_1_1_2,
  input      [0:0]    port_key_1_1_3,
  input      [0:0]    port_key_1_1_4,
  input      [0:0]    port_key_1_1_5,
  input      [0:0]    port_key_1_1_6,
  input      [0:0]    port_key_1_1_7,
  input      [0:0]    port_key_2_0_0,
  input      [0:0]    port_key_2_0_1,
  input      [0:0]    port_key_2_0_2,
  input      [0:0]    port_key_2_0_3,
  input      [0:0]    port_key_2_0_4,
  input      [0:0]    port_key_2_0_5,
  input      [0:0]    port_key_2_0_6,
  input      [0:0]    port_key_2_0_7,
  input      [0:0]    port_key_2_1_0,
  input      [0:0]    port_key_2_1_1,
  input      [0:0]    port_key_2_1_2,
  input      [0:0]    port_key_2_1_3,
  input      [0:0]    port_key_2_1_4,
  input      [0:0]    port_key_2_1_5,
  input      [0:0]    port_key_2_1_6,
  input      [0:0]    port_key_2_1_7,
  input      [0:0]    port_key_3_0_0,
  input      [0:0]    port_key_3_0_1,
  input      [0:0]    port_key_3_0_2,
  input      [0:0]    port_key_3_0_3,
  input      [0:0]    port_key_3_0_4,
  input      [0:0]    port_key_3_0_5,
  input      [0:0]    port_key_3_0_6,
  input      [0:0]    port_key_3_0_7,
  input      [0:0]    port_key_3_1_0,
  input      [0:0]    port_key_3_1_1,
  input      [0:0]    port_key_3_1_2,
  input      [0:0]    port_key_3_1_3,
  input      [0:0]    port_key_3_1_4,
  input      [0:0]    port_key_3_1_5,
  input      [0:0]    port_key_3_1_6,
  input      [0:0]    port_key_3_1_7,
  input      [0:0]    port_key_4_0_0,
  input      [0:0]    port_key_4_0_1,
  input      [0:0]    port_key_4_0_2,
  input      [0:0]    port_key_4_0_3,
  input      [0:0]    port_key_4_0_4,
  input      [0:0]    port_key_4_0_5,
  input      [0:0]    port_key_4_0_6,
  input      [0:0]    port_key_4_0_7,
  input      [0:0]    port_key_4_1_0,
  input      [0:0]    port_key_4_1_1,
  input      [0:0]    port_key_4_1_2,
  input      [0:0]    port_key_4_1_3,
  input      [0:0]    port_key_4_1_4,
  input      [0:0]    port_key_4_1_5,
  input      [0:0]    port_key_4_1_6,
  input      [0:0]    port_key_4_1_7,
  input      [0:0]    port_key_5_0_0,
  input      [0:0]    port_key_5_0_1,
  input      [0:0]    port_key_5_0_2,
  input      [0:0]    port_key_5_0_3,
  input      [0:0]    port_key_5_0_4,
  input      [0:0]    port_key_5_0_5,
  input      [0:0]    port_key_5_0_6,
  input      [0:0]    port_key_5_0_7,
  input      [0:0]    port_key_5_1_0,
  input      [0:0]    port_key_5_1_1,
  input      [0:0]    port_key_5_1_2,
  input      [0:0]    port_key_5_1_3,
  input      [0:0]    port_key_5_1_4,
  input      [0:0]    port_key_5_1_5,
  input      [0:0]    port_key_5_1_6,
  input      [0:0]    port_key_5_1_7,
  input      [0:0]    port_key_6_0_0,
  input      [0:0]    port_key_6_0_1,
  input      [0:0]    port_key_6_0_2,
  input      [0:0]    port_key_6_0_3,
  input      [0:0]    port_key_6_0_4,
  input      [0:0]    port_key_6_0_5,
  input      [0:0]    port_key_6_0_6,
  input      [0:0]    port_key_6_0_7,
  input      [0:0]    port_key_6_1_0,
  input      [0:0]    port_key_6_1_1,
  input      [0:0]    port_key_6_1_2,
  input      [0:0]    port_key_6_1_3,
  input      [0:0]    port_key_6_1_4,
  input      [0:0]    port_key_6_1_5,
  input      [0:0]    port_key_6_1_6,
  input      [0:0]    port_key_6_1_7,
  input      [0:0]    port_key_7_0_0,
  input      [0:0]    port_key_7_0_1,
  input      [0:0]    port_key_7_0_2,
  input      [0:0]    port_key_7_0_3,
  input      [0:0]    port_key_7_0_4,
  input      [0:0]    port_key_7_0_5,
  input      [0:0]    port_key_7_0_6,
  input      [0:0]    port_key_7_0_7,
  input      [0:0]    port_key_7_1_0,
  input      [0:0]    port_key_7_1_1,
  input      [0:0]    port_key_7_1_2,
  input      [0:0]    port_key_7_1_3,
  input      [0:0]    port_key_7_1_4,
  input      [0:0]    port_key_7_1_5,
  input      [0:0]    port_key_7_1_6,
  input      [0:0]    port_key_7_1_7,
  input      [0:0]    port_key_8_0_0,
  input      [0:0]    port_key_8_0_1,
  input      [0:0]    port_key_8_0_2,
  input      [0:0]    port_key_8_0_3,
  input      [0:0]    port_key_8_0_4,
  input      [0:0]    port_key_8_0_5,
  input      [0:0]    port_key_8_0_6,
  input      [0:0]    port_key_8_0_7,
  input      [0:0]    port_key_8_1_0,
  input      [0:0]    port_key_8_1_1,
  input      [0:0]    port_key_8_1_2,
  input      [0:0]    port_key_8_1_3,
  input      [0:0]    port_key_8_1_4,
  input      [0:0]    port_key_8_1_5,
  input      [0:0]    port_key_8_1_6,
  input      [0:0]    port_key_8_1_7,
  input      [0:0]    port_key_9_0_0,
  input      [0:0]    port_key_9_0_1,
  input      [0:0]    port_key_9_0_2,
  input      [0:0]    port_key_9_0_3,
  input      [0:0]    port_key_9_0_4,
  input      [0:0]    port_key_9_0_5,
  input      [0:0]    port_key_9_0_6,
  input      [0:0]    port_key_9_0_7,
  input      [0:0]    port_key_9_1_0,
  input      [0:0]    port_key_9_1_1,
  input      [0:0]    port_key_9_1_2,
  input      [0:0]    port_key_9_1_3,
  input      [0:0]    port_key_9_1_4,
  input      [0:0]    port_key_9_1_5,
  input      [0:0]    port_key_9_1_6,
  input      [0:0]    port_key_9_1_7,
  input      [0:0]    port_key_10_0_0,
  input      [0:0]    port_key_10_0_1,
  input      [0:0]    port_key_10_0_2,
  input      [0:0]    port_key_10_0_3,
  input      [0:0]    port_key_10_0_4,
  input      [0:0]    port_key_10_0_5,
  input      [0:0]    port_key_10_0_6,
  input      [0:0]    port_key_10_0_7,
  input      [0:0]    port_key_10_1_0,
  input      [0:0]    port_key_10_1_1,
  input      [0:0]    port_key_10_1_2,
  input      [0:0]    port_key_10_1_3,
  input      [0:0]    port_key_10_1_4,
  input      [0:0]    port_key_10_1_5,
  input      [0:0]    port_key_10_1_6,
  input      [0:0]    port_key_10_1_7,
  input      [0:0]    port_key_11_0_0,
  input      [0:0]    port_key_11_0_1,
  input      [0:0]    port_key_11_0_2,
  input      [0:0]    port_key_11_0_3,
  input      [0:0]    port_key_11_0_4,
  input      [0:0]    port_key_11_0_5,
  input      [0:0]    port_key_11_0_6,
  input      [0:0]    port_key_11_0_7,
  input      [0:0]    port_key_11_1_0,
  input      [0:0]    port_key_11_1_1,
  input      [0:0]    port_key_11_1_2,
  input      [0:0]    port_key_11_1_3,
  input      [0:0]    port_key_11_1_4,
  input      [0:0]    port_key_11_1_5,
  input      [0:0]    port_key_11_1_6,
  input      [0:0]    port_key_11_1_7,
  input      [0:0]    port_key_12_0_0,
  input      [0:0]    port_key_12_0_1,
  input      [0:0]    port_key_12_0_2,
  input      [0:0]    port_key_12_0_3,
  input      [0:0]    port_key_12_0_4,
  input      [0:0]    port_key_12_0_5,
  input      [0:0]    port_key_12_0_6,
  input      [0:0]    port_key_12_0_7,
  input      [0:0]    port_key_12_1_0,
  input      [0:0]    port_key_12_1_1,
  input      [0:0]    port_key_12_1_2,
  input      [0:0]    port_key_12_1_3,
  input      [0:0]    port_key_12_1_4,
  input      [0:0]    port_key_12_1_5,
  input      [0:0]    port_key_12_1_6,
  input      [0:0]    port_key_12_1_7,
  input      [0:0]    port_key_13_0_0,
  input      [0:0]    port_key_13_0_1,
  input      [0:0]    port_key_13_0_2,
  input      [0:0]    port_key_13_0_3,
  input      [0:0]    port_key_13_0_4,
  input      [0:0]    port_key_13_0_5,
  input      [0:0]    port_key_13_0_6,
  input      [0:0]    port_key_13_0_7,
  input      [0:0]    port_key_13_1_0,
  input      [0:0]    port_key_13_1_1,
  input      [0:0]    port_key_13_1_2,
  input      [0:0]    port_key_13_1_3,
  input      [0:0]    port_key_13_1_4,
  input      [0:0]    port_key_13_1_5,
  input      [0:0]    port_key_13_1_6,
  input      [0:0]    port_key_13_1_7,
  input      [0:0]    port_key_14_0_0,
  input      [0:0]    port_key_14_0_1,
  input      [0:0]    port_key_14_0_2,
  input      [0:0]    port_key_14_0_3,
  input      [0:0]    port_key_14_0_4,
  input      [0:0]    port_key_14_0_5,
  input      [0:0]    port_key_14_0_6,
  input      [0:0]    port_key_14_0_7,
  input      [0:0]    port_key_14_1_0,
  input      [0:0]    port_key_14_1_1,
  input      [0:0]    port_key_14_1_2,
  input      [0:0]    port_key_14_1_3,
  input      [0:0]    port_key_14_1_4,
  input      [0:0]    port_key_14_1_5,
  input      [0:0]    port_key_14_1_6,
  input      [0:0]    port_key_14_1_7,
  input      [0:0]    port_key_15_0_0,
  input      [0:0]    port_key_15_0_1,
  input      [0:0]    port_key_15_0_2,
  input      [0:0]    port_key_15_0_3,
  input      [0:0]    port_key_15_0_4,
  input      [0:0]    port_key_15_0_5,
  input      [0:0]    port_key_15_0_6,
  input      [0:0]    port_key_15_0_7,
  input      [0:0]    port_key_15_1_0,
  input      [0:0]    port_key_15_1_1,
  input      [0:0]    port_key_15_1_2,
  input      [0:0]    port_key_15_1_3,
  input      [0:0]    port_key_15_1_4,
  input      [0:0]    port_key_15_1_5,
  input      [0:0]    port_key_15_1_6,
  input      [0:0]    port_key_15_1_7,
  input               port_rand_0_0,
  input               port_rand_0_1,
  input               port_rand_0_2,
  input               port_rand_0_3,
  input               port_rand_0_4,
  input               port_rand_0_5,
  input               port_rand_0_6,
  input               port_rand_0_7,
  input               port_rand_0_8,
  input               port_rand_0_9,
  input               port_rand_0_10,
  input               port_rand_0_11,
  input               port_rand_0_12,
  input               port_rand_0_13,
  input               port_rand_0_14,
  input               port_rand_0_15,
  input               port_rand_0_16,
  input               port_rand_0_17,
  input               port_rand_0_18,
  input               port_rand_0_19,
  input               port_rand_0_20,
  input               port_rand_0_21,
  input               port_rand_0_22,
  input               port_rand_0_23,
  input               port_rand_0_24,
  input               port_rand_0_25,
  input               port_rand_0_26,
  input               port_rand_0_27,
  input               port_rand_0_28,
  input               port_rand_0_29,
  input               port_rand_0_30,
  input               port_rand_0_31,
  input               port_rand_0_32,
  input               port_rand_0_33,
  input               port_rand_0_34,
  input               port_rand_0_35,
  input               port_rand_0_36,
  input               port_rand_0_37,
  input               port_rand_0_38,
  input               port_rand_0_39,
  input               port_rand_0_40,
  input               port_rand_0_41,
  input               port_rand_0_42,
  input               port_rand_0_43,
  input               port_rand_0_44,
  input               port_rand_0_45,
  input               port_rand_0_46,
  input               port_rand_0_47,
  input               port_rand_0_48,
  input               port_rand_0_49,
  input               port_rand_0_50,
  input               port_rand_0_51,
  input               port_rand_0_52,
  input               port_rand_0_53,
  input               port_rand_1_0,
  input               port_rand_1_1,
  input               port_rand_1_2,
  input               port_rand_1_3,
  input               port_rand_1_4,
  input               port_rand_1_5,
  input               port_rand_1_6,
  input               port_rand_1_7,
  input               port_rand_1_8,
  input               port_rand_1_9,
  input               port_rand_1_10,
  input               port_rand_1_11,
  input               port_rand_1_12,
  input               port_rand_1_13,
  input               port_rand_1_14,
  input               port_rand_1_15,
  input               port_rand_1_16,
  input               port_rand_1_17,
  input               port_rand_1_18,
  input               port_rand_1_19,
  input               port_rand_1_20,
  input               port_rand_1_21,
  input               port_rand_1_22,
  input               port_rand_1_23,
  input               port_rand_1_24,
  input               port_rand_1_25,
  input               port_rand_1_26,
  input               port_rand_1_27,
  input               port_rand_1_28,
  input               port_rand_1_29,
  input               port_rand_1_30,
  input               port_rand_1_31,
  input               port_rand_1_32,
  input               port_rand_1_33,
  input               port_rand_1_34,
  input               port_rand_1_35,
  input               port_rand_1_36,
  input               port_rand_1_37,
  input               port_rand_1_38,
  input               port_rand_1_39,
  input               port_rand_1_40,
  input               port_rand_1_41,
  input               port_rand_1_42,
  input               port_rand_1_43,
  input               port_rand_1_44,
  input               port_rand_1_45,
  input               port_rand_1_46,
  input               port_rand_1_47,
  input               port_rand_1_48,
  input               port_rand_1_49,
  input               port_rand_1_50,
  input               port_rand_1_51,
  input               port_rand_1_52,
  input               port_rand_1_53,
  input               port_rand_2_0,
  input               port_rand_2_1,
  input               port_rand_2_2,
  input               port_rand_2_3,
  input               port_rand_2_4,
  input               port_rand_2_5,
  input               port_rand_2_6,
  input               port_rand_2_7,
  input               port_rand_2_8,
  input               port_rand_2_9,
  input               port_rand_2_10,
  input               port_rand_2_11,
  input               port_rand_2_12,
  input               port_rand_2_13,
  input               port_rand_2_14,
  input               port_rand_2_15,
  input               port_rand_2_16,
  input               port_rand_2_17,
  input               port_rand_2_18,
  input               port_rand_2_19,
  input               port_rand_2_20,
  input               port_rand_2_21,
  input               port_rand_2_22,
  input               port_rand_2_23,
  input               port_rand_2_24,
  input               port_rand_2_25,
  input               port_rand_2_26,
  input               port_rand_2_27,
  input               port_rand_2_28,
  input               port_rand_2_29,
  input               port_rand_2_30,
  input               port_rand_2_31,
  input               port_rand_2_32,
  input               port_rand_2_33,
  input               port_rand_2_34,
  input               port_rand_2_35,
  input               port_rand_2_36,
  input               port_rand_2_37,
  input               port_rand_2_38,
  input               port_rand_2_39,
  input               port_rand_2_40,
  input               port_rand_2_41,
  input               port_rand_2_42,
  input               port_rand_2_43,
  input               port_rand_2_44,
  input               port_rand_2_45,
  input               port_rand_2_46,
  input               port_rand_2_47,
  input               port_rand_2_48,
  input               port_rand_2_49,
  input               port_rand_2_50,
  input               port_rand_2_51,
  input               port_rand_2_52,
  input               port_rand_2_53,
  input               port_rand_3_0,
  input               port_rand_3_1,
  input               port_rand_3_2,
  input               port_rand_3_3,
  input               port_rand_3_4,
  input               port_rand_3_5,
  input               port_rand_3_6,
  input               port_rand_3_7,
  input               port_rand_3_8,
  input               port_rand_3_9,
  input               port_rand_3_10,
  input               port_rand_3_11,
  input               port_rand_3_12,
  input               port_rand_3_13,
  input               port_rand_3_14,
  input               port_rand_3_15,
  input               port_rand_3_16,
  input               port_rand_3_17,
  input               port_rand_3_18,
  input               port_rand_3_19,
  input               port_rand_3_20,
  input               port_rand_3_21,
  input               port_rand_3_22,
  input               port_rand_3_23,
  input               port_rand_3_24,
  input               port_rand_3_25,
  input               port_rand_3_26,
  input               port_rand_3_27,
  input               port_rand_3_28,
  input               port_rand_3_29,
  input               port_rand_3_30,
  input               port_rand_3_31,
  input               port_rand_3_32,
  input               port_rand_3_33,
  input               port_rand_3_34,
  input               port_rand_3_35,
  input               port_rand_3_36,
  input               port_rand_3_37,
  input               port_rand_3_38,
  input               port_rand_3_39,
  input               port_rand_3_40,
  input               port_rand_3_41,
  input               port_rand_3_42,
  input               port_rand_3_43,
  input               port_rand_3_44,
  input               port_rand_3_45,
  input               port_rand_3_46,
  input               port_rand_3_47,
  input               port_rand_3_48,
  input               port_rand_3_49,
  input               port_rand_3_50,
  input               port_rand_3_51,
  input               port_rand_3_52,
  input               port_rand_3_53,
  input               port_rand_4_0,
  input               port_rand_4_1,
  input               port_rand_4_2,
  input               port_rand_4_3,
  input               port_rand_4_4,
  input               port_rand_4_5,
  input               port_rand_4_6,
  input               port_rand_4_7,
  input               port_rand_4_8,
  input               port_rand_4_9,
  input               port_rand_4_10,
  input               port_rand_4_11,
  input               port_rand_4_12,
  input               port_rand_4_13,
  input               port_rand_4_14,
  input               port_rand_4_15,
  input               port_rand_4_16,
  input               port_rand_4_17,
  input               port_rand_4_18,
  input               port_rand_4_19,
  input               port_rand_4_20,
  input               port_rand_4_21,
  input               port_rand_4_22,
  input               port_rand_4_23,
  input               port_rand_4_24,
  input               port_rand_4_25,
  input               port_rand_4_26,
  input               port_rand_4_27,
  input               port_rand_4_28,
  input               port_rand_4_29,
  input               port_rand_4_30,
  input               port_rand_4_31,
  input               port_rand_4_32,
  input               port_rand_4_33,
  input               port_rand_4_34,
  input               port_rand_4_35,
  input               port_rand_4_36,
  input               port_rand_4_37,
  input               port_rand_4_38,
  input               port_rand_4_39,
  input               port_rand_4_40,
  input               port_rand_4_41,
  input               port_rand_4_42,
  input               port_rand_4_43,
  input               port_rand_4_44,
  input               port_rand_4_45,
  input               port_rand_4_46,
  input               port_rand_4_47,
  input               port_rand_4_48,
  input               port_rand_4_49,
  input               port_rand_4_50,
  input               port_rand_4_51,
  input               port_rand_4_52,
  input               port_rand_4_53,
  input               port_rand_5_0,
  input               port_rand_5_1,
  input               port_rand_5_2,
  input               port_rand_5_3,
  input               port_rand_5_4,
  input               port_rand_5_5,
  input               port_rand_5_6,
  input               port_rand_5_7,
  input               port_rand_5_8,
  input               port_rand_5_9,
  input               port_rand_5_10,
  input               port_rand_5_11,
  input               port_rand_5_12,
  input               port_rand_5_13,
  input               port_rand_5_14,
  input               port_rand_5_15,
  input               port_rand_5_16,
  input               port_rand_5_17,
  input               port_rand_5_18,
  input               port_rand_5_19,
  input               port_rand_5_20,
  input               port_rand_5_21,
  input               port_rand_5_22,
  input               port_rand_5_23,
  input               port_rand_5_24,
  input               port_rand_5_25,
  input               port_rand_5_26,
  input               port_rand_5_27,
  input               port_rand_5_28,
  input               port_rand_5_29,
  input               port_rand_5_30,
  input               port_rand_5_31,
  input               port_rand_5_32,
  input               port_rand_5_33,
  input               port_rand_5_34,
  input               port_rand_5_35,
  input               port_rand_5_36,
  input               port_rand_5_37,
  input               port_rand_5_38,
  input               port_rand_5_39,
  input               port_rand_5_40,
  input               port_rand_5_41,
  input               port_rand_5_42,
  input               port_rand_5_43,
  input               port_rand_5_44,
  input               port_rand_5_45,
  input               port_rand_5_46,
  input               port_rand_5_47,
  input               port_rand_5_48,
  input               port_rand_5_49,
  input               port_rand_5_50,
  input               port_rand_5_51,
  input               port_rand_5_52,
  input               port_rand_5_53,
  input               port_rand_6_0,
  input               port_rand_6_1,
  input               port_rand_6_2,
  input               port_rand_6_3,
  input               port_rand_6_4,
  input               port_rand_6_5,
  input               port_rand_6_6,
  input               port_rand_6_7,
  input               port_rand_6_8,
  input               port_rand_6_9,
  input               port_rand_6_10,
  input               port_rand_6_11,
  input               port_rand_6_12,
  input               port_rand_6_13,
  input               port_rand_6_14,
  input               port_rand_6_15,
  input               port_rand_6_16,
  input               port_rand_6_17,
  input               port_rand_6_18,
  input               port_rand_6_19,
  input               port_rand_6_20,
  input               port_rand_6_21,
  input               port_rand_6_22,
  input               port_rand_6_23,
  input               port_rand_6_24,
  input               port_rand_6_25,
  input               port_rand_6_26,
  input               port_rand_6_27,
  input               port_rand_6_28,
  input               port_rand_6_29,
  input               port_rand_6_30,
  input               port_rand_6_31,
  input               port_rand_6_32,
  input               port_rand_6_33,
  input               port_rand_6_34,
  input               port_rand_6_35,
  input               port_rand_6_36,
  input               port_rand_6_37,
  input               port_rand_6_38,
  input               port_rand_6_39,
  input               port_rand_6_40,
  input               port_rand_6_41,
  input               port_rand_6_42,
  input               port_rand_6_43,
  input               port_rand_6_44,
  input               port_rand_6_45,
  input               port_rand_6_46,
  input               port_rand_6_47,
  input               port_rand_6_48,
  input               port_rand_6_49,
  input               port_rand_6_50,
  input               port_rand_6_51,
  input               port_rand_6_52,
  input               port_rand_6_53,
  input               port_rand_7_0,
  input               port_rand_7_1,
  input               port_rand_7_2,
  input               port_rand_7_3,
  input               port_rand_7_4,
  input               port_rand_7_5,
  input               port_rand_7_6,
  input               port_rand_7_7,
  input               port_rand_7_8,
  input               port_rand_7_9,
  input               port_rand_7_10,
  input               port_rand_7_11,
  input               port_rand_7_12,
  input               port_rand_7_13,
  input               port_rand_7_14,
  input               port_rand_7_15,
  input               port_rand_7_16,
  input               port_rand_7_17,
  input               port_rand_7_18,
  input               port_rand_7_19,
  input               port_rand_7_20,
  input               port_rand_7_21,
  input               port_rand_7_22,
  input               port_rand_7_23,
  input               port_rand_7_24,
  input               port_rand_7_25,
  input               port_rand_7_26,
  input               port_rand_7_27,
  input               port_rand_7_28,
  input               port_rand_7_29,
  input               port_rand_7_30,
  input               port_rand_7_31,
  input               port_rand_7_32,
  input               port_rand_7_33,
  input               port_rand_7_34,
  input               port_rand_7_35,
  input               port_rand_7_36,
  input               port_rand_7_37,
  input               port_rand_7_38,
  input               port_rand_7_39,
  input               port_rand_7_40,
  input               port_rand_7_41,
  input               port_rand_7_42,
  input               port_rand_7_43,
  input               port_rand_7_44,
  input               port_rand_7_45,
  input               port_rand_7_46,
  input               port_rand_7_47,
  input               port_rand_7_48,
  input               port_rand_7_49,
  input               port_rand_7_50,
  input               port_rand_7_51,
  input               port_rand_7_52,
  input               port_rand_7_53,
  input               port_rand_8_0,
  input               port_rand_8_1,
  input               port_rand_8_2,
  input               port_rand_8_3,
  input               port_rand_8_4,
  input               port_rand_8_5,
  input               port_rand_8_6,
  input               port_rand_8_7,
  input               port_rand_8_8,
  input               port_rand_8_9,
  input               port_rand_8_10,
  input               port_rand_8_11,
  input               port_rand_8_12,
  input               port_rand_8_13,
  input               port_rand_8_14,
  input               port_rand_8_15,
  input               port_rand_8_16,
  input               port_rand_8_17,
  input               port_rand_8_18,
  input               port_rand_8_19,
  input               port_rand_8_20,
  input               port_rand_8_21,
  input               port_rand_8_22,
  input               port_rand_8_23,
  input               port_rand_8_24,
  input               port_rand_8_25,
  input               port_rand_8_26,
  input               port_rand_8_27,
  input               port_rand_8_28,
  input               port_rand_8_29,
  input               port_rand_8_30,
  input               port_rand_8_31,
  input               port_rand_8_32,
  input               port_rand_8_33,
  input               port_rand_8_34,
  input               port_rand_8_35,
  input               port_rand_8_36,
  input               port_rand_8_37,
  input               port_rand_8_38,
  input               port_rand_8_39,
  input               port_rand_8_40,
  input               port_rand_8_41,
  input               port_rand_8_42,
  input               port_rand_8_43,
  input               port_rand_8_44,
  input               port_rand_8_45,
  input               port_rand_8_46,
  input               port_rand_8_47,
  input               port_rand_8_48,
  input               port_rand_8_49,
  input               port_rand_8_50,
  input               port_rand_8_51,
  input               port_rand_8_52,
  input               port_rand_8_53,
  input               port_rand_9_0,
  input               port_rand_9_1,
  input               port_rand_9_2,
  input               port_rand_9_3,
  input               port_rand_9_4,
  input               port_rand_9_5,
  input               port_rand_9_6,
  input               port_rand_9_7,
  input               port_rand_9_8,
  input               port_rand_9_9,
  input               port_rand_9_10,
  input               port_rand_9_11,
  input               port_rand_9_12,
  input               port_rand_9_13,
  input               port_rand_9_14,
  input               port_rand_9_15,
  input               port_rand_9_16,
  input               port_rand_9_17,
  input               port_rand_9_18,
  input               port_rand_9_19,
  input               port_rand_9_20,
  input               port_rand_9_21,
  input               port_rand_9_22,
  input               port_rand_9_23,
  input               port_rand_9_24,
  input               port_rand_9_25,
  input               port_rand_9_26,
  input               port_rand_9_27,
  input               port_rand_9_28,
  input               port_rand_9_29,
  input               port_rand_9_30,
  input               port_rand_9_31,
  input               port_rand_9_32,
  input               port_rand_9_33,
  input               port_rand_9_34,
  input               port_rand_9_35,
  input               port_rand_9_36,
  input               port_rand_9_37,
  input               port_rand_9_38,
  input               port_rand_9_39,
  input               port_rand_9_40,
  input               port_rand_9_41,
  input               port_rand_9_42,
  input               port_rand_9_43,
  input               port_rand_9_44,
  input               port_rand_9_45,
  input               port_rand_9_46,
  input               port_rand_9_47,
  input               port_rand_9_48,
  input               port_rand_9_49,
  input               port_rand_9_50,
  input               port_rand_9_51,
  input               port_rand_9_52,
  input               port_rand_9_53,
  input               port_rand_10_0,
  input               port_rand_10_1,
  input               port_rand_10_2,
  input               port_rand_10_3,
  input               port_rand_10_4,
  input               port_rand_10_5,
  input               port_rand_10_6,
  input               port_rand_10_7,
  input               port_rand_10_8,
  input               port_rand_10_9,
  input               port_rand_10_10,
  input               port_rand_10_11,
  input               port_rand_10_12,
  input               port_rand_10_13,
  input               port_rand_10_14,
  input               port_rand_10_15,
  input               port_rand_10_16,
  input               port_rand_10_17,
  input               port_rand_10_18,
  input               port_rand_10_19,
  input               port_rand_10_20,
  input               port_rand_10_21,
  input               port_rand_10_22,
  input               port_rand_10_23,
  input               port_rand_10_24,
  input               port_rand_10_25,
  input               port_rand_10_26,
  input               port_rand_10_27,
  input               port_rand_10_28,
  input               port_rand_10_29,
  input               port_rand_10_30,
  input               port_rand_10_31,
  input               port_rand_10_32,
  input               port_rand_10_33,
  input               port_rand_10_34,
  input               port_rand_10_35,
  input               port_rand_10_36,
  input               port_rand_10_37,
  input               port_rand_10_38,
  input               port_rand_10_39,
  input               port_rand_10_40,
  input               port_rand_10_41,
  input               port_rand_10_42,
  input               port_rand_10_43,
  input               port_rand_10_44,
  input               port_rand_10_45,
  input               port_rand_10_46,
  input               port_rand_10_47,
  input               port_rand_10_48,
  input               port_rand_10_49,
  input               port_rand_10_50,
  input               port_rand_10_51,
  input               port_rand_10_52,
  input               port_rand_10_53,
  input               port_rand_11_0,
  input               port_rand_11_1,
  input               port_rand_11_2,
  input               port_rand_11_3,
  input               port_rand_11_4,
  input               port_rand_11_5,
  input               port_rand_11_6,
  input               port_rand_11_7,
  input               port_rand_11_8,
  input               port_rand_11_9,
  input               port_rand_11_10,
  input               port_rand_11_11,
  input               port_rand_11_12,
  input               port_rand_11_13,
  input               port_rand_11_14,
  input               port_rand_11_15,
  input               port_rand_11_16,
  input               port_rand_11_17,
  input               port_rand_11_18,
  input               port_rand_11_19,
  input               port_rand_11_20,
  input               port_rand_11_21,
  input               port_rand_11_22,
  input               port_rand_11_23,
  input               port_rand_11_24,
  input               port_rand_11_25,
  input               port_rand_11_26,
  input               port_rand_11_27,
  input               port_rand_11_28,
  input               port_rand_11_29,
  input               port_rand_11_30,
  input               port_rand_11_31,
  input               port_rand_11_32,
  input               port_rand_11_33,
  input               port_rand_11_34,
  input               port_rand_11_35,
  input               port_rand_11_36,
  input               port_rand_11_37,
  input               port_rand_11_38,
  input               port_rand_11_39,
  input               port_rand_11_40,
  input               port_rand_11_41,
  input               port_rand_11_42,
  input               port_rand_11_43,
  input               port_rand_11_44,
  input               port_rand_11_45,
  input               port_rand_11_46,
  input               port_rand_11_47,
  input               port_rand_11_48,
  input               port_rand_11_49,
  input               port_rand_11_50,
  input               port_rand_11_51,
  input               port_rand_11_52,
  input               port_rand_11_53,
  input               port_rand_12_0,
  input               port_rand_12_1,
  input               port_rand_12_2,
  input               port_rand_12_3,
  input               port_rand_12_4,
  input               port_rand_12_5,
  input               port_rand_12_6,
  input               port_rand_12_7,
  input               port_rand_12_8,
  input               port_rand_12_9,
  input               port_rand_12_10,
  input               port_rand_12_11,
  input               port_rand_12_12,
  input               port_rand_12_13,
  input               port_rand_12_14,
  input               port_rand_12_15,
  input               port_rand_12_16,
  input               port_rand_12_17,
  input               port_rand_12_18,
  input               port_rand_12_19,
  input               port_rand_12_20,
  input               port_rand_12_21,
  input               port_rand_12_22,
  input               port_rand_12_23,
  input               port_rand_12_24,
  input               port_rand_12_25,
  input               port_rand_12_26,
  input               port_rand_12_27,
  input               port_rand_12_28,
  input               port_rand_12_29,
  input               port_rand_12_30,
  input               port_rand_12_31,
  input               port_rand_12_32,
  input               port_rand_12_33,
  input               port_rand_12_34,
  input               port_rand_12_35,
  input               port_rand_12_36,
  input               port_rand_12_37,
  input               port_rand_12_38,
  input               port_rand_12_39,
  input               port_rand_12_40,
  input               port_rand_12_41,
  input               port_rand_12_42,
  input               port_rand_12_43,
  input               port_rand_12_44,
  input               port_rand_12_45,
  input               port_rand_12_46,
  input               port_rand_12_47,
  input               port_rand_12_48,
  input               port_rand_12_49,
  input               port_rand_12_50,
  input               port_rand_12_51,
  input               port_rand_12_52,
  input               port_rand_12_53,
  input               port_rand_13_0,
  input               port_rand_13_1,
  input               port_rand_13_2,
  input               port_rand_13_3,
  input               port_rand_13_4,
  input               port_rand_13_5,
  input               port_rand_13_6,
  input               port_rand_13_7,
  input               port_rand_13_8,
  input               port_rand_13_9,
  input               port_rand_13_10,
  input               port_rand_13_11,
  input               port_rand_13_12,
  input               port_rand_13_13,
  input               port_rand_13_14,
  input               port_rand_13_15,
  input               port_rand_13_16,
  input               port_rand_13_17,
  input               port_rand_13_18,
  input               port_rand_13_19,
  input               port_rand_13_20,
  input               port_rand_13_21,
  input               port_rand_13_22,
  input               port_rand_13_23,
  input               port_rand_13_24,
  input               port_rand_13_25,
  input               port_rand_13_26,
  input               port_rand_13_27,
  input               port_rand_13_28,
  input               port_rand_13_29,
  input               port_rand_13_30,
  input               port_rand_13_31,
  input               port_rand_13_32,
  input               port_rand_13_33,
  input               port_rand_13_34,
  input               port_rand_13_35,
  input               port_rand_13_36,
  input               port_rand_13_37,
  input               port_rand_13_38,
  input               port_rand_13_39,
  input               port_rand_13_40,
  input               port_rand_13_41,
  input               port_rand_13_42,
  input               port_rand_13_43,
  input               port_rand_13_44,
  input               port_rand_13_45,
  input               port_rand_13_46,
  input               port_rand_13_47,
  input               port_rand_13_48,
  input               port_rand_13_49,
  input               port_rand_13_50,
  input               port_rand_13_51,
  input               port_rand_13_52,
  input               port_rand_13_53,
  input               port_rand_14_0,
  input               port_rand_14_1,
  input               port_rand_14_2,
  input               port_rand_14_3,
  input               port_rand_14_4,
  input               port_rand_14_5,
  input               port_rand_14_6,
  input               port_rand_14_7,
  input               port_rand_14_8,
  input               port_rand_14_9,
  input               port_rand_14_10,
  input               port_rand_14_11,
  input               port_rand_14_12,
  input               port_rand_14_13,
  input               port_rand_14_14,
  input               port_rand_14_15,
  input               port_rand_14_16,
  input               port_rand_14_17,
  input               port_rand_14_18,
  input               port_rand_14_19,
  input               port_rand_14_20,
  input               port_rand_14_21,
  input               port_rand_14_22,
  input               port_rand_14_23,
  input               port_rand_14_24,
  input               port_rand_14_25,
  input               port_rand_14_26,
  input               port_rand_14_27,
  input               port_rand_14_28,
  input               port_rand_14_29,
  input               port_rand_14_30,
  input               port_rand_14_31,
  input               port_rand_14_32,
  input               port_rand_14_33,
  input               port_rand_14_34,
  input               port_rand_14_35,
  input               port_rand_14_36,
  input               port_rand_14_37,
  input               port_rand_14_38,
  input               port_rand_14_39,
  input               port_rand_14_40,
  input               port_rand_14_41,
  input               port_rand_14_42,
  input               port_rand_14_43,
  input               port_rand_14_44,
  input               port_rand_14_45,
  input               port_rand_14_46,
  input               port_rand_14_47,
  input               port_rand_14_48,
  input               port_rand_14_49,
  input               port_rand_14_50,
  input               port_rand_14_51,
  input               port_rand_14_52,
  input               port_rand_14_53,
  input               port_rand_15_0,
  input               port_rand_15_1,
  input               port_rand_15_2,
  input               port_rand_15_3,
  input               port_rand_15_4,
  input               port_rand_15_5,
  input               port_rand_15_6,
  input               port_rand_15_7,
  input               port_rand_15_8,
  input               port_rand_15_9,
  input               port_rand_15_10,
  input               port_rand_15_11,
  input               port_rand_15_12,
  input               port_rand_15_13,
  input               port_rand_15_14,
  input               port_rand_15_15,
  input               port_rand_15_16,
  input               port_rand_15_17,
  input               port_rand_15_18,
  input               port_rand_15_19,
  input               port_rand_15_20,
  input               port_rand_15_21,
  input               port_rand_15_22,
  input               port_rand_15_23,
  input               port_rand_15_24,
  input               port_rand_15_25,
  input               port_rand_15_26,
  input               port_rand_15_27,
  input               port_rand_15_28,
  input               port_rand_15_29,
  input               port_rand_15_30,
  input               port_rand_15_31,
  input               port_rand_15_32,
  input               port_rand_15_33,
  input               port_rand_15_34,
  input               port_rand_15_35,
  input               port_rand_15_36,
  input               port_rand_15_37,
  input               port_rand_15_38,
  input               port_rand_15_39,
  input               port_rand_15_40,
  input               port_rand_15_41,
  input               port_rand_15_42,
  input               port_rand_15_43,
  input               port_rand_15_44,
  input               port_rand_15_45,
  input               port_rand_15_46,
  input               port_rand_15_47,
  input               port_rand_15_48,
  input               port_rand_15_49,
  input               port_rand_15_50,
  input               port_rand_15_51,
  input               port_rand_15_52,
  input               port_rand_15_53,
  output     [0:0]    port_state_out_0_0_0,
  output     [0:0]    port_state_out_0_0_1,
  output     [0:0]    port_state_out_0_0_2,
  output     [0:0]    port_state_out_0_0_3,
  output     [0:0]    port_state_out_0_0_4,
  output     [0:0]    port_state_out_0_0_5,
  output     [0:0]    port_state_out_0_0_6,
  output     [0:0]    port_state_out_0_0_7,
  output     [0:0]    port_state_out_0_1_0,
  output     [0:0]    port_state_out_0_1_1,
  output     [0:0]    port_state_out_0_1_2,
  output     [0:0]    port_state_out_0_1_3,
  output     [0:0]    port_state_out_0_1_4,
  output     [0:0]    port_state_out_0_1_5,
  output     [0:0]    port_state_out_0_1_6,
  output     [0:0]    port_state_out_0_1_7,
  output     [0:0]    port_state_out_1_0_0,
  output     [0:0]    port_state_out_1_0_1,
  output     [0:0]    port_state_out_1_0_2,
  output     [0:0]    port_state_out_1_0_3,
  output     [0:0]    port_state_out_1_0_4,
  output     [0:0]    port_state_out_1_0_5,
  output     [0:0]    port_state_out_1_0_6,
  output     [0:0]    port_state_out_1_0_7,
  output     [0:0]    port_state_out_1_1_0,
  output     [0:0]    port_state_out_1_1_1,
  output     [0:0]    port_state_out_1_1_2,
  output     [0:0]    port_state_out_1_1_3,
  output     [0:0]    port_state_out_1_1_4,
  output     [0:0]    port_state_out_1_1_5,
  output     [0:0]    port_state_out_1_1_6,
  output     [0:0]    port_state_out_1_1_7,
  output     [0:0]    port_state_out_2_0_0,
  output     [0:0]    port_state_out_2_0_1,
  output     [0:0]    port_state_out_2_0_2,
  output     [0:0]    port_state_out_2_0_3,
  output     [0:0]    port_state_out_2_0_4,
  output     [0:0]    port_state_out_2_0_5,
  output     [0:0]    port_state_out_2_0_6,
  output     [0:0]    port_state_out_2_0_7,
  output     [0:0]    port_state_out_2_1_0,
  output     [0:0]    port_state_out_2_1_1,
  output     [0:0]    port_state_out_2_1_2,
  output     [0:0]    port_state_out_2_1_3,
  output     [0:0]    port_state_out_2_1_4,
  output     [0:0]    port_state_out_2_1_5,
  output     [0:0]    port_state_out_2_1_6,
  output     [0:0]    port_state_out_2_1_7,
  output     [0:0]    port_state_out_3_0_0,
  output     [0:0]    port_state_out_3_0_1,
  output     [0:0]    port_state_out_3_0_2,
  output     [0:0]    port_state_out_3_0_3,
  output     [0:0]    port_state_out_3_0_4,
  output     [0:0]    port_state_out_3_0_5,
  output     [0:0]    port_state_out_3_0_6,
  output     [0:0]    port_state_out_3_0_7,
  output     [0:0]    port_state_out_3_1_0,
  output     [0:0]    port_state_out_3_1_1,
  output     [0:0]    port_state_out_3_1_2,
  output     [0:0]    port_state_out_3_1_3,
  output     [0:0]    port_state_out_3_1_4,
  output     [0:0]    port_state_out_3_1_5,
  output     [0:0]    port_state_out_3_1_6,
  output     [0:0]    port_state_out_3_1_7,
  output     [0:0]    port_state_out_4_0_0,
  output     [0:0]    port_state_out_4_0_1,
  output     [0:0]    port_state_out_4_0_2,
  output     [0:0]    port_state_out_4_0_3,
  output     [0:0]    port_state_out_4_0_4,
  output     [0:0]    port_state_out_4_0_5,
  output     [0:0]    port_state_out_4_0_6,
  output     [0:0]    port_state_out_4_0_7,
  output     [0:0]    port_state_out_4_1_0,
  output     [0:0]    port_state_out_4_1_1,
  output     [0:0]    port_state_out_4_1_2,
  output     [0:0]    port_state_out_4_1_3,
  output     [0:0]    port_state_out_4_1_4,
  output     [0:0]    port_state_out_4_1_5,
  output     [0:0]    port_state_out_4_1_6,
  output     [0:0]    port_state_out_4_1_7,
  output     [0:0]    port_state_out_5_0_0,
  output     [0:0]    port_state_out_5_0_1,
  output     [0:0]    port_state_out_5_0_2,
  output     [0:0]    port_state_out_5_0_3,
  output     [0:0]    port_state_out_5_0_4,
  output     [0:0]    port_state_out_5_0_5,
  output     [0:0]    port_state_out_5_0_6,
  output     [0:0]    port_state_out_5_0_7,
  output     [0:0]    port_state_out_5_1_0,
  output     [0:0]    port_state_out_5_1_1,
  output     [0:0]    port_state_out_5_1_2,
  output     [0:0]    port_state_out_5_1_3,
  output     [0:0]    port_state_out_5_1_4,
  output     [0:0]    port_state_out_5_1_5,
  output     [0:0]    port_state_out_5_1_6,
  output     [0:0]    port_state_out_5_1_7,
  output     [0:0]    port_state_out_6_0_0,
  output     [0:0]    port_state_out_6_0_1,
  output     [0:0]    port_state_out_6_0_2,
  output     [0:0]    port_state_out_6_0_3,
  output     [0:0]    port_state_out_6_0_4,
  output     [0:0]    port_state_out_6_0_5,
  output     [0:0]    port_state_out_6_0_6,
  output     [0:0]    port_state_out_6_0_7,
  output     [0:0]    port_state_out_6_1_0,
  output     [0:0]    port_state_out_6_1_1,
  output     [0:0]    port_state_out_6_1_2,
  output     [0:0]    port_state_out_6_1_3,
  output     [0:0]    port_state_out_6_1_4,
  output     [0:0]    port_state_out_6_1_5,
  output     [0:0]    port_state_out_6_1_6,
  output     [0:0]    port_state_out_6_1_7,
  output     [0:0]    port_state_out_7_0_0,
  output     [0:0]    port_state_out_7_0_1,
  output     [0:0]    port_state_out_7_0_2,
  output     [0:0]    port_state_out_7_0_3,
  output     [0:0]    port_state_out_7_0_4,
  output     [0:0]    port_state_out_7_0_5,
  output     [0:0]    port_state_out_7_0_6,
  output     [0:0]    port_state_out_7_0_7,
  output     [0:0]    port_state_out_7_1_0,
  output     [0:0]    port_state_out_7_1_1,
  output     [0:0]    port_state_out_7_1_2,
  output     [0:0]    port_state_out_7_1_3,
  output     [0:0]    port_state_out_7_1_4,
  output     [0:0]    port_state_out_7_1_5,
  output     [0:0]    port_state_out_7_1_6,
  output     [0:0]    port_state_out_7_1_7,
  output     [0:0]    port_state_out_8_0_0,
  output     [0:0]    port_state_out_8_0_1,
  output     [0:0]    port_state_out_8_0_2,
  output     [0:0]    port_state_out_8_0_3,
  output     [0:0]    port_state_out_8_0_4,
  output     [0:0]    port_state_out_8_0_5,
  output     [0:0]    port_state_out_8_0_6,
  output     [0:0]    port_state_out_8_0_7,
  output     [0:0]    port_state_out_8_1_0,
  output     [0:0]    port_state_out_8_1_1,
  output     [0:0]    port_state_out_8_1_2,
  output     [0:0]    port_state_out_8_1_3,
  output     [0:0]    port_state_out_8_1_4,
  output     [0:0]    port_state_out_8_1_5,
  output     [0:0]    port_state_out_8_1_6,
  output     [0:0]    port_state_out_8_1_7,
  output     [0:0]    port_state_out_9_0_0,
  output     [0:0]    port_state_out_9_0_1,
  output     [0:0]    port_state_out_9_0_2,
  output     [0:0]    port_state_out_9_0_3,
  output     [0:0]    port_state_out_9_0_4,
  output     [0:0]    port_state_out_9_0_5,
  output     [0:0]    port_state_out_9_0_6,
  output     [0:0]    port_state_out_9_0_7,
  output     [0:0]    port_state_out_9_1_0,
  output     [0:0]    port_state_out_9_1_1,
  output     [0:0]    port_state_out_9_1_2,
  output     [0:0]    port_state_out_9_1_3,
  output     [0:0]    port_state_out_9_1_4,
  output     [0:0]    port_state_out_9_1_5,
  output     [0:0]    port_state_out_9_1_6,
  output     [0:0]    port_state_out_9_1_7,
  output     [0:0]    port_state_out_10_0_0,
  output     [0:0]    port_state_out_10_0_1,
  output     [0:0]    port_state_out_10_0_2,
  output     [0:0]    port_state_out_10_0_3,
  output     [0:0]    port_state_out_10_0_4,
  output     [0:0]    port_state_out_10_0_5,
  output     [0:0]    port_state_out_10_0_6,
  output     [0:0]    port_state_out_10_0_7,
  output     [0:0]    port_state_out_10_1_0,
  output     [0:0]    port_state_out_10_1_1,
  output     [0:0]    port_state_out_10_1_2,
  output     [0:0]    port_state_out_10_1_3,
  output     [0:0]    port_state_out_10_1_4,
  output     [0:0]    port_state_out_10_1_5,
  output     [0:0]    port_state_out_10_1_6,
  output     [0:0]    port_state_out_10_1_7,
  output     [0:0]    port_state_out_11_0_0,
  output     [0:0]    port_state_out_11_0_1,
  output     [0:0]    port_state_out_11_0_2,
  output     [0:0]    port_state_out_11_0_3,
  output     [0:0]    port_state_out_11_0_4,
  output     [0:0]    port_state_out_11_0_5,
  output     [0:0]    port_state_out_11_0_6,
  output     [0:0]    port_state_out_11_0_7,
  output     [0:0]    port_state_out_11_1_0,
  output     [0:0]    port_state_out_11_1_1,
  output     [0:0]    port_state_out_11_1_2,
  output     [0:0]    port_state_out_11_1_3,
  output     [0:0]    port_state_out_11_1_4,
  output     [0:0]    port_state_out_11_1_5,
  output     [0:0]    port_state_out_11_1_6,
  output     [0:0]    port_state_out_11_1_7,
  output     [0:0]    port_state_out_12_0_0,
  output     [0:0]    port_state_out_12_0_1,
  output     [0:0]    port_state_out_12_0_2,
  output     [0:0]    port_state_out_12_0_3,
  output     [0:0]    port_state_out_12_0_4,
  output     [0:0]    port_state_out_12_0_5,
  output     [0:0]    port_state_out_12_0_6,
  output     [0:0]    port_state_out_12_0_7,
  output     [0:0]    port_state_out_12_1_0,
  output     [0:0]    port_state_out_12_1_1,
  output     [0:0]    port_state_out_12_1_2,
  output     [0:0]    port_state_out_12_1_3,
  output     [0:0]    port_state_out_12_1_4,
  output     [0:0]    port_state_out_12_1_5,
  output     [0:0]    port_state_out_12_1_6,
  output     [0:0]    port_state_out_12_1_7,
  output     [0:0]    port_state_out_13_0_0,
  output     [0:0]    port_state_out_13_0_1,
  output     [0:0]    port_state_out_13_0_2,
  output     [0:0]    port_state_out_13_0_3,
  output     [0:0]    port_state_out_13_0_4,
  output     [0:0]    port_state_out_13_0_5,
  output     [0:0]    port_state_out_13_0_6,
  output     [0:0]    port_state_out_13_0_7,
  output     [0:0]    port_state_out_13_1_0,
  output     [0:0]    port_state_out_13_1_1,
  output     [0:0]    port_state_out_13_1_2,
  output     [0:0]    port_state_out_13_1_3,
  output     [0:0]    port_state_out_13_1_4,
  output     [0:0]    port_state_out_13_1_5,
  output     [0:0]    port_state_out_13_1_6,
  output     [0:0]    port_state_out_13_1_7,
  output     [0:0]    port_state_out_14_0_0,
  output     [0:0]    port_state_out_14_0_1,
  output     [0:0]    port_state_out_14_0_2,
  output     [0:0]    port_state_out_14_0_3,
  output     [0:0]    port_state_out_14_0_4,
  output     [0:0]    port_state_out_14_0_5,
  output     [0:0]    port_state_out_14_0_6,
  output     [0:0]    port_state_out_14_0_7,
  output     [0:0]    port_state_out_14_1_0,
  output     [0:0]    port_state_out_14_1_1,
  output     [0:0]    port_state_out_14_1_2,
  output     [0:0]    port_state_out_14_1_3,
  output     [0:0]    port_state_out_14_1_4,
  output     [0:0]    port_state_out_14_1_5,
  output     [0:0]    port_state_out_14_1_6,
  output     [0:0]    port_state_out_14_1_7,
  output     [0:0]    port_state_out_15_0_0,
  output     [0:0]    port_state_out_15_0_1,
  output     [0:0]    port_state_out_15_0_2,
  output     [0:0]    port_state_out_15_0_3,
  output     [0:0]    port_state_out_15_0_4,
  output     [0:0]    port_state_out_15_0_5,
  output     [0:0]    port_state_out_15_0_6,
  output     [0:0]    port_state_out_15_0_7,
  output     [0:0]    port_state_out_15_1_0,
  output     [0:0]    port_state_out_15_1_1,
  output     [0:0]    port_state_out_15_1_2,
  output     [0:0]    port_state_out_15_1_3,
  output     [0:0]    port_state_out_15_1_4,
  output     [0:0]    port_state_out_15_1_5,
  output     [0:0]    port_state_out_15_1_6,
  output     [0:0]    port_state_out_15_1_7,
  input               clk,
  input               reset
);

  wire       [0:0]    keyAdd_port_state_out_0_0_0;
  wire       [0:0]    keyAdd_port_state_out_0_0_1;
  wire       [0:0]    keyAdd_port_state_out_0_0_2;
  wire       [0:0]    keyAdd_port_state_out_0_0_3;
  wire       [0:0]    keyAdd_port_state_out_0_0_4;
  wire       [0:0]    keyAdd_port_state_out_0_0_5;
  wire       [0:0]    keyAdd_port_state_out_0_0_6;
  wire       [0:0]    keyAdd_port_state_out_0_0_7;
  wire       [0:0]    keyAdd_port_state_out_0_1_0;
  wire       [0:0]    keyAdd_port_state_out_0_1_1;
  wire       [0:0]    keyAdd_port_state_out_0_1_2;
  wire       [0:0]    keyAdd_port_state_out_0_1_3;
  wire       [0:0]    keyAdd_port_state_out_0_1_4;
  wire       [0:0]    keyAdd_port_state_out_0_1_5;
  wire       [0:0]    keyAdd_port_state_out_0_1_6;
  wire       [0:0]    keyAdd_port_state_out_0_1_7;
  wire       [0:0]    keyAdd_port_state_out_1_0_0;
  wire       [0:0]    keyAdd_port_state_out_1_0_1;
  wire       [0:0]    keyAdd_port_state_out_1_0_2;
  wire       [0:0]    keyAdd_port_state_out_1_0_3;
  wire       [0:0]    keyAdd_port_state_out_1_0_4;
  wire       [0:0]    keyAdd_port_state_out_1_0_5;
  wire       [0:0]    keyAdd_port_state_out_1_0_6;
  wire       [0:0]    keyAdd_port_state_out_1_0_7;
  wire       [0:0]    keyAdd_port_state_out_1_1_0;
  wire       [0:0]    keyAdd_port_state_out_1_1_1;
  wire       [0:0]    keyAdd_port_state_out_1_1_2;
  wire       [0:0]    keyAdd_port_state_out_1_1_3;
  wire       [0:0]    keyAdd_port_state_out_1_1_4;
  wire       [0:0]    keyAdd_port_state_out_1_1_5;
  wire       [0:0]    keyAdd_port_state_out_1_1_6;
  wire       [0:0]    keyAdd_port_state_out_1_1_7;
  wire       [0:0]    keyAdd_port_state_out_2_0_0;
  wire       [0:0]    keyAdd_port_state_out_2_0_1;
  wire       [0:0]    keyAdd_port_state_out_2_0_2;
  wire       [0:0]    keyAdd_port_state_out_2_0_3;
  wire       [0:0]    keyAdd_port_state_out_2_0_4;
  wire       [0:0]    keyAdd_port_state_out_2_0_5;
  wire       [0:0]    keyAdd_port_state_out_2_0_6;
  wire       [0:0]    keyAdd_port_state_out_2_0_7;
  wire       [0:0]    keyAdd_port_state_out_2_1_0;
  wire       [0:0]    keyAdd_port_state_out_2_1_1;
  wire       [0:0]    keyAdd_port_state_out_2_1_2;
  wire       [0:0]    keyAdd_port_state_out_2_1_3;
  wire       [0:0]    keyAdd_port_state_out_2_1_4;
  wire       [0:0]    keyAdd_port_state_out_2_1_5;
  wire       [0:0]    keyAdd_port_state_out_2_1_6;
  wire       [0:0]    keyAdd_port_state_out_2_1_7;
  wire       [0:0]    keyAdd_port_state_out_3_0_0;
  wire       [0:0]    keyAdd_port_state_out_3_0_1;
  wire       [0:0]    keyAdd_port_state_out_3_0_2;
  wire       [0:0]    keyAdd_port_state_out_3_0_3;
  wire       [0:0]    keyAdd_port_state_out_3_0_4;
  wire       [0:0]    keyAdd_port_state_out_3_0_5;
  wire       [0:0]    keyAdd_port_state_out_3_0_6;
  wire       [0:0]    keyAdd_port_state_out_3_0_7;
  wire       [0:0]    keyAdd_port_state_out_3_1_0;
  wire       [0:0]    keyAdd_port_state_out_3_1_1;
  wire       [0:0]    keyAdd_port_state_out_3_1_2;
  wire       [0:0]    keyAdd_port_state_out_3_1_3;
  wire       [0:0]    keyAdd_port_state_out_3_1_4;
  wire       [0:0]    keyAdd_port_state_out_3_1_5;
  wire       [0:0]    keyAdd_port_state_out_3_1_6;
  wire       [0:0]    keyAdd_port_state_out_3_1_7;
  wire       [0:0]    keyAdd_port_state_out_4_0_0;
  wire       [0:0]    keyAdd_port_state_out_4_0_1;
  wire       [0:0]    keyAdd_port_state_out_4_0_2;
  wire       [0:0]    keyAdd_port_state_out_4_0_3;
  wire       [0:0]    keyAdd_port_state_out_4_0_4;
  wire       [0:0]    keyAdd_port_state_out_4_0_5;
  wire       [0:0]    keyAdd_port_state_out_4_0_6;
  wire       [0:0]    keyAdd_port_state_out_4_0_7;
  wire       [0:0]    keyAdd_port_state_out_4_1_0;
  wire       [0:0]    keyAdd_port_state_out_4_1_1;
  wire       [0:0]    keyAdd_port_state_out_4_1_2;
  wire       [0:0]    keyAdd_port_state_out_4_1_3;
  wire       [0:0]    keyAdd_port_state_out_4_1_4;
  wire       [0:0]    keyAdd_port_state_out_4_1_5;
  wire       [0:0]    keyAdd_port_state_out_4_1_6;
  wire       [0:0]    keyAdd_port_state_out_4_1_7;
  wire       [0:0]    keyAdd_port_state_out_5_0_0;
  wire       [0:0]    keyAdd_port_state_out_5_0_1;
  wire       [0:0]    keyAdd_port_state_out_5_0_2;
  wire       [0:0]    keyAdd_port_state_out_5_0_3;
  wire       [0:0]    keyAdd_port_state_out_5_0_4;
  wire       [0:0]    keyAdd_port_state_out_5_0_5;
  wire       [0:0]    keyAdd_port_state_out_5_0_6;
  wire       [0:0]    keyAdd_port_state_out_5_0_7;
  wire       [0:0]    keyAdd_port_state_out_5_1_0;
  wire       [0:0]    keyAdd_port_state_out_5_1_1;
  wire       [0:0]    keyAdd_port_state_out_5_1_2;
  wire       [0:0]    keyAdd_port_state_out_5_1_3;
  wire       [0:0]    keyAdd_port_state_out_5_1_4;
  wire       [0:0]    keyAdd_port_state_out_5_1_5;
  wire       [0:0]    keyAdd_port_state_out_5_1_6;
  wire       [0:0]    keyAdd_port_state_out_5_1_7;
  wire       [0:0]    keyAdd_port_state_out_6_0_0;
  wire       [0:0]    keyAdd_port_state_out_6_0_1;
  wire       [0:0]    keyAdd_port_state_out_6_0_2;
  wire       [0:0]    keyAdd_port_state_out_6_0_3;
  wire       [0:0]    keyAdd_port_state_out_6_0_4;
  wire       [0:0]    keyAdd_port_state_out_6_0_5;
  wire       [0:0]    keyAdd_port_state_out_6_0_6;
  wire       [0:0]    keyAdd_port_state_out_6_0_7;
  wire       [0:0]    keyAdd_port_state_out_6_1_0;
  wire       [0:0]    keyAdd_port_state_out_6_1_1;
  wire       [0:0]    keyAdd_port_state_out_6_1_2;
  wire       [0:0]    keyAdd_port_state_out_6_1_3;
  wire       [0:0]    keyAdd_port_state_out_6_1_4;
  wire       [0:0]    keyAdd_port_state_out_6_1_5;
  wire       [0:0]    keyAdd_port_state_out_6_1_6;
  wire       [0:0]    keyAdd_port_state_out_6_1_7;
  wire       [0:0]    keyAdd_port_state_out_7_0_0;
  wire       [0:0]    keyAdd_port_state_out_7_0_1;
  wire       [0:0]    keyAdd_port_state_out_7_0_2;
  wire       [0:0]    keyAdd_port_state_out_7_0_3;
  wire       [0:0]    keyAdd_port_state_out_7_0_4;
  wire       [0:0]    keyAdd_port_state_out_7_0_5;
  wire       [0:0]    keyAdd_port_state_out_7_0_6;
  wire       [0:0]    keyAdd_port_state_out_7_0_7;
  wire       [0:0]    keyAdd_port_state_out_7_1_0;
  wire       [0:0]    keyAdd_port_state_out_7_1_1;
  wire       [0:0]    keyAdd_port_state_out_7_1_2;
  wire       [0:0]    keyAdd_port_state_out_7_1_3;
  wire       [0:0]    keyAdd_port_state_out_7_1_4;
  wire       [0:0]    keyAdd_port_state_out_7_1_5;
  wire       [0:0]    keyAdd_port_state_out_7_1_6;
  wire       [0:0]    keyAdd_port_state_out_7_1_7;
  wire       [0:0]    keyAdd_port_state_out_8_0_0;
  wire       [0:0]    keyAdd_port_state_out_8_0_1;
  wire       [0:0]    keyAdd_port_state_out_8_0_2;
  wire       [0:0]    keyAdd_port_state_out_8_0_3;
  wire       [0:0]    keyAdd_port_state_out_8_0_4;
  wire       [0:0]    keyAdd_port_state_out_8_0_5;
  wire       [0:0]    keyAdd_port_state_out_8_0_6;
  wire       [0:0]    keyAdd_port_state_out_8_0_7;
  wire       [0:0]    keyAdd_port_state_out_8_1_0;
  wire       [0:0]    keyAdd_port_state_out_8_1_1;
  wire       [0:0]    keyAdd_port_state_out_8_1_2;
  wire       [0:0]    keyAdd_port_state_out_8_1_3;
  wire       [0:0]    keyAdd_port_state_out_8_1_4;
  wire       [0:0]    keyAdd_port_state_out_8_1_5;
  wire       [0:0]    keyAdd_port_state_out_8_1_6;
  wire       [0:0]    keyAdd_port_state_out_8_1_7;
  wire       [0:0]    keyAdd_port_state_out_9_0_0;
  wire       [0:0]    keyAdd_port_state_out_9_0_1;
  wire       [0:0]    keyAdd_port_state_out_9_0_2;
  wire       [0:0]    keyAdd_port_state_out_9_0_3;
  wire       [0:0]    keyAdd_port_state_out_9_0_4;
  wire       [0:0]    keyAdd_port_state_out_9_0_5;
  wire       [0:0]    keyAdd_port_state_out_9_0_6;
  wire       [0:0]    keyAdd_port_state_out_9_0_7;
  wire       [0:0]    keyAdd_port_state_out_9_1_0;
  wire       [0:0]    keyAdd_port_state_out_9_1_1;
  wire       [0:0]    keyAdd_port_state_out_9_1_2;
  wire       [0:0]    keyAdd_port_state_out_9_1_3;
  wire       [0:0]    keyAdd_port_state_out_9_1_4;
  wire       [0:0]    keyAdd_port_state_out_9_1_5;
  wire       [0:0]    keyAdd_port_state_out_9_1_6;
  wire       [0:0]    keyAdd_port_state_out_9_1_7;
  wire       [0:0]    keyAdd_port_state_out_10_0_0;
  wire       [0:0]    keyAdd_port_state_out_10_0_1;
  wire       [0:0]    keyAdd_port_state_out_10_0_2;
  wire       [0:0]    keyAdd_port_state_out_10_0_3;
  wire       [0:0]    keyAdd_port_state_out_10_0_4;
  wire       [0:0]    keyAdd_port_state_out_10_0_5;
  wire       [0:0]    keyAdd_port_state_out_10_0_6;
  wire       [0:0]    keyAdd_port_state_out_10_0_7;
  wire       [0:0]    keyAdd_port_state_out_10_1_0;
  wire       [0:0]    keyAdd_port_state_out_10_1_1;
  wire       [0:0]    keyAdd_port_state_out_10_1_2;
  wire       [0:0]    keyAdd_port_state_out_10_1_3;
  wire       [0:0]    keyAdd_port_state_out_10_1_4;
  wire       [0:0]    keyAdd_port_state_out_10_1_5;
  wire       [0:0]    keyAdd_port_state_out_10_1_6;
  wire       [0:0]    keyAdd_port_state_out_10_1_7;
  wire       [0:0]    keyAdd_port_state_out_11_0_0;
  wire       [0:0]    keyAdd_port_state_out_11_0_1;
  wire       [0:0]    keyAdd_port_state_out_11_0_2;
  wire       [0:0]    keyAdd_port_state_out_11_0_3;
  wire       [0:0]    keyAdd_port_state_out_11_0_4;
  wire       [0:0]    keyAdd_port_state_out_11_0_5;
  wire       [0:0]    keyAdd_port_state_out_11_0_6;
  wire       [0:0]    keyAdd_port_state_out_11_0_7;
  wire       [0:0]    keyAdd_port_state_out_11_1_0;
  wire       [0:0]    keyAdd_port_state_out_11_1_1;
  wire       [0:0]    keyAdd_port_state_out_11_1_2;
  wire       [0:0]    keyAdd_port_state_out_11_1_3;
  wire       [0:0]    keyAdd_port_state_out_11_1_4;
  wire       [0:0]    keyAdd_port_state_out_11_1_5;
  wire       [0:0]    keyAdd_port_state_out_11_1_6;
  wire       [0:0]    keyAdd_port_state_out_11_1_7;
  wire       [0:0]    keyAdd_port_state_out_12_0_0;
  wire       [0:0]    keyAdd_port_state_out_12_0_1;
  wire       [0:0]    keyAdd_port_state_out_12_0_2;
  wire       [0:0]    keyAdd_port_state_out_12_0_3;
  wire       [0:0]    keyAdd_port_state_out_12_0_4;
  wire       [0:0]    keyAdd_port_state_out_12_0_5;
  wire       [0:0]    keyAdd_port_state_out_12_0_6;
  wire       [0:0]    keyAdd_port_state_out_12_0_7;
  wire       [0:0]    keyAdd_port_state_out_12_1_0;
  wire       [0:0]    keyAdd_port_state_out_12_1_1;
  wire       [0:0]    keyAdd_port_state_out_12_1_2;
  wire       [0:0]    keyAdd_port_state_out_12_1_3;
  wire       [0:0]    keyAdd_port_state_out_12_1_4;
  wire       [0:0]    keyAdd_port_state_out_12_1_5;
  wire       [0:0]    keyAdd_port_state_out_12_1_6;
  wire       [0:0]    keyAdd_port_state_out_12_1_7;
  wire       [0:0]    keyAdd_port_state_out_13_0_0;
  wire       [0:0]    keyAdd_port_state_out_13_0_1;
  wire       [0:0]    keyAdd_port_state_out_13_0_2;
  wire       [0:0]    keyAdd_port_state_out_13_0_3;
  wire       [0:0]    keyAdd_port_state_out_13_0_4;
  wire       [0:0]    keyAdd_port_state_out_13_0_5;
  wire       [0:0]    keyAdd_port_state_out_13_0_6;
  wire       [0:0]    keyAdd_port_state_out_13_0_7;
  wire       [0:0]    keyAdd_port_state_out_13_1_0;
  wire       [0:0]    keyAdd_port_state_out_13_1_1;
  wire       [0:0]    keyAdd_port_state_out_13_1_2;
  wire       [0:0]    keyAdd_port_state_out_13_1_3;
  wire       [0:0]    keyAdd_port_state_out_13_1_4;
  wire       [0:0]    keyAdd_port_state_out_13_1_5;
  wire       [0:0]    keyAdd_port_state_out_13_1_6;
  wire       [0:0]    keyAdd_port_state_out_13_1_7;
  wire       [0:0]    keyAdd_port_state_out_14_0_0;
  wire       [0:0]    keyAdd_port_state_out_14_0_1;
  wire       [0:0]    keyAdd_port_state_out_14_0_2;
  wire       [0:0]    keyAdd_port_state_out_14_0_3;
  wire       [0:0]    keyAdd_port_state_out_14_0_4;
  wire       [0:0]    keyAdd_port_state_out_14_0_5;
  wire       [0:0]    keyAdd_port_state_out_14_0_6;
  wire       [0:0]    keyAdd_port_state_out_14_0_7;
  wire       [0:0]    keyAdd_port_state_out_14_1_0;
  wire       [0:0]    keyAdd_port_state_out_14_1_1;
  wire       [0:0]    keyAdd_port_state_out_14_1_2;
  wire       [0:0]    keyAdd_port_state_out_14_1_3;
  wire       [0:0]    keyAdd_port_state_out_14_1_4;
  wire       [0:0]    keyAdd_port_state_out_14_1_5;
  wire       [0:0]    keyAdd_port_state_out_14_1_6;
  wire       [0:0]    keyAdd_port_state_out_14_1_7;
  wire       [0:0]    keyAdd_port_state_out_15_0_0;
  wire       [0:0]    keyAdd_port_state_out_15_0_1;
  wire       [0:0]    keyAdd_port_state_out_15_0_2;
  wire       [0:0]    keyAdd_port_state_out_15_0_3;
  wire       [0:0]    keyAdd_port_state_out_15_0_4;
  wire       [0:0]    keyAdd_port_state_out_15_0_5;
  wire       [0:0]    keyAdd_port_state_out_15_0_6;
  wire       [0:0]    keyAdd_port_state_out_15_0_7;
  wire       [0:0]    keyAdd_port_state_out_15_1_0;
  wire       [0:0]    keyAdd_port_state_out_15_1_1;
  wire       [0:0]    keyAdd_port_state_out_15_1_2;
  wire       [0:0]    keyAdd_port_state_out_15_1_3;
  wire       [0:0]    keyAdd_port_state_out_15_1_4;
  wire       [0:0]    keyAdd_port_state_out_15_1_5;
  wire       [0:0]    keyAdd_port_state_out_15_1_6;
  wire       [0:0]    keyAdd_port_state_out_15_1_7;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_16_port_o_0_0;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_16_port_o_0_1;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_16_port_o_0_2;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_16_port_o_0_3;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_16_port_o_0_4;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_16_port_o_0_5;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_16_port_o_0_6;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_16_port_o_0_7;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_16_port_o_1_0;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_16_port_o_1_1;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_16_port_o_1_2;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_16_port_o_1_3;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_16_port_o_1_4;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_16_port_o_1_5;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_16_port_o_1_6;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_16_port_o_1_7;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_17_port_o_0_0;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_17_port_o_0_1;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_17_port_o_0_2;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_17_port_o_0_3;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_17_port_o_0_4;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_17_port_o_0_5;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_17_port_o_0_6;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_17_port_o_0_7;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_17_port_o_1_0;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_17_port_o_1_1;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_17_port_o_1_2;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_17_port_o_1_3;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_17_port_o_1_4;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_17_port_o_1_5;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_17_port_o_1_6;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_17_port_o_1_7;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_18_port_o_0_0;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_18_port_o_0_1;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_18_port_o_0_2;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_18_port_o_0_3;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_18_port_o_0_4;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_18_port_o_0_5;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_18_port_o_0_6;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_18_port_o_0_7;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_18_port_o_1_0;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_18_port_o_1_1;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_18_port_o_1_2;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_18_port_o_1_3;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_18_port_o_1_4;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_18_port_o_1_5;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_18_port_o_1_6;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_18_port_o_1_7;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_19_port_o_0_0;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_19_port_o_0_1;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_19_port_o_0_2;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_19_port_o_0_3;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_19_port_o_0_4;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_19_port_o_0_5;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_19_port_o_0_6;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_19_port_o_0_7;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_19_port_o_1_0;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_19_port_o_1_1;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_19_port_o_1_2;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_19_port_o_1_3;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_19_port_o_1_4;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_19_port_o_1_5;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_19_port_o_1_6;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_19_port_o_1_7;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_20_port_o_0_0;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_20_port_o_0_1;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_20_port_o_0_2;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_20_port_o_0_3;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_20_port_o_0_4;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_20_port_o_0_5;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_20_port_o_0_6;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_20_port_o_0_7;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_20_port_o_1_0;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_20_port_o_1_1;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_20_port_o_1_2;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_20_port_o_1_3;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_20_port_o_1_4;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_20_port_o_1_5;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_20_port_o_1_6;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_20_port_o_1_7;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_21_port_o_0_0;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_21_port_o_0_1;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_21_port_o_0_2;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_21_port_o_0_3;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_21_port_o_0_4;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_21_port_o_0_5;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_21_port_o_0_6;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_21_port_o_0_7;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_21_port_o_1_0;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_21_port_o_1_1;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_21_port_o_1_2;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_21_port_o_1_3;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_21_port_o_1_4;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_21_port_o_1_5;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_21_port_o_1_6;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_21_port_o_1_7;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_22_port_o_0_0;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_22_port_o_0_1;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_22_port_o_0_2;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_22_port_o_0_3;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_22_port_o_0_4;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_22_port_o_0_5;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_22_port_o_0_6;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_22_port_o_0_7;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_22_port_o_1_0;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_22_port_o_1_1;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_22_port_o_1_2;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_22_port_o_1_3;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_22_port_o_1_4;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_22_port_o_1_5;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_22_port_o_1_6;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_22_port_o_1_7;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_23_port_o_0_0;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_23_port_o_0_1;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_23_port_o_0_2;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_23_port_o_0_3;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_23_port_o_0_4;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_23_port_o_0_5;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_23_port_o_0_6;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_23_port_o_0_7;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_23_port_o_1_0;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_23_port_o_1_1;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_23_port_o_1_2;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_23_port_o_1_3;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_23_port_o_1_4;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_23_port_o_1_5;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_23_port_o_1_6;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_23_port_o_1_7;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_24_port_o_0_0;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_24_port_o_0_1;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_24_port_o_0_2;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_24_port_o_0_3;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_24_port_o_0_4;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_24_port_o_0_5;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_24_port_o_0_6;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_24_port_o_0_7;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_24_port_o_1_0;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_24_port_o_1_1;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_24_port_o_1_2;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_24_port_o_1_3;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_24_port_o_1_4;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_24_port_o_1_5;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_24_port_o_1_6;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_24_port_o_1_7;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_25_port_o_0_0;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_25_port_o_0_1;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_25_port_o_0_2;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_25_port_o_0_3;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_25_port_o_0_4;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_25_port_o_0_5;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_25_port_o_0_6;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_25_port_o_0_7;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_25_port_o_1_0;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_25_port_o_1_1;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_25_port_o_1_2;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_25_port_o_1_3;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_25_port_o_1_4;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_25_port_o_1_5;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_25_port_o_1_6;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_25_port_o_1_7;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_26_port_o_0_0;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_26_port_o_0_1;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_26_port_o_0_2;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_26_port_o_0_3;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_26_port_o_0_4;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_26_port_o_0_5;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_26_port_o_0_6;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_26_port_o_0_7;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_26_port_o_1_0;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_26_port_o_1_1;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_26_port_o_1_2;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_26_port_o_1_3;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_26_port_o_1_4;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_26_port_o_1_5;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_26_port_o_1_6;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_26_port_o_1_7;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_27_port_o_0_0;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_27_port_o_0_1;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_27_port_o_0_2;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_27_port_o_0_3;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_27_port_o_0_4;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_27_port_o_0_5;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_27_port_o_0_6;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_27_port_o_0_7;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_27_port_o_1_0;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_27_port_o_1_1;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_27_port_o_1_2;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_27_port_o_1_3;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_27_port_o_1_4;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_27_port_o_1_5;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_27_port_o_1_6;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_27_port_o_1_7;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_28_port_o_0_0;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_28_port_o_0_1;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_28_port_o_0_2;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_28_port_o_0_3;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_28_port_o_0_4;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_28_port_o_0_5;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_28_port_o_0_6;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_28_port_o_0_7;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_28_port_o_1_0;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_28_port_o_1_1;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_28_port_o_1_2;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_28_port_o_1_3;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_28_port_o_1_4;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_28_port_o_1_5;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_28_port_o_1_6;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_28_port_o_1_7;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_29_port_o_0_0;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_29_port_o_0_1;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_29_port_o_0_2;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_29_port_o_0_3;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_29_port_o_0_4;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_29_port_o_0_5;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_29_port_o_0_6;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_29_port_o_0_7;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_29_port_o_1_0;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_29_port_o_1_1;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_29_port_o_1_2;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_29_port_o_1_3;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_29_port_o_1_4;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_29_port_o_1_5;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_29_port_o_1_6;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_29_port_o_1_7;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_30_port_o_0_0;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_30_port_o_0_1;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_30_port_o_0_2;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_30_port_o_0_3;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_30_port_o_0_4;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_30_port_o_0_5;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_30_port_o_0_6;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_30_port_o_0_7;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_30_port_o_1_0;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_30_port_o_1_1;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_30_port_o_1_2;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_30_port_o_1_3;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_30_port_o_1_4;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_30_port_o_1_5;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_30_port_o_1_6;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_30_port_o_1_7;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_31_port_o_0_0;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_31_port_o_0_1;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_31_port_o_0_2;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_31_port_o_0_3;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_31_port_o_0_4;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_31_port_o_0_5;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_31_port_o_0_6;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_31_port_o_0_7;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_31_port_o_1_0;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_31_port_o_1_1;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_31_port_o_1_2;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_31_port_o_1_3;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_31_port_o_1_4;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_31_port_o_1_5;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_31_port_o_1_6;
  wire       [0:0]    sbox_AES_Canright_CMS_2shares_31_port_o_1_7;
  wire       [0:0]    shiftRows_port_state_out_0_0_0;
  wire       [0:0]    shiftRows_port_state_out_0_0_1;
  wire       [0:0]    shiftRows_port_state_out_0_0_2;
  wire       [0:0]    shiftRows_port_state_out_0_0_3;
  wire       [0:0]    shiftRows_port_state_out_0_0_4;
  wire       [0:0]    shiftRows_port_state_out_0_0_5;
  wire       [0:0]    shiftRows_port_state_out_0_0_6;
  wire       [0:0]    shiftRows_port_state_out_0_0_7;
  wire       [0:0]    shiftRows_port_state_out_0_1_0;
  wire       [0:0]    shiftRows_port_state_out_0_1_1;
  wire       [0:0]    shiftRows_port_state_out_0_1_2;
  wire       [0:0]    shiftRows_port_state_out_0_1_3;
  wire       [0:0]    shiftRows_port_state_out_0_1_4;
  wire       [0:0]    shiftRows_port_state_out_0_1_5;
  wire       [0:0]    shiftRows_port_state_out_0_1_6;
  wire       [0:0]    shiftRows_port_state_out_0_1_7;
  wire       [0:0]    shiftRows_port_state_out_1_0_0;
  wire       [0:0]    shiftRows_port_state_out_1_0_1;
  wire       [0:0]    shiftRows_port_state_out_1_0_2;
  wire       [0:0]    shiftRows_port_state_out_1_0_3;
  wire       [0:0]    shiftRows_port_state_out_1_0_4;
  wire       [0:0]    shiftRows_port_state_out_1_0_5;
  wire       [0:0]    shiftRows_port_state_out_1_0_6;
  wire       [0:0]    shiftRows_port_state_out_1_0_7;
  wire       [0:0]    shiftRows_port_state_out_1_1_0;
  wire       [0:0]    shiftRows_port_state_out_1_1_1;
  wire       [0:0]    shiftRows_port_state_out_1_1_2;
  wire       [0:0]    shiftRows_port_state_out_1_1_3;
  wire       [0:0]    shiftRows_port_state_out_1_1_4;
  wire       [0:0]    shiftRows_port_state_out_1_1_5;
  wire       [0:0]    shiftRows_port_state_out_1_1_6;
  wire       [0:0]    shiftRows_port_state_out_1_1_7;
  wire       [0:0]    shiftRows_port_state_out_2_0_0;
  wire       [0:0]    shiftRows_port_state_out_2_0_1;
  wire       [0:0]    shiftRows_port_state_out_2_0_2;
  wire       [0:0]    shiftRows_port_state_out_2_0_3;
  wire       [0:0]    shiftRows_port_state_out_2_0_4;
  wire       [0:0]    shiftRows_port_state_out_2_0_5;
  wire       [0:0]    shiftRows_port_state_out_2_0_6;
  wire       [0:0]    shiftRows_port_state_out_2_0_7;
  wire       [0:0]    shiftRows_port_state_out_2_1_0;
  wire       [0:0]    shiftRows_port_state_out_2_1_1;
  wire       [0:0]    shiftRows_port_state_out_2_1_2;
  wire       [0:0]    shiftRows_port_state_out_2_1_3;
  wire       [0:0]    shiftRows_port_state_out_2_1_4;
  wire       [0:0]    shiftRows_port_state_out_2_1_5;
  wire       [0:0]    shiftRows_port_state_out_2_1_6;
  wire       [0:0]    shiftRows_port_state_out_2_1_7;
  wire       [0:0]    shiftRows_port_state_out_3_0_0;
  wire       [0:0]    shiftRows_port_state_out_3_0_1;
  wire       [0:0]    shiftRows_port_state_out_3_0_2;
  wire       [0:0]    shiftRows_port_state_out_3_0_3;
  wire       [0:0]    shiftRows_port_state_out_3_0_4;
  wire       [0:0]    shiftRows_port_state_out_3_0_5;
  wire       [0:0]    shiftRows_port_state_out_3_0_6;
  wire       [0:0]    shiftRows_port_state_out_3_0_7;
  wire       [0:0]    shiftRows_port_state_out_3_1_0;
  wire       [0:0]    shiftRows_port_state_out_3_1_1;
  wire       [0:0]    shiftRows_port_state_out_3_1_2;
  wire       [0:0]    shiftRows_port_state_out_3_1_3;
  wire       [0:0]    shiftRows_port_state_out_3_1_4;
  wire       [0:0]    shiftRows_port_state_out_3_1_5;
  wire       [0:0]    shiftRows_port_state_out_3_1_6;
  wire       [0:0]    shiftRows_port_state_out_3_1_7;
  wire       [0:0]    shiftRows_port_state_out_4_0_0;
  wire       [0:0]    shiftRows_port_state_out_4_0_1;
  wire       [0:0]    shiftRows_port_state_out_4_0_2;
  wire       [0:0]    shiftRows_port_state_out_4_0_3;
  wire       [0:0]    shiftRows_port_state_out_4_0_4;
  wire       [0:0]    shiftRows_port_state_out_4_0_5;
  wire       [0:0]    shiftRows_port_state_out_4_0_6;
  wire       [0:0]    shiftRows_port_state_out_4_0_7;
  wire       [0:0]    shiftRows_port_state_out_4_1_0;
  wire       [0:0]    shiftRows_port_state_out_4_1_1;
  wire       [0:0]    shiftRows_port_state_out_4_1_2;
  wire       [0:0]    shiftRows_port_state_out_4_1_3;
  wire       [0:0]    shiftRows_port_state_out_4_1_4;
  wire       [0:0]    shiftRows_port_state_out_4_1_5;
  wire       [0:0]    shiftRows_port_state_out_4_1_6;
  wire       [0:0]    shiftRows_port_state_out_4_1_7;
  wire       [0:0]    shiftRows_port_state_out_5_0_0;
  wire       [0:0]    shiftRows_port_state_out_5_0_1;
  wire       [0:0]    shiftRows_port_state_out_5_0_2;
  wire       [0:0]    shiftRows_port_state_out_5_0_3;
  wire       [0:0]    shiftRows_port_state_out_5_0_4;
  wire       [0:0]    shiftRows_port_state_out_5_0_5;
  wire       [0:0]    shiftRows_port_state_out_5_0_6;
  wire       [0:0]    shiftRows_port_state_out_5_0_7;
  wire       [0:0]    shiftRows_port_state_out_5_1_0;
  wire       [0:0]    shiftRows_port_state_out_5_1_1;
  wire       [0:0]    shiftRows_port_state_out_5_1_2;
  wire       [0:0]    shiftRows_port_state_out_5_1_3;
  wire       [0:0]    shiftRows_port_state_out_5_1_4;
  wire       [0:0]    shiftRows_port_state_out_5_1_5;
  wire       [0:0]    shiftRows_port_state_out_5_1_6;
  wire       [0:0]    shiftRows_port_state_out_5_1_7;
  wire       [0:0]    shiftRows_port_state_out_6_0_0;
  wire       [0:0]    shiftRows_port_state_out_6_0_1;
  wire       [0:0]    shiftRows_port_state_out_6_0_2;
  wire       [0:0]    shiftRows_port_state_out_6_0_3;
  wire       [0:0]    shiftRows_port_state_out_6_0_4;
  wire       [0:0]    shiftRows_port_state_out_6_0_5;
  wire       [0:0]    shiftRows_port_state_out_6_0_6;
  wire       [0:0]    shiftRows_port_state_out_6_0_7;
  wire       [0:0]    shiftRows_port_state_out_6_1_0;
  wire       [0:0]    shiftRows_port_state_out_6_1_1;
  wire       [0:0]    shiftRows_port_state_out_6_1_2;
  wire       [0:0]    shiftRows_port_state_out_6_1_3;
  wire       [0:0]    shiftRows_port_state_out_6_1_4;
  wire       [0:0]    shiftRows_port_state_out_6_1_5;
  wire       [0:0]    shiftRows_port_state_out_6_1_6;
  wire       [0:0]    shiftRows_port_state_out_6_1_7;
  wire       [0:0]    shiftRows_port_state_out_7_0_0;
  wire       [0:0]    shiftRows_port_state_out_7_0_1;
  wire       [0:0]    shiftRows_port_state_out_7_0_2;
  wire       [0:0]    shiftRows_port_state_out_7_0_3;
  wire       [0:0]    shiftRows_port_state_out_7_0_4;
  wire       [0:0]    shiftRows_port_state_out_7_0_5;
  wire       [0:0]    shiftRows_port_state_out_7_0_6;
  wire       [0:0]    shiftRows_port_state_out_7_0_7;
  wire       [0:0]    shiftRows_port_state_out_7_1_0;
  wire       [0:0]    shiftRows_port_state_out_7_1_1;
  wire       [0:0]    shiftRows_port_state_out_7_1_2;
  wire       [0:0]    shiftRows_port_state_out_7_1_3;
  wire       [0:0]    shiftRows_port_state_out_7_1_4;
  wire       [0:0]    shiftRows_port_state_out_7_1_5;
  wire       [0:0]    shiftRows_port_state_out_7_1_6;
  wire       [0:0]    shiftRows_port_state_out_7_1_7;
  wire       [0:0]    shiftRows_port_state_out_8_0_0;
  wire       [0:0]    shiftRows_port_state_out_8_0_1;
  wire       [0:0]    shiftRows_port_state_out_8_0_2;
  wire       [0:0]    shiftRows_port_state_out_8_0_3;
  wire       [0:0]    shiftRows_port_state_out_8_0_4;
  wire       [0:0]    shiftRows_port_state_out_8_0_5;
  wire       [0:0]    shiftRows_port_state_out_8_0_6;
  wire       [0:0]    shiftRows_port_state_out_8_0_7;
  wire       [0:0]    shiftRows_port_state_out_8_1_0;
  wire       [0:0]    shiftRows_port_state_out_8_1_1;
  wire       [0:0]    shiftRows_port_state_out_8_1_2;
  wire       [0:0]    shiftRows_port_state_out_8_1_3;
  wire       [0:0]    shiftRows_port_state_out_8_1_4;
  wire       [0:0]    shiftRows_port_state_out_8_1_5;
  wire       [0:0]    shiftRows_port_state_out_8_1_6;
  wire       [0:0]    shiftRows_port_state_out_8_1_7;
  wire       [0:0]    shiftRows_port_state_out_9_0_0;
  wire       [0:0]    shiftRows_port_state_out_9_0_1;
  wire       [0:0]    shiftRows_port_state_out_9_0_2;
  wire       [0:0]    shiftRows_port_state_out_9_0_3;
  wire       [0:0]    shiftRows_port_state_out_9_0_4;
  wire       [0:0]    shiftRows_port_state_out_9_0_5;
  wire       [0:0]    shiftRows_port_state_out_9_0_6;
  wire       [0:0]    shiftRows_port_state_out_9_0_7;
  wire       [0:0]    shiftRows_port_state_out_9_1_0;
  wire       [0:0]    shiftRows_port_state_out_9_1_1;
  wire       [0:0]    shiftRows_port_state_out_9_1_2;
  wire       [0:0]    shiftRows_port_state_out_9_1_3;
  wire       [0:0]    shiftRows_port_state_out_9_1_4;
  wire       [0:0]    shiftRows_port_state_out_9_1_5;
  wire       [0:0]    shiftRows_port_state_out_9_1_6;
  wire       [0:0]    shiftRows_port_state_out_9_1_7;
  wire       [0:0]    shiftRows_port_state_out_10_0_0;
  wire       [0:0]    shiftRows_port_state_out_10_0_1;
  wire       [0:0]    shiftRows_port_state_out_10_0_2;
  wire       [0:0]    shiftRows_port_state_out_10_0_3;
  wire       [0:0]    shiftRows_port_state_out_10_0_4;
  wire       [0:0]    shiftRows_port_state_out_10_0_5;
  wire       [0:0]    shiftRows_port_state_out_10_0_6;
  wire       [0:0]    shiftRows_port_state_out_10_0_7;
  wire       [0:0]    shiftRows_port_state_out_10_1_0;
  wire       [0:0]    shiftRows_port_state_out_10_1_1;
  wire       [0:0]    shiftRows_port_state_out_10_1_2;
  wire       [0:0]    shiftRows_port_state_out_10_1_3;
  wire       [0:0]    shiftRows_port_state_out_10_1_4;
  wire       [0:0]    shiftRows_port_state_out_10_1_5;
  wire       [0:0]    shiftRows_port_state_out_10_1_6;
  wire       [0:0]    shiftRows_port_state_out_10_1_7;
  wire       [0:0]    shiftRows_port_state_out_11_0_0;
  wire       [0:0]    shiftRows_port_state_out_11_0_1;
  wire       [0:0]    shiftRows_port_state_out_11_0_2;
  wire       [0:0]    shiftRows_port_state_out_11_0_3;
  wire       [0:0]    shiftRows_port_state_out_11_0_4;
  wire       [0:0]    shiftRows_port_state_out_11_0_5;
  wire       [0:0]    shiftRows_port_state_out_11_0_6;
  wire       [0:0]    shiftRows_port_state_out_11_0_7;
  wire       [0:0]    shiftRows_port_state_out_11_1_0;
  wire       [0:0]    shiftRows_port_state_out_11_1_1;
  wire       [0:0]    shiftRows_port_state_out_11_1_2;
  wire       [0:0]    shiftRows_port_state_out_11_1_3;
  wire       [0:0]    shiftRows_port_state_out_11_1_4;
  wire       [0:0]    shiftRows_port_state_out_11_1_5;
  wire       [0:0]    shiftRows_port_state_out_11_1_6;
  wire       [0:0]    shiftRows_port_state_out_11_1_7;
  wire       [0:0]    shiftRows_port_state_out_12_0_0;
  wire       [0:0]    shiftRows_port_state_out_12_0_1;
  wire       [0:0]    shiftRows_port_state_out_12_0_2;
  wire       [0:0]    shiftRows_port_state_out_12_0_3;
  wire       [0:0]    shiftRows_port_state_out_12_0_4;
  wire       [0:0]    shiftRows_port_state_out_12_0_5;
  wire       [0:0]    shiftRows_port_state_out_12_0_6;
  wire       [0:0]    shiftRows_port_state_out_12_0_7;
  wire       [0:0]    shiftRows_port_state_out_12_1_0;
  wire       [0:0]    shiftRows_port_state_out_12_1_1;
  wire       [0:0]    shiftRows_port_state_out_12_1_2;
  wire       [0:0]    shiftRows_port_state_out_12_1_3;
  wire       [0:0]    shiftRows_port_state_out_12_1_4;
  wire       [0:0]    shiftRows_port_state_out_12_1_5;
  wire       [0:0]    shiftRows_port_state_out_12_1_6;
  wire       [0:0]    shiftRows_port_state_out_12_1_7;
  wire       [0:0]    shiftRows_port_state_out_13_0_0;
  wire       [0:0]    shiftRows_port_state_out_13_0_1;
  wire       [0:0]    shiftRows_port_state_out_13_0_2;
  wire       [0:0]    shiftRows_port_state_out_13_0_3;
  wire       [0:0]    shiftRows_port_state_out_13_0_4;
  wire       [0:0]    shiftRows_port_state_out_13_0_5;
  wire       [0:0]    shiftRows_port_state_out_13_0_6;
  wire       [0:0]    shiftRows_port_state_out_13_0_7;
  wire       [0:0]    shiftRows_port_state_out_13_1_0;
  wire       [0:0]    shiftRows_port_state_out_13_1_1;
  wire       [0:0]    shiftRows_port_state_out_13_1_2;
  wire       [0:0]    shiftRows_port_state_out_13_1_3;
  wire       [0:0]    shiftRows_port_state_out_13_1_4;
  wire       [0:0]    shiftRows_port_state_out_13_1_5;
  wire       [0:0]    shiftRows_port_state_out_13_1_6;
  wire       [0:0]    shiftRows_port_state_out_13_1_7;
  wire       [0:0]    shiftRows_port_state_out_14_0_0;
  wire       [0:0]    shiftRows_port_state_out_14_0_1;
  wire       [0:0]    shiftRows_port_state_out_14_0_2;
  wire       [0:0]    shiftRows_port_state_out_14_0_3;
  wire       [0:0]    shiftRows_port_state_out_14_0_4;
  wire       [0:0]    shiftRows_port_state_out_14_0_5;
  wire       [0:0]    shiftRows_port_state_out_14_0_6;
  wire       [0:0]    shiftRows_port_state_out_14_0_7;
  wire       [0:0]    shiftRows_port_state_out_14_1_0;
  wire       [0:0]    shiftRows_port_state_out_14_1_1;
  wire       [0:0]    shiftRows_port_state_out_14_1_2;
  wire       [0:0]    shiftRows_port_state_out_14_1_3;
  wire       [0:0]    shiftRows_port_state_out_14_1_4;
  wire       [0:0]    shiftRows_port_state_out_14_1_5;
  wire       [0:0]    shiftRows_port_state_out_14_1_6;
  wire       [0:0]    shiftRows_port_state_out_14_1_7;
  wire       [0:0]    shiftRows_port_state_out_15_0_0;
  wire       [0:0]    shiftRows_port_state_out_15_0_1;
  wire       [0:0]    shiftRows_port_state_out_15_0_2;
  wire       [0:0]    shiftRows_port_state_out_15_0_3;
  wire       [0:0]    shiftRows_port_state_out_15_0_4;
  wire       [0:0]    shiftRows_port_state_out_15_0_5;
  wire       [0:0]    shiftRows_port_state_out_15_0_6;
  wire       [0:0]    shiftRows_port_state_out_15_0_7;
  wire       [0:0]    shiftRows_port_state_out_15_1_0;
  wire       [0:0]    shiftRows_port_state_out_15_1_1;
  wire       [0:0]    shiftRows_port_state_out_15_1_2;
  wire       [0:0]    shiftRows_port_state_out_15_1_3;
  wire       [0:0]    shiftRows_port_state_out_15_1_4;
  wire       [0:0]    shiftRows_port_state_out_15_1_5;
  wire       [0:0]    shiftRows_port_state_out_15_1_6;
  wire       [0:0]    shiftRows_port_state_out_15_1_7;
  wire       [0:0]    mixColumns_port_state_out_0_0_0;
  wire       [0:0]    mixColumns_port_state_out_0_0_1;
  wire       [0:0]    mixColumns_port_state_out_0_0_2;
  wire       [0:0]    mixColumns_port_state_out_0_0_3;
  wire       [0:0]    mixColumns_port_state_out_0_0_4;
  wire       [0:0]    mixColumns_port_state_out_0_0_5;
  wire       [0:0]    mixColumns_port_state_out_0_0_6;
  wire       [0:0]    mixColumns_port_state_out_0_0_7;
  wire       [0:0]    mixColumns_port_state_out_0_1_0;
  wire       [0:0]    mixColumns_port_state_out_0_1_1;
  wire       [0:0]    mixColumns_port_state_out_0_1_2;
  wire       [0:0]    mixColumns_port_state_out_0_1_3;
  wire       [0:0]    mixColumns_port_state_out_0_1_4;
  wire       [0:0]    mixColumns_port_state_out_0_1_5;
  wire       [0:0]    mixColumns_port_state_out_0_1_6;
  wire       [0:0]    mixColumns_port_state_out_0_1_7;
  wire       [0:0]    mixColumns_port_state_out_1_0_0;
  wire       [0:0]    mixColumns_port_state_out_1_0_1;
  wire       [0:0]    mixColumns_port_state_out_1_0_2;
  wire       [0:0]    mixColumns_port_state_out_1_0_3;
  wire       [0:0]    mixColumns_port_state_out_1_0_4;
  wire       [0:0]    mixColumns_port_state_out_1_0_5;
  wire       [0:0]    mixColumns_port_state_out_1_0_6;
  wire       [0:0]    mixColumns_port_state_out_1_0_7;
  wire       [0:0]    mixColumns_port_state_out_1_1_0;
  wire       [0:0]    mixColumns_port_state_out_1_1_1;
  wire       [0:0]    mixColumns_port_state_out_1_1_2;
  wire       [0:0]    mixColumns_port_state_out_1_1_3;
  wire       [0:0]    mixColumns_port_state_out_1_1_4;
  wire       [0:0]    mixColumns_port_state_out_1_1_5;
  wire       [0:0]    mixColumns_port_state_out_1_1_6;
  wire       [0:0]    mixColumns_port_state_out_1_1_7;
  wire       [0:0]    mixColumns_port_state_out_2_0_0;
  wire       [0:0]    mixColumns_port_state_out_2_0_1;
  wire       [0:0]    mixColumns_port_state_out_2_0_2;
  wire       [0:0]    mixColumns_port_state_out_2_0_3;
  wire       [0:0]    mixColumns_port_state_out_2_0_4;
  wire       [0:0]    mixColumns_port_state_out_2_0_5;
  wire       [0:0]    mixColumns_port_state_out_2_0_6;
  wire       [0:0]    mixColumns_port_state_out_2_0_7;
  wire       [0:0]    mixColumns_port_state_out_2_1_0;
  wire       [0:0]    mixColumns_port_state_out_2_1_1;
  wire       [0:0]    mixColumns_port_state_out_2_1_2;
  wire       [0:0]    mixColumns_port_state_out_2_1_3;
  wire       [0:0]    mixColumns_port_state_out_2_1_4;
  wire       [0:0]    mixColumns_port_state_out_2_1_5;
  wire       [0:0]    mixColumns_port_state_out_2_1_6;
  wire       [0:0]    mixColumns_port_state_out_2_1_7;
  wire       [0:0]    mixColumns_port_state_out_3_0_0;
  wire       [0:0]    mixColumns_port_state_out_3_0_1;
  wire       [0:0]    mixColumns_port_state_out_3_0_2;
  wire       [0:0]    mixColumns_port_state_out_3_0_3;
  wire       [0:0]    mixColumns_port_state_out_3_0_4;
  wire       [0:0]    mixColumns_port_state_out_3_0_5;
  wire       [0:0]    mixColumns_port_state_out_3_0_6;
  wire       [0:0]    mixColumns_port_state_out_3_0_7;
  wire       [0:0]    mixColumns_port_state_out_3_1_0;
  wire       [0:0]    mixColumns_port_state_out_3_1_1;
  wire       [0:0]    mixColumns_port_state_out_3_1_2;
  wire       [0:0]    mixColumns_port_state_out_3_1_3;
  wire       [0:0]    mixColumns_port_state_out_3_1_4;
  wire       [0:0]    mixColumns_port_state_out_3_1_5;
  wire       [0:0]    mixColumns_port_state_out_3_1_6;
  wire       [0:0]    mixColumns_port_state_out_3_1_7;
  wire       [0:0]    mixColumns_port_state_out_4_0_0;
  wire       [0:0]    mixColumns_port_state_out_4_0_1;
  wire       [0:0]    mixColumns_port_state_out_4_0_2;
  wire       [0:0]    mixColumns_port_state_out_4_0_3;
  wire       [0:0]    mixColumns_port_state_out_4_0_4;
  wire       [0:0]    mixColumns_port_state_out_4_0_5;
  wire       [0:0]    mixColumns_port_state_out_4_0_6;
  wire       [0:0]    mixColumns_port_state_out_4_0_7;
  wire       [0:0]    mixColumns_port_state_out_4_1_0;
  wire       [0:0]    mixColumns_port_state_out_4_1_1;
  wire       [0:0]    mixColumns_port_state_out_4_1_2;
  wire       [0:0]    mixColumns_port_state_out_4_1_3;
  wire       [0:0]    mixColumns_port_state_out_4_1_4;
  wire       [0:0]    mixColumns_port_state_out_4_1_5;
  wire       [0:0]    mixColumns_port_state_out_4_1_6;
  wire       [0:0]    mixColumns_port_state_out_4_1_7;
  wire       [0:0]    mixColumns_port_state_out_5_0_0;
  wire       [0:0]    mixColumns_port_state_out_5_0_1;
  wire       [0:0]    mixColumns_port_state_out_5_0_2;
  wire       [0:0]    mixColumns_port_state_out_5_0_3;
  wire       [0:0]    mixColumns_port_state_out_5_0_4;
  wire       [0:0]    mixColumns_port_state_out_5_0_5;
  wire       [0:0]    mixColumns_port_state_out_5_0_6;
  wire       [0:0]    mixColumns_port_state_out_5_0_7;
  wire       [0:0]    mixColumns_port_state_out_5_1_0;
  wire       [0:0]    mixColumns_port_state_out_5_1_1;
  wire       [0:0]    mixColumns_port_state_out_5_1_2;
  wire       [0:0]    mixColumns_port_state_out_5_1_3;
  wire       [0:0]    mixColumns_port_state_out_5_1_4;
  wire       [0:0]    mixColumns_port_state_out_5_1_5;
  wire       [0:0]    mixColumns_port_state_out_5_1_6;
  wire       [0:0]    mixColumns_port_state_out_5_1_7;
  wire       [0:0]    mixColumns_port_state_out_6_0_0;
  wire       [0:0]    mixColumns_port_state_out_6_0_1;
  wire       [0:0]    mixColumns_port_state_out_6_0_2;
  wire       [0:0]    mixColumns_port_state_out_6_0_3;
  wire       [0:0]    mixColumns_port_state_out_6_0_4;
  wire       [0:0]    mixColumns_port_state_out_6_0_5;
  wire       [0:0]    mixColumns_port_state_out_6_0_6;
  wire       [0:0]    mixColumns_port_state_out_6_0_7;
  wire       [0:0]    mixColumns_port_state_out_6_1_0;
  wire       [0:0]    mixColumns_port_state_out_6_1_1;
  wire       [0:0]    mixColumns_port_state_out_6_1_2;
  wire       [0:0]    mixColumns_port_state_out_6_1_3;
  wire       [0:0]    mixColumns_port_state_out_6_1_4;
  wire       [0:0]    mixColumns_port_state_out_6_1_5;
  wire       [0:0]    mixColumns_port_state_out_6_1_6;
  wire       [0:0]    mixColumns_port_state_out_6_1_7;
  wire       [0:0]    mixColumns_port_state_out_7_0_0;
  wire       [0:0]    mixColumns_port_state_out_7_0_1;
  wire       [0:0]    mixColumns_port_state_out_7_0_2;
  wire       [0:0]    mixColumns_port_state_out_7_0_3;
  wire       [0:0]    mixColumns_port_state_out_7_0_4;
  wire       [0:0]    mixColumns_port_state_out_7_0_5;
  wire       [0:0]    mixColumns_port_state_out_7_0_6;
  wire       [0:0]    mixColumns_port_state_out_7_0_7;
  wire       [0:0]    mixColumns_port_state_out_7_1_0;
  wire       [0:0]    mixColumns_port_state_out_7_1_1;
  wire       [0:0]    mixColumns_port_state_out_7_1_2;
  wire       [0:0]    mixColumns_port_state_out_7_1_3;
  wire       [0:0]    mixColumns_port_state_out_7_1_4;
  wire       [0:0]    mixColumns_port_state_out_7_1_5;
  wire       [0:0]    mixColumns_port_state_out_7_1_6;
  wire       [0:0]    mixColumns_port_state_out_7_1_7;
  wire       [0:0]    mixColumns_port_state_out_8_0_0;
  wire       [0:0]    mixColumns_port_state_out_8_0_1;
  wire       [0:0]    mixColumns_port_state_out_8_0_2;
  wire       [0:0]    mixColumns_port_state_out_8_0_3;
  wire       [0:0]    mixColumns_port_state_out_8_0_4;
  wire       [0:0]    mixColumns_port_state_out_8_0_5;
  wire       [0:0]    mixColumns_port_state_out_8_0_6;
  wire       [0:0]    mixColumns_port_state_out_8_0_7;
  wire       [0:0]    mixColumns_port_state_out_8_1_0;
  wire       [0:0]    mixColumns_port_state_out_8_1_1;
  wire       [0:0]    mixColumns_port_state_out_8_1_2;
  wire       [0:0]    mixColumns_port_state_out_8_1_3;
  wire       [0:0]    mixColumns_port_state_out_8_1_4;
  wire       [0:0]    mixColumns_port_state_out_8_1_5;
  wire       [0:0]    mixColumns_port_state_out_8_1_6;
  wire       [0:0]    mixColumns_port_state_out_8_1_7;
  wire       [0:0]    mixColumns_port_state_out_9_0_0;
  wire       [0:0]    mixColumns_port_state_out_9_0_1;
  wire       [0:0]    mixColumns_port_state_out_9_0_2;
  wire       [0:0]    mixColumns_port_state_out_9_0_3;
  wire       [0:0]    mixColumns_port_state_out_9_0_4;
  wire       [0:0]    mixColumns_port_state_out_9_0_5;
  wire       [0:0]    mixColumns_port_state_out_9_0_6;
  wire       [0:0]    mixColumns_port_state_out_9_0_7;
  wire       [0:0]    mixColumns_port_state_out_9_1_0;
  wire       [0:0]    mixColumns_port_state_out_9_1_1;
  wire       [0:0]    mixColumns_port_state_out_9_1_2;
  wire       [0:0]    mixColumns_port_state_out_9_1_3;
  wire       [0:0]    mixColumns_port_state_out_9_1_4;
  wire       [0:0]    mixColumns_port_state_out_9_1_5;
  wire       [0:0]    mixColumns_port_state_out_9_1_6;
  wire       [0:0]    mixColumns_port_state_out_9_1_7;
  wire       [0:0]    mixColumns_port_state_out_10_0_0;
  wire       [0:0]    mixColumns_port_state_out_10_0_1;
  wire       [0:0]    mixColumns_port_state_out_10_0_2;
  wire       [0:0]    mixColumns_port_state_out_10_0_3;
  wire       [0:0]    mixColumns_port_state_out_10_0_4;
  wire       [0:0]    mixColumns_port_state_out_10_0_5;
  wire       [0:0]    mixColumns_port_state_out_10_0_6;
  wire       [0:0]    mixColumns_port_state_out_10_0_7;
  wire       [0:0]    mixColumns_port_state_out_10_1_0;
  wire       [0:0]    mixColumns_port_state_out_10_1_1;
  wire       [0:0]    mixColumns_port_state_out_10_1_2;
  wire       [0:0]    mixColumns_port_state_out_10_1_3;
  wire       [0:0]    mixColumns_port_state_out_10_1_4;
  wire       [0:0]    mixColumns_port_state_out_10_1_5;
  wire       [0:0]    mixColumns_port_state_out_10_1_6;
  wire       [0:0]    mixColumns_port_state_out_10_1_7;
  wire       [0:0]    mixColumns_port_state_out_11_0_0;
  wire       [0:0]    mixColumns_port_state_out_11_0_1;
  wire       [0:0]    mixColumns_port_state_out_11_0_2;
  wire       [0:0]    mixColumns_port_state_out_11_0_3;
  wire       [0:0]    mixColumns_port_state_out_11_0_4;
  wire       [0:0]    mixColumns_port_state_out_11_0_5;
  wire       [0:0]    mixColumns_port_state_out_11_0_6;
  wire       [0:0]    mixColumns_port_state_out_11_0_7;
  wire       [0:0]    mixColumns_port_state_out_11_1_0;
  wire       [0:0]    mixColumns_port_state_out_11_1_1;
  wire       [0:0]    mixColumns_port_state_out_11_1_2;
  wire       [0:0]    mixColumns_port_state_out_11_1_3;
  wire       [0:0]    mixColumns_port_state_out_11_1_4;
  wire       [0:0]    mixColumns_port_state_out_11_1_5;
  wire       [0:0]    mixColumns_port_state_out_11_1_6;
  wire       [0:0]    mixColumns_port_state_out_11_1_7;
  wire       [0:0]    mixColumns_port_state_out_12_0_0;
  wire       [0:0]    mixColumns_port_state_out_12_0_1;
  wire       [0:0]    mixColumns_port_state_out_12_0_2;
  wire       [0:0]    mixColumns_port_state_out_12_0_3;
  wire       [0:0]    mixColumns_port_state_out_12_0_4;
  wire       [0:0]    mixColumns_port_state_out_12_0_5;
  wire       [0:0]    mixColumns_port_state_out_12_0_6;
  wire       [0:0]    mixColumns_port_state_out_12_0_7;
  wire       [0:0]    mixColumns_port_state_out_12_1_0;
  wire       [0:0]    mixColumns_port_state_out_12_1_1;
  wire       [0:0]    mixColumns_port_state_out_12_1_2;
  wire       [0:0]    mixColumns_port_state_out_12_1_3;
  wire       [0:0]    mixColumns_port_state_out_12_1_4;
  wire       [0:0]    mixColumns_port_state_out_12_1_5;
  wire       [0:0]    mixColumns_port_state_out_12_1_6;
  wire       [0:0]    mixColumns_port_state_out_12_1_7;
  wire       [0:0]    mixColumns_port_state_out_13_0_0;
  wire       [0:0]    mixColumns_port_state_out_13_0_1;
  wire       [0:0]    mixColumns_port_state_out_13_0_2;
  wire       [0:0]    mixColumns_port_state_out_13_0_3;
  wire       [0:0]    mixColumns_port_state_out_13_0_4;
  wire       [0:0]    mixColumns_port_state_out_13_0_5;
  wire       [0:0]    mixColumns_port_state_out_13_0_6;
  wire       [0:0]    mixColumns_port_state_out_13_0_7;
  wire       [0:0]    mixColumns_port_state_out_13_1_0;
  wire       [0:0]    mixColumns_port_state_out_13_1_1;
  wire       [0:0]    mixColumns_port_state_out_13_1_2;
  wire       [0:0]    mixColumns_port_state_out_13_1_3;
  wire       [0:0]    mixColumns_port_state_out_13_1_4;
  wire       [0:0]    mixColumns_port_state_out_13_1_5;
  wire       [0:0]    mixColumns_port_state_out_13_1_6;
  wire       [0:0]    mixColumns_port_state_out_13_1_7;
  wire       [0:0]    mixColumns_port_state_out_14_0_0;
  wire       [0:0]    mixColumns_port_state_out_14_0_1;
  wire       [0:0]    mixColumns_port_state_out_14_0_2;
  wire       [0:0]    mixColumns_port_state_out_14_0_3;
  wire       [0:0]    mixColumns_port_state_out_14_0_4;
  wire       [0:0]    mixColumns_port_state_out_14_0_5;
  wire       [0:0]    mixColumns_port_state_out_14_0_6;
  wire       [0:0]    mixColumns_port_state_out_14_0_7;
  wire       [0:0]    mixColumns_port_state_out_14_1_0;
  wire       [0:0]    mixColumns_port_state_out_14_1_1;
  wire       [0:0]    mixColumns_port_state_out_14_1_2;
  wire       [0:0]    mixColumns_port_state_out_14_1_3;
  wire       [0:0]    mixColumns_port_state_out_14_1_4;
  wire       [0:0]    mixColumns_port_state_out_14_1_5;
  wire       [0:0]    mixColumns_port_state_out_14_1_6;
  wire       [0:0]    mixColumns_port_state_out_14_1_7;
  wire       [0:0]    mixColumns_port_state_out_15_0_0;
  wire       [0:0]    mixColumns_port_state_out_15_0_1;
  wire       [0:0]    mixColumns_port_state_out_15_0_2;
  wire       [0:0]    mixColumns_port_state_out_15_0_3;
  wire       [0:0]    mixColumns_port_state_out_15_0_4;
  wire       [0:0]    mixColumns_port_state_out_15_0_5;
  wire       [0:0]    mixColumns_port_state_out_15_0_6;
  wire       [0:0]    mixColumns_port_state_out_15_0_7;
  wire       [0:0]    mixColumns_port_state_out_15_1_0;
  wire       [0:0]    mixColumns_port_state_out_15_1_1;
  wire       [0:0]    mixColumns_port_state_out_15_1_2;
  wire       [0:0]    mixColumns_port_state_out_15_1_3;
  wire       [0:0]    mixColumns_port_state_out_15_1_4;
  wire       [0:0]    mixColumns_port_state_out_15_1_5;
  wire       [0:0]    mixColumns_port_state_out_15_1_6;
  wire       [0:0]    mixColumns_port_state_out_15_1_7;
  wire       [0:0]    subBytes_out_0_0_0;
  wire       [0:0]    subBytes_out_0_0_1;
  wire       [0:0]    subBytes_out_0_0_2;
  wire       [0:0]    subBytes_out_0_0_3;
  wire       [0:0]    subBytes_out_0_0_4;
  wire       [0:0]    subBytes_out_0_0_5;
  wire       [0:0]    subBytes_out_0_0_6;
  wire       [0:0]    subBytes_out_0_0_7;
  wire       [0:0]    subBytes_out_0_1_0;
  wire       [0:0]    subBytes_out_0_1_1;
  wire       [0:0]    subBytes_out_0_1_2;
  wire       [0:0]    subBytes_out_0_1_3;
  wire       [0:0]    subBytes_out_0_1_4;
  wire       [0:0]    subBytes_out_0_1_5;
  wire       [0:0]    subBytes_out_0_1_6;
  wire       [0:0]    subBytes_out_0_1_7;
  wire       [0:0]    subBytes_out_1_0_0;
  wire       [0:0]    subBytes_out_1_0_1;
  wire       [0:0]    subBytes_out_1_0_2;
  wire       [0:0]    subBytes_out_1_0_3;
  wire       [0:0]    subBytes_out_1_0_4;
  wire       [0:0]    subBytes_out_1_0_5;
  wire       [0:0]    subBytes_out_1_0_6;
  wire       [0:0]    subBytes_out_1_0_7;
  wire       [0:0]    subBytes_out_1_1_0;
  wire       [0:0]    subBytes_out_1_1_1;
  wire       [0:0]    subBytes_out_1_1_2;
  wire       [0:0]    subBytes_out_1_1_3;
  wire       [0:0]    subBytes_out_1_1_4;
  wire       [0:0]    subBytes_out_1_1_5;
  wire       [0:0]    subBytes_out_1_1_6;
  wire       [0:0]    subBytes_out_1_1_7;
  wire       [0:0]    subBytes_out_2_0_0;
  wire       [0:0]    subBytes_out_2_0_1;
  wire       [0:0]    subBytes_out_2_0_2;
  wire       [0:0]    subBytes_out_2_0_3;
  wire       [0:0]    subBytes_out_2_0_4;
  wire       [0:0]    subBytes_out_2_0_5;
  wire       [0:0]    subBytes_out_2_0_6;
  wire       [0:0]    subBytes_out_2_0_7;
  wire       [0:0]    subBytes_out_2_1_0;
  wire       [0:0]    subBytes_out_2_1_1;
  wire       [0:0]    subBytes_out_2_1_2;
  wire       [0:0]    subBytes_out_2_1_3;
  wire       [0:0]    subBytes_out_2_1_4;
  wire       [0:0]    subBytes_out_2_1_5;
  wire       [0:0]    subBytes_out_2_1_6;
  wire       [0:0]    subBytes_out_2_1_7;
  wire       [0:0]    subBytes_out_3_0_0;
  wire       [0:0]    subBytes_out_3_0_1;
  wire       [0:0]    subBytes_out_3_0_2;
  wire       [0:0]    subBytes_out_3_0_3;
  wire       [0:0]    subBytes_out_3_0_4;
  wire       [0:0]    subBytes_out_3_0_5;
  wire       [0:0]    subBytes_out_3_0_6;
  wire       [0:0]    subBytes_out_3_0_7;
  wire       [0:0]    subBytes_out_3_1_0;
  wire       [0:0]    subBytes_out_3_1_1;
  wire       [0:0]    subBytes_out_3_1_2;
  wire       [0:0]    subBytes_out_3_1_3;
  wire       [0:0]    subBytes_out_3_1_4;
  wire       [0:0]    subBytes_out_3_1_5;
  wire       [0:0]    subBytes_out_3_1_6;
  wire       [0:0]    subBytes_out_3_1_7;
  wire       [0:0]    subBytes_out_4_0_0;
  wire       [0:0]    subBytes_out_4_0_1;
  wire       [0:0]    subBytes_out_4_0_2;
  wire       [0:0]    subBytes_out_4_0_3;
  wire       [0:0]    subBytes_out_4_0_4;
  wire       [0:0]    subBytes_out_4_0_5;
  wire       [0:0]    subBytes_out_4_0_6;
  wire       [0:0]    subBytes_out_4_0_7;
  wire       [0:0]    subBytes_out_4_1_0;
  wire       [0:0]    subBytes_out_4_1_1;
  wire       [0:0]    subBytes_out_4_1_2;
  wire       [0:0]    subBytes_out_4_1_3;
  wire       [0:0]    subBytes_out_4_1_4;
  wire       [0:0]    subBytes_out_4_1_5;
  wire       [0:0]    subBytes_out_4_1_6;
  wire       [0:0]    subBytes_out_4_1_7;
  wire       [0:0]    subBytes_out_5_0_0;
  wire       [0:0]    subBytes_out_5_0_1;
  wire       [0:0]    subBytes_out_5_0_2;
  wire       [0:0]    subBytes_out_5_0_3;
  wire       [0:0]    subBytes_out_5_0_4;
  wire       [0:0]    subBytes_out_5_0_5;
  wire       [0:0]    subBytes_out_5_0_6;
  wire       [0:0]    subBytes_out_5_0_7;
  wire       [0:0]    subBytes_out_5_1_0;
  wire       [0:0]    subBytes_out_5_1_1;
  wire       [0:0]    subBytes_out_5_1_2;
  wire       [0:0]    subBytes_out_5_1_3;
  wire       [0:0]    subBytes_out_5_1_4;
  wire       [0:0]    subBytes_out_5_1_5;
  wire       [0:0]    subBytes_out_5_1_6;
  wire       [0:0]    subBytes_out_5_1_7;
  wire       [0:0]    subBytes_out_6_0_0;
  wire       [0:0]    subBytes_out_6_0_1;
  wire       [0:0]    subBytes_out_6_0_2;
  wire       [0:0]    subBytes_out_6_0_3;
  wire       [0:0]    subBytes_out_6_0_4;
  wire       [0:0]    subBytes_out_6_0_5;
  wire       [0:0]    subBytes_out_6_0_6;
  wire       [0:0]    subBytes_out_6_0_7;
  wire       [0:0]    subBytes_out_6_1_0;
  wire       [0:0]    subBytes_out_6_1_1;
  wire       [0:0]    subBytes_out_6_1_2;
  wire       [0:0]    subBytes_out_6_1_3;
  wire       [0:0]    subBytes_out_6_1_4;
  wire       [0:0]    subBytes_out_6_1_5;
  wire       [0:0]    subBytes_out_6_1_6;
  wire       [0:0]    subBytes_out_6_1_7;
  wire       [0:0]    subBytes_out_7_0_0;
  wire       [0:0]    subBytes_out_7_0_1;
  wire       [0:0]    subBytes_out_7_0_2;
  wire       [0:0]    subBytes_out_7_0_3;
  wire       [0:0]    subBytes_out_7_0_4;
  wire       [0:0]    subBytes_out_7_0_5;
  wire       [0:0]    subBytes_out_7_0_6;
  wire       [0:0]    subBytes_out_7_0_7;
  wire       [0:0]    subBytes_out_7_1_0;
  wire       [0:0]    subBytes_out_7_1_1;
  wire       [0:0]    subBytes_out_7_1_2;
  wire       [0:0]    subBytes_out_7_1_3;
  wire       [0:0]    subBytes_out_7_1_4;
  wire       [0:0]    subBytes_out_7_1_5;
  wire       [0:0]    subBytes_out_7_1_6;
  wire       [0:0]    subBytes_out_7_1_7;
  wire       [0:0]    subBytes_out_8_0_0;
  wire       [0:0]    subBytes_out_8_0_1;
  wire       [0:0]    subBytes_out_8_0_2;
  wire       [0:0]    subBytes_out_8_0_3;
  wire       [0:0]    subBytes_out_8_0_4;
  wire       [0:0]    subBytes_out_8_0_5;
  wire       [0:0]    subBytes_out_8_0_6;
  wire       [0:0]    subBytes_out_8_0_7;
  wire       [0:0]    subBytes_out_8_1_0;
  wire       [0:0]    subBytes_out_8_1_1;
  wire       [0:0]    subBytes_out_8_1_2;
  wire       [0:0]    subBytes_out_8_1_3;
  wire       [0:0]    subBytes_out_8_1_4;
  wire       [0:0]    subBytes_out_8_1_5;
  wire       [0:0]    subBytes_out_8_1_6;
  wire       [0:0]    subBytes_out_8_1_7;
  wire       [0:0]    subBytes_out_9_0_0;
  wire       [0:0]    subBytes_out_9_0_1;
  wire       [0:0]    subBytes_out_9_0_2;
  wire       [0:0]    subBytes_out_9_0_3;
  wire       [0:0]    subBytes_out_9_0_4;
  wire       [0:0]    subBytes_out_9_0_5;
  wire       [0:0]    subBytes_out_9_0_6;
  wire       [0:0]    subBytes_out_9_0_7;
  wire       [0:0]    subBytes_out_9_1_0;
  wire       [0:0]    subBytes_out_9_1_1;
  wire       [0:0]    subBytes_out_9_1_2;
  wire       [0:0]    subBytes_out_9_1_3;
  wire       [0:0]    subBytes_out_9_1_4;
  wire       [0:0]    subBytes_out_9_1_5;
  wire       [0:0]    subBytes_out_9_1_6;
  wire       [0:0]    subBytes_out_9_1_7;
  wire       [0:0]    subBytes_out_10_0_0;
  wire       [0:0]    subBytes_out_10_0_1;
  wire       [0:0]    subBytes_out_10_0_2;
  wire       [0:0]    subBytes_out_10_0_3;
  wire       [0:0]    subBytes_out_10_0_4;
  wire       [0:0]    subBytes_out_10_0_5;
  wire       [0:0]    subBytes_out_10_0_6;
  wire       [0:0]    subBytes_out_10_0_7;
  wire       [0:0]    subBytes_out_10_1_0;
  wire       [0:0]    subBytes_out_10_1_1;
  wire       [0:0]    subBytes_out_10_1_2;
  wire       [0:0]    subBytes_out_10_1_3;
  wire       [0:0]    subBytes_out_10_1_4;
  wire       [0:0]    subBytes_out_10_1_5;
  wire       [0:0]    subBytes_out_10_1_6;
  wire       [0:0]    subBytes_out_10_1_7;
  wire       [0:0]    subBytes_out_11_0_0;
  wire       [0:0]    subBytes_out_11_0_1;
  wire       [0:0]    subBytes_out_11_0_2;
  wire       [0:0]    subBytes_out_11_0_3;
  wire       [0:0]    subBytes_out_11_0_4;
  wire       [0:0]    subBytes_out_11_0_5;
  wire       [0:0]    subBytes_out_11_0_6;
  wire       [0:0]    subBytes_out_11_0_7;
  wire       [0:0]    subBytes_out_11_1_0;
  wire       [0:0]    subBytes_out_11_1_1;
  wire       [0:0]    subBytes_out_11_1_2;
  wire       [0:0]    subBytes_out_11_1_3;
  wire       [0:0]    subBytes_out_11_1_4;
  wire       [0:0]    subBytes_out_11_1_5;
  wire       [0:0]    subBytes_out_11_1_6;
  wire       [0:0]    subBytes_out_11_1_7;
  wire       [0:0]    subBytes_out_12_0_0;
  wire       [0:0]    subBytes_out_12_0_1;
  wire       [0:0]    subBytes_out_12_0_2;
  wire       [0:0]    subBytes_out_12_0_3;
  wire       [0:0]    subBytes_out_12_0_4;
  wire       [0:0]    subBytes_out_12_0_5;
  wire       [0:0]    subBytes_out_12_0_6;
  wire       [0:0]    subBytes_out_12_0_7;
  wire       [0:0]    subBytes_out_12_1_0;
  wire       [0:0]    subBytes_out_12_1_1;
  wire       [0:0]    subBytes_out_12_1_2;
  wire       [0:0]    subBytes_out_12_1_3;
  wire       [0:0]    subBytes_out_12_1_4;
  wire       [0:0]    subBytes_out_12_1_5;
  wire       [0:0]    subBytes_out_12_1_6;
  wire       [0:0]    subBytes_out_12_1_7;
  wire       [0:0]    subBytes_out_13_0_0;
  wire       [0:0]    subBytes_out_13_0_1;
  wire       [0:0]    subBytes_out_13_0_2;
  wire       [0:0]    subBytes_out_13_0_3;
  wire       [0:0]    subBytes_out_13_0_4;
  wire       [0:0]    subBytes_out_13_0_5;
  wire       [0:0]    subBytes_out_13_0_6;
  wire       [0:0]    subBytes_out_13_0_7;
  wire       [0:0]    subBytes_out_13_1_0;
  wire       [0:0]    subBytes_out_13_1_1;
  wire       [0:0]    subBytes_out_13_1_2;
  wire       [0:0]    subBytes_out_13_1_3;
  wire       [0:0]    subBytes_out_13_1_4;
  wire       [0:0]    subBytes_out_13_1_5;
  wire       [0:0]    subBytes_out_13_1_6;
  wire       [0:0]    subBytes_out_13_1_7;
  wire       [0:0]    subBytes_out_14_0_0;
  wire       [0:0]    subBytes_out_14_0_1;
  wire       [0:0]    subBytes_out_14_0_2;
  wire       [0:0]    subBytes_out_14_0_3;
  wire       [0:0]    subBytes_out_14_0_4;
  wire       [0:0]    subBytes_out_14_0_5;
  wire       [0:0]    subBytes_out_14_0_6;
  wire       [0:0]    subBytes_out_14_0_7;
  wire       [0:0]    subBytes_out_14_1_0;
  wire       [0:0]    subBytes_out_14_1_1;
  wire       [0:0]    subBytes_out_14_1_2;
  wire       [0:0]    subBytes_out_14_1_3;
  wire       [0:0]    subBytes_out_14_1_4;
  wire       [0:0]    subBytes_out_14_1_5;
  wire       [0:0]    subBytes_out_14_1_6;
  wire       [0:0]    subBytes_out_14_1_7;
  wire       [0:0]    subBytes_out_15_0_0;
  wire       [0:0]    subBytes_out_15_0_1;
  wire       [0:0]    subBytes_out_15_0_2;
  wire       [0:0]    subBytes_out_15_0_3;
  wire       [0:0]    subBytes_out_15_0_4;
  wire       [0:0]    subBytes_out_15_0_5;
  wire       [0:0]    subBytes_out_15_0_6;
  wire       [0:0]    subBytes_out_15_0_7;
  wire       [0:0]    subBytes_out_15_1_0;
  wire       [0:0]    subBytes_out_15_1_1;
  wire       [0:0]    subBytes_out_15_1_2;
  wire       [0:0]    subBytes_out_15_1_3;
  wire       [0:0]    subBytes_out_15_1_4;
  wire       [0:0]    subBytes_out_15_1_5;
  wire       [0:0]    subBytes_out_15_1_6;
  wire       [0:0]    subBytes_out_15_1_7;
  reg        [0:0]    roundReg_0_0_0;
  reg        [0:0]    roundReg_0_0_1;
  reg        [0:0]    roundReg_0_0_2;
  reg        [0:0]    roundReg_0_0_3;
  reg        [0:0]    roundReg_0_0_4;
  reg        [0:0]    roundReg_0_0_5;
  reg        [0:0]    roundReg_0_0_6;
  reg        [0:0]    roundReg_0_0_7;
  reg        [0:0]    roundReg_0_1_0;
  reg        [0:0]    roundReg_0_1_1;
  reg        [0:0]    roundReg_0_1_2;
  reg        [0:0]    roundReg_0_1_3;
  reg        [0:0]    roundReg_0_1_4;
  reg        [0:0]    roundReg_0_1_5;
  reg        [0:0]    roundReg_0_1_6;
  reg        [0:0]    roundReg_0_1_7;
  reg        [0:0]    roundReg_1_0_0;
  reg        [0:0]    roundReg_1_0_1;
  reg        [0:0]    roundReg_1_0_2;
  reg        [0:0]    roundReg_1_0_3;
  reg        [0:0]    roundReg_1_0_4;
  reg        [0:0]    roundReg_1_0_5;
  reg        [0:0]    roundReg_1_0_6;
  reg        [0:0]    roundReg_1_0_7;
  reg        [0:0]    roundReg_1_1_0;
  reg        [0:0]    roundReg_1_1_1;
  reg        [0:0]    roundReg_1_1_2;
  reg        [0:0]    roundReg_1_1_3;
  reg        [0:0]    roundReg_1_1_4;
  reg        [0:0]    roundReg_1_1_5;
  reg        [0:0]    roundReg_1_1_6;
  reg        [0:0]    roundReg_1_1_7;
  reg        [0:0]    roundReg_2_0_0;
  reg        [0:0]    roundReg_2_0_1;
  reg        [0:0]    roundReg_2_0_2;
  reg        [0:0]    roundReg_2_0_3;
  reg        [0:0]    roundReg_2_0_4;
  reg        [0:0]    roundReg_2_0_5;
  reg        [0:0]    roundReg_2_0_6;
  reg        [0:0]    roundReg_2_0_7;
  reg        [0:0]    roundReg_2_1_0;
  reg        [0:0]    roundReg_2_1_1;
  reg        [0:0]    roundReg_2_1_2;
  reg        [0:0]    roundReg_2_1_3;
  reg        [0:0]    roundReg_2_1_4;
  reg        [0:0]    roundReg_2_1_5;
  reg        [0:0]    roundReg_2_1_6;
  reg        [0:0]    roundReg_2_1_7;
  reg        [0:0]    roundReg_3_0_0;
  reg        [0:0]    roundReg_3_0_1;
  reg        [0:0]    roundReg_3_0_2;
  reg        [0:0]    roundReg_3_0_3;
  reg        [0:0]    roundReg_3_0_4;
  reg        [0:0]    roundReg_3_0_5;
  reg        [0:0]    roundReg_3_0_6;
  reg        [0:0]    roundReg_3_0_7;
  reg        [0:0]    roundReg_3_1_0;
  reg        [0:0]    roundReg_3_1_1;
  reg        [0:0]    roundReg_3_1_2;
  reg        [0:0]    roundReg_3_1_3;
  reg        [0:0]    roundReg_3_1_4;
  reg        [0:0]    roundReg_3_1_5;
  reg        [0:0]    roundReg_3_1_6;
  reg        [0:0]    roundReg_3_1_7;
  reg        [0:0]    roundReg_4_0_0;
  reg        [0:0]    roundReg_4_0_1;
  reg        [0:0]    roundReg_4_0_2;
  reg        [0:0]    roundReg_4_0_3;
  reg        [0:0]    roundReg_4_0_4;
  reg        [0:0]    roundReg_4_0_5;
  reg        [0:0]    roundReg_4_0_6;
  reg        [0:0]    roundReg_4_0_7;
  reg        [0:0]    roundReg_4_1_0;
  reg        [0:0]    roundReg_4_1_1;
  reg        [0:0]    roundReg_4_1_2;
  reg        [0:0]    roundReg_4_1_3;
  reg        [0:0]    roundReg_4_1_4;
  reg        [0:0]    roundReg_4_1_5;
  reg        [0:0]    roundReg_4_1_6;
  reg        [0:0]    roundReg_4_1_7;
  reg        [0:0]    roundReg_5_0_0;
  reg        [0:0]    roundReg_5_0_1;
  reg        [0:0]    roundReg_5_0_2;
  reg        [0:0]    roundReg_5_0_3;
  reg        [0:0]    roundReg_5_0_4;
  reg        [0:0]    roundReg_5_0_5;
  reg        [0:0]    roundReg_5_0_6;
  reg        [0:0]    roundReg_5_0_7;
  reg        [0:0]    roundReg_5_1_0;
  reg        [0:0]    roundReg_5_1_1;
  reg        [0:0]    roundReg_5_1_2;
  reg        [0:0]    roundReg_5_1_3;
  reg        [0:0]    roundReg_5_1_4;
  reg        [0:0]    roundReg_5_1_5;
  reg        [0:0]    roundReg_5_1_6;
  reg        [0:0]    roundReg_5_1_7;
  reg        [0:0]    roundReg_6_0_0;
  reg        [0:0]    roundReg_6_0_1;
  reg        [0:0]    roundReg_6_0_2;
  reg        [0:0]    roundReg_6_0_3;
  reg        [0:0]    roundReg_6_0_4;
  reg        [0:0]    roundReg_6_0_5;
  reg        [0:0]    roundReg_6_0_6;
  reg        [0:0]    roundReg_6_0_7;
  reg        [0:0]    roundReg_6_1_0;
  reg        [0:0]    roundReg_6_1_1;
  reg        [0:0]    roundReg_6_1_2;
  reg        [0:0]    roundReg_6_1_3;
  reg        [0:0]    roundReg_6_1_4;
  reg        [0:0]    roundReg_6_1_5;
  reg        [0:0]    roundReg_6_1_6;
  reg        [0:0]    roundReg_6_1_7;
  reg        [0:0]    roundReg_7_0_0;
  reg        [0:0]    roundReg_7_0_1;
  reg        [0:0]    roundReg_7_0_2;
  reg        [0:0]    roundReg_7_0_3;
  reg        [0:0]    roundReg_7_0_4;
  reg        [0:0]    roundReg_7_0_5;
  reg        [0:0]    roundReg_7_0_6;
  reg        [0:0]    roundReg_7_0_7;
  reg        [0:0]    roundReg_7_1_0;
  reg        [0:0]    roundReg_7_1_1;
  reg        [0:0]    roundReg_7_1_2;
  reg        [0:0]    roundReg_7_1_3;
  reg        [0:0]    roundReg_7_1_4;
  reg        [0:0]    roundReg_7_1_5;
  reg        [0:0]    roundReg_7_1_6;
  reg        [0:0]    roundReg_7_1_7;
  reg        [0:0]    roundReg_8_0_0;
  reg        [0:0]    roundReg_8_0_1;
  reg        [0:0]    roundReg_8_0_2;
  reg        [0:0]    roundReg_8_0_3;
  reg        [0:0]    roundReg_8_0_4;
  reg        [0:0]    roundReg_8_0_5;
  reg        [0:0]    roundReg_8_0_6;
  reg        [0:0]    roundReg_8_0_7;
  reg        [0:0]    roundReg_8_1_0;
  reg        [0:0]    roundReg_8_1_1;
  reg        [0:0]    roundReg_8_1_2;
  reg        [0:0]    roundReg_8_1_3;
  reg        [0:0]    roundReg_8_1_4;
  reg        [0:0]    roundReg_8_1_5;
  reg        [0:0]    roundReg_8_1_6;
  reg        [0:0]    roundReg_8_1_7;
  reg        [0:0]    roundReg_9_0_0;
  reg        [0:0]    roundReg_9_0_1;
  reg        [0:0]    roundReg_9_0_2;
  reg        [0:0]    roundReg_9_0_3;
  reg        [0:0]    roundReg_9_0_4;
  reg        [0:0]    roundReg_9_0_5;
  reg        [0:0]    roundReg_9_0_6;
  reg        [0:0]    roundReg_9_0_7;
  reg        [0:0]    roundReg_9_1_0;
  reg        [0:0]    roundReg_9_1_1;
  reg        [0:0]    roundReg_9_1_2;
  reg        [0:0]    roundReg_9_1_3;
  reg        [0:0]    roundReg_9_1_4;
  reg        [0:0]    roundReg_9_1_5;
  reg        [0:0]    roundReg_9_1_6;
  reg        [0:0]    roundReg_9_1_7;
  reg        [0:0]    roundReg_10_0_0;
  reg        [0:0]    roundReg_10_0_1;
  reg        [0:0]    roundReg_10_0_2;
  reg        [0:0]    roundReg_10_0_3;
  reg        [0:0]    roundReg_10_0_4;
  reg        [0:0]    roundReg_10_0_5;
  reg        [0:0]    roundReg_10_0_6;
  reg        [0:0]    roundReg_10_0_7;
  reg        [0:0]    roundReg_10_1_0;
  reg        [0:0]    roundReg_10_1_1;
  reg        [0:0]    roundReg_10_1_2;
  reg        [0:0]    roundReg_10_1_3;
  reg        [0:0]    roundReg_10_1_4;
  reg        [0:0]    roundReg_10_1_5;
  reg        [0:0]    roundReg_10_1_6;
  reg        [0:0]    roundReg_10_1_7;
  reg        [0:0]    roundReg_11_0_0;
  reg        [0:0]    roundReg_11_0_1;
  reg        [0:0]    roundReg_11_0_2;
  reg        [0:0]    roundReg_11_0_3;
  reg        [0:0]    roundReg_11_0_4;
  reg        [0:0]    roundReg_11_0_5;
  reg        [0:0]    roundReg_11_0_6;
  reg        [0:0]    roundReg_11_0_7;
  reg        [0:0]    roundReg_11_1_0;
  reg        [0:0]    roundReg_11_1_1;
  reg        [0:0]    roundReg_11_1_2;
  reg        [0:0]    roundReg_11_1_3;
  reg        [0:0]    roundReg_11_1_4;
  reg        [0:0]    roundReg_11_1_5;
  reg        [0:0]    roundReg_11_1_6;
  reg        [0:0]    roundReg_11_1_7;
  reg        [0:0]    roundReg_12_0_0;
  reg        [0:0]    roundReg_12_0_1;
  reg        [0:0]    roundReg_12_0_2;
  reg        [0:0]    roundReg_12_0_3;
  reg        [0:0]    roundReg_12_0_4;
  reg        [0:0]    roundReg_12_0_5;
  reg        [0:0]    roundReg_12_0_6;
  reg        [0:0]    roundReg_12_0_7;
  reg        [0:0]    roundReg_12_1_0;
  reg        [0:0]    roundReg_12_1_1;
  reg        [0:0]    roundReg_12_1_2;
  reg        [0:0]    roundReg_12_1_3;
  reg        [0:0]    roundReg_12_1_4;
  reg        [0:0]    roundReg_12_1_5;
  reg        [0:0]    roundReg_12_1_6;
  reg        [0:0]    roundReg_12_1_7;
  reg        [0:0]    roundReg_13_0_0;
  reg        [0:0]    roundReg_13_0_1;
  reg        [0:0]    roundReg_13_0_2;
  reg        [0:0]    roundReg_13_0_3;
  reg        [0:0]    roundReg_13_0_4;
  reg        [0:0]    roundReg_13_0_5;
  reg        [0:0]    roundReg_13_0_6;
  reg        [0:0]    roundReg_13_0_7;
  reg        [0:0]    roundReg_13_1_0;
  reg        [0:0]    roundReg_13_1_1;
  reg        [0:0]    roundReg_13_1_2;
  reg        [0:0]    roundReg_13_1_3;
  reg        [0:0]    roundReg_13_1_4;
  reg        [0:0]    roundReg_13_1_5;
  reg        [0:0]    roundReg_13_1_6;
  reg        [0:0]    roundReg_13_1_7;
  reg        [0:0]    roundReg_14_0_0;
  reg        [0:0]    roundReg_14_0_1;
  reg        [0:0]    roundReg_14_0_2;
  reg        [0:0]    roundReg_14_0_3;
  reg        [0:0]    roundReg_14_0_4;
  reg        [0:0]    roundReg_14_0_5;
  reg        [0:0]    roundReg_14_0_6;
  reg        [0:0]    roundReg_14_0_7;
  reg        [0:0]    roundReg_14_1_0;
  reg        [0:0]    roundReg_14_1_1;
  reg        [0:0]    roundReg_14_1_2;
  reg        [0:0]    roundReg_14_1_3;
  reg        [0:0]    roundReg_14_1_4;
  reg        [0:0]    roundReg_14_1_5;
  reg        [0:0]    roundReg_14_1_6;
  reg        [0:0]    roundReg_14_1_7;
  reg        [0:0]    roundReg_15_0_0;
  reg        [0:0]    roundReg_15_0_1;
  reg        [0:0]    roundReg_15_0_2;
  reg        [0:0]    roundReg_15_0_3;
  reg        [0:0]    roundReg_15_0_4;
  reg        [0:0]    roundReg_15_0_5;
  reg        [0:0]    roundReg_15_0_6;
  reg        [0:0]    roundReg_15_0_7;
  reg        [0:0]    roundReg_15_1_0;
  reg        [0:0]    roundReg_15_1_1;
  reg        [0:0]    roundReg_15_1_2;
  reg        [0:0]    roundReg_15_1_3;
  reg        [0:0]    roundReg_15_1_4;
  reg        [0:0]    roundReg_15_1_5;
  reg        [0:0]    roundReg_15_1_6;
  reg        [0:0]    roundReg_15_1_7;

  AES_KeyAddition keyAdd (
    .port_state_in_0_0_0   (port_state_in_0_0_0         ), //i
    .port_state_in_0_0_1   (port_state_in_0_0_1         ), //i
    .port_state_in_0_0_2   (port_state_in_0_0_2         ), //i
    .port_state_in_0_0_3   (port_state_in_0_0_3         ), //i
    .port_state_in_0_0_4   (port_state_in_0_0_4         ), //i
    .port_state_in_0_0_5   (port_state_in_0_0_5         ), //i
    .port_state_in_0_0_6   (port_state_in_0_0_6         ), //i
    .port_state_in_0_0_7   (port_state_in_0_0_7         ), //i
    .port_state_in_0_1_0   (port_state_in_0_1_0         ), //i
    .port_state_in_0_1_1   (port_state_in_0_1_1         ), //i
    .port_state_in_0_1_2   (port_state_in_0_1_2         ), //i
    .port_state_in_0_1_3   (port_state_in_0_1_3         ), //i
    .port_state_in_0_1_4   (port_state_in_0_1_4         ), //i
    .port_state_in_0_1_5   (port_state_in_0_1_5         ), //i
    .port_state_in_0_1_6   (port_state_in_0_1_6         ), //i
    .port_state_in_0_1_7   (port_state_in_0_1_7         ), //i
    .port_state_in_1_0_0   (port_state_in_1_0_0         ), //i
    .port_state_in_1_0_1   (port_state_in_1_0_1         ), //i
    .port_state_in_1_0_2   (port_state_in_1_0_2         ), //i
    .port_state_in_1_0_3   (port_state_in_1_0_3         ), //i
    .port_state_in_1_0_4   (port_state_in_1_0_4         ), //i
    .port_state_in_1_0_5   (port_state_in_1_0_5         ), //i
    .port_state_in_1_0_6   (port_state_in_1_0_6         ), //i
    .port_state_in_1_0_7   (port_state_in_1_0_7         ), //i
    .port_state_in_1_1_0   (port_state_in_1_1_0         ), //i
    .port_state_in_1_1_1   (port_state_in_1_1_1         ), //i
    .port_state_in_1_1_2   (port_state_in_1_1_2         ), //i
    .port_state_in_1_1_3   (port_state_in_1_1_3         ), //i
    .port_state_in_1_1_4   (port_state_in_1_1_4         ), //i
    .port_state_in_1_1_5   (port_state_in_1_1_5         ), //i
    .port_state_in_1_1_6   (port_state_in_1_1_6         ), //i
    .port_state_in_1_1_7   (port_state_in_1_1_7         ), //i
    .port_state_in_2_0_0   (port_state_in_2_0_0         ), //i
    .port_state_in_2_0_1   (port_state_in_2_0_1         ), //i
    .port_state_in_2_0_2   (port_state_in_2_0_2         ), //i
    .port_state_in_2_0_3   (port_state_in_2_0_3         ), //i
    .port_state_in_2_0_4   (port_state_in_2_0_4         ), //i
    .port_state_in_2_0_5   (port_state_in_2_0_5         ), //i
    .port_state_in_2_0_6   (port_state_in_2_0_6         ), //i
    .port_state_in_2_0_7   (port_state_in_2_0_7         ), //i
    .port_state_in_2_1_0   (port_state_in_2_1_0         ), //i
    .port_state_in_2_1_1   (port_state_in_2_1_1         ), //i
    .port_state_in_2_1_2   (port_state_in_2_1_2         ), //i
    .port_state_in_2_1_3   (port_state_in_2_1_3         ), //i
    .port_state_in_2_1_4   (port_state_in_2_1_4         ), //i
    .port_state_in_2_1_5   (port_state_in_2_1_5         ), //i
    .port_state_in_2_1_6   (port_state_in_2_1_6         ), //i
    .port_state_in_2_1_7   (port_state_in_2_1_7         ), //i
    .port_state_in_3_0_0   (port_state_in_3_0_0         ), //i
    .port_state_in_3_0_1   (port_state_in_3_0_1         ), //i
    .port_state_in_3_0_2   (port_state_in_3_0_2         ), //i
    .port_state_in_3_0_3   (port_state_in_3_0_3         ), //i
    .port_state_in_3_0_4   (port_state_in_3_0_4         ), //i
    .port_state_in_3_0_5   (port_state_in_3_0_5         ), //i
    .port_state_in_3_0_6   (port_state_in_3_0_6         ), //i
    .port_state_in_3_0_7   (port_state_in_3_0_7         ), //i
    .port_state_in_3_1_0   (port_state_in_3_1_0         ), //i
    .port_state_in_3_1_1   (port_state_in_3_1_1         ), //i
    .port_state_in_3_1_2   (port_state_in_3_1_2         ), //i
    .port_state_in_3_1_3   (port_state_in_3_1_3         ), //i
    .port_state_in_3_1_4   (port_state_in_3_1_4         ), //i
    .port_state_in_3_1_5   (port_state_in_3_1_5         ), //i
    .port_state_in_3_1_6   (port_state_in_3_1_6         ), //i
    .port_state_in_3_1_7   (port_state_in_3_1_7         ), //i
    .port_state_in_4_0_0   (port_state_in_4_0_0         ), //i
    .port_state_in_4_0_1   (port_state_in_4_0_1         ), //i
    .port_state_in_4_0_2   (port_state_in_4_0_2         ), //i
    .port_state_in_4_0_3   (port_state_in_4_0_3         ), //i
    .port_state_in_4_0_4   (port_state_in_4_0_4         ), //i
    .port_state_in_4_0_5   (port_state_in_4_0_5         ), //i
    .port_state_in_4_0_6   (port_state_in_4_0_6         ), //i
    .port_state_in_4_0_7   (port_state_in_4_0_7         ), //i
    .port_state_in_4_1_0   (port_state_in_4_1_0         ), //i
    .port_state_in_4_1_1   (port_state_in_4_1_1         ), //i
    .port_state_in_4_1_2   (port_state_in_4_1_2         ), //i
    .port_state_in_4_1_3   (port_state_in_4_1_3         ), //i
    .port_state_in_4_1_4   (port_state_in_4_1_4         ), //i
    .port_state_in_4_1_5   (port_state_in_4_1_5         ), //i
    .port_state_in_4_1_6   (port_state_in_4_1_6         ), //i
    .port_state_in_4_1_7   (port_state_in_4_1_7         ), //i
    .port_state_in_5_0_0   (port_state_in_5_0_0         ), //i
    .port_state_in_5_0_1   (port_state_in_5_0_1         ), //i
    .port_state_in_5_0_2   (port_state_in_5_0_2         ), //i
    .port_state_in_5_0_3   (port_state_in_5_0_3         ), //i
    .port_state_in_5_0_4   (port_state_in_5_0_4         ), //i
    .port_state_in_5_0_5   (port_state_in_5_0_5         ), //i
    .port_state_in_5_0_6   (port_state_in_5_0_6         ), //i
    .port_state_in_5_0_7   (port_state_in_5_0_7         ), //i
    .port_state_in_5_1_0   (port_state_in_5_1_0         ), //i
    .port_state_in_5_1_1   (port_state_in_5_1_1         ), //i
    .port_state_in_5_1_2   (port_state_in_5_1_2         ), //i
    .port_state_in_5_1_3   (port_state_in_5_1_3         ), //i
    .port_state_in_5_1_4   (port_state_in_5_1_4         ), //i
    .port_state_in_5_1_5   (port_state_in_5_1_5         ), //i
    .port_state_in_5_1_6   (port_state_in_5_1_6         ), //i
    .port_state_in_5_1_7   (port_state_in_5_1_7         ), //i
    .port_state_in_6_0_0   (port_state_in_6_0_0         ), //i
    .port_state_in_6_0_1   (port_state_in_6_0_1         ), //i
    .port_state_in_6_0_2   (port_state_in_6_0_2         ), //i
    .port_state_in_6_0_3   (port_state_in_6_0_3         ), //i
    .port_state_in_6_0_4   (port_state_in_6_0_4         ), //i
    .port_state_in_6_0_5   (port_state_in_6_0_5         ), //i
    .port_state_in_6_0_6   (port_state_in_6_0_6         ), //i
    .port_state_in_6_0_7   (port_state_in_6_0_7         ), //i
    .port_state_in_6_1_0   (port_state_in_6_1_0         ), //i
    .port_state_in_6_1_1   (port_state_in_6_1_1         ), //i
    .port_state_in_6_1_2   (port_state_in_6_1_2         ), //i
    .port_state_in_6_1_3   (port_state_in_6_1_3         ), //i
    .port_state_in_6_1_4   (port_state_in_6_1_4         ), //i
    .port_state_in_6_1_5   (port_state_in_6_1_5         ), //i
    .port_state_in_6_1_6   (port_state_in_6_1_6         ), //i
    .port_state_in_6_1_7   (port_state_in_6_1_7         ), //i
    .port_state_in_7_0_0   (port_state_in_7_0_0         ), //i
    .port_state_in_7_0_1   (port_state_in_7_0_1         ), //i
    .port_state_in_7_0_2   (port_state_in_7_0_2         ), //i
    .port_state_in_7_0_3   (port_state_in_7_0_3         ), //i
    .port_state_in_7_0_4   (port_state_in_7_0_4         ), //i
    .port_state_in_7_0_5   (port_state_in_7_0_5         ), //i
    .port_state_in_7_0_6   (port_state_in_7_0_6         ), //i
    .port_state_in_7_0_7   (port_state_in_7_0_7         ), //i
    .port_state_in_7_1_0   (port_state_in_7_1_0         ), //i
    .port_state_in_7_1_1   (port_state_in_7_1_1         ), //i
    .port_state_in_7_1_2   (port_state_in_7_1_2         ), //i
    .port_state_in_7_1_3   (port_state_in_7_1_3         ), //i
    .port_state_in_7_1_4   (port_state_in_7_1_4         ), //i
    .port_state_in_7_1_5   (port_state_in_7_1_5         ), //i
    .port_state_in_7_1_6   (port_state_in_7_1_6         ), //i
    .port_state_in_7_1_7   (port_state_in_7_1_7         ), //i
    .port_state_in_8_0_0   (port_state_in_8_0_0         ), //i
    .port_state_in_8_0_1   (port_state_in_8_0_1         ), //i
    .port_state_in_8_0_2   (port_state_in_8_0_2         ), //i
    .port_state_in_8_0_3   (port_state_in_8_0_3         ), //i
    .port_state_in_8_0_4   (port_state_in_8_0_4         ), //i
    .port_state_in_8_0_5   (port_state_in_8_0_5         ), //i
    .port_state_in_8_0_6   (port_state_in_8_0_6         ), //i
    .port_state_in_8_0_7   (port_state_in_8_0_7         ), //i
    .port_state_in_8_1_0   (port_state_in_8_1_0         ), //i
    .port_state_in_8_1_1   (port_state_in_8_1_1         ), //i
    .port_state_in_8_1_2   (port_state_in_8_1_2         ), //i
    .port_state_in_8_1_3   (port_state_in_8_1_3         ), //i
    .port_state_in_8_1_4   (port_state_in_8_1_4         ), //i
    .port_state_in_8_1_5   (port_state_in_8_1_5         ), //i
    .port_state_in_8_1_6   (port_state_in_8_1_6         ), //i
    .port_state_in_8_1_7   (port_state_in_8_1_7         ), //i
    .port_state_in_9_0_0   (port_state_in_9_0_0         ), //i
    .port_state_in_9_0_1   (port_state_in_9_0_1         ), //i
    .port_state_in_9_0_2   (port_state_in_9_0_2         ), //i
    .port_state_in_9_0_3   (port_state_in_9_0_3         ), //i
    .port_state_in_9_0_4   (port_state_in_9_0_4         ), //i
    .port_state_in_9_0_5   (port_state_in_9_0_5         ), //i
    .port_state_in_9_0_6   (port_state_in_9_0_6         ), //i
    .port_state_in_9_0_7   (port_state_in_9_0_7         ), //i
    .port_state_in_9_1_0   (port_state_in_9_1_0         ), //i
    .port_state_in_9_1_1   (port_state_in_9_1_1         ), //i
    .port_state_in_9_1_2   (port_state_in_9_1_2         ), //i
    .port_state_in_9_1_3   (port_state_in_9_1_3         ), //i
    .port_state_in_9_1_4   (port_state_in_9_1_4         ), //i
    .port_state_in_9_1_5   (port_state_in_9_1_5         ), //i
    .port_state_in_9_1_6   (port_state_in_9_1_6         ), //i
    .port_state_in_9_1_7   (port_state_in_9_1_7         ), //i
    .port_state_in_10_0_0  (port_state_in_10_0_0        ), //i
    .port_state_in_10_0_1  (port_state_in_10_0_1        ), //i
    .port_state_in_10_0_2  (port_state_in_10_0_2        ), //i
    .port_state_in_10_0_3  (port_state_in_10_0_3        ), //i
    .port_state_in_10_0_4  (port_state_in_10_0_4        ), //i
    .port_state_in_10_0_5  (port_state_in_10_0_5        ), //i
    .port_state_in_10_0_6  (port_state_in_10_0_6        ), //i
    .port_state_in_10_0_7  (port_state_in_10_0_7        ), //i
    .port_state_in_10_1_0  (port_state_in_10_1_0        ), //i
    .port_state_in_10_1_1  (port_state_in_10_1_1        ), //i
    .port_state_in_10_1_2  (port_state_in_10_1_2        ), //i
    .port_state_in_10_1_3  (port_state_in_10_1_3        ), //i
    .port_state_in_10_1_4  (port_state_in_10_1_4        ), //i
    .port_state_in_10_1_5  (port_state_in_10_1_5        ), //i
    .port_state_in_10_1_6  (port_state_in_10_1_6        ), //i
    .port_state_in_10_1_7  (port_state_in_10_1_7        ), //i
    .port_state_in_11_0_0  (port_state_in_11_0_0        ), //i
    .port_state_in_11_0_1  (port_state_in_11_0_1        ), //i
    .port_state_in_11_0_2  (port_state_in_11_0_2        ), //i
    .port_state_in_11_0_3  (port_state_in_11_0_3        ), //i
    .port_state_in_11_0_4  (port_state_in_11_0_4        ), //i
    .port_state_in_11_0_5  (port_state_in_11_0_5        ), //i
    .port_state_in_11_0_6  (port_state_in_11_0_6        ), //i
    .port_state_in_11_0_7  (port_state_in_11_0_7        ), //i
    .port_state_in_11_1_0  (port_state_in_11_1_0        ), //i
    .port_state_in_11_1_1  (port_state_in_11_1_1        ), //i
    .port_state_in_11_1_2  (port_state_in_11_1_2        ), //i
    .port_state_in_11_1_3  (port_state_in_11_1_3        ), //i
    .port_state_in_11_1_4  (port_state_in_11_1_4        ), //i
    .port_state_in_11_1_5  (port_state_in_11_1_5        ), //i
    .port_state_in_11_1_6  (port_state_in_11_1_6        ), //i
    .port_state_in_11_1_7  (port_state_in_11_1_7        ), //i
    .port_state_in_12_0_0  (port_state_in_12_0_0        ), //i
    .port_state_in_12_0_1  (port_state_in_12_0_1        ), //i
    .port_state_in_12_0_2  (port_state_in_12_0_2        ), //i
    .port_state_in_12_0_3  (port_state_in_12_0_3        ), //i
    .port_state_in_12_0_4  (port_state_in_12_0_4        ), //i
    .port_state_in_12_0_5  (port_state_in_12_0_5        ), //i
    .port_state_in_12_0_6  (port_state_in_12_0_6        ), //i
    .port_state_in_12_0_7  (port_state_in_12_0_7        ), //i
    .port_state_in_12_1_0  (port_state_in_12_1_0        ), //i
    .port_state_in_12_1_1  (port_state_in_12_1_1        ), //i
    .port_state_in_12_1_2  (port_state_in_12_1_2        ), //i
    .port_state_in_12_1_3  (port_state_in_12_1_3        ), //i
    .port_state_in_12_1_4  (port_state_in_12_1_4        ), //i
    .port_state_in_12_1_5  (port_state_in_12_1_5        ), //i
    .port_state_in_12_1_6  (port_state_in_12_1_6        ), //i
    .port_state_in_12_1_7  (port_state_in_12_1_7        ), //i
    .port_state_in_13_0_0  (port_state_in_13_0_0        ), //i
    .port_state_in_13_0_1  (port_state_in_13_0_1        ), //i
    .port_state_in_13_0_2  (port_state_in_13_0_2        ), //i
    .port_state_in_13_0_3  (port_state_in_13_0_3        ), //i
    .port_state_in_13_0_4  (port_state_in_13_0_4        ), //i
    .port_state_in_13_0_5  (port_state_in_13_0_5        ), //i
    .port_state_in_13_0_6  (port_state_in_13_0_6        ), //i
    .port_state_in_13_0_7  (port_state_in_13_0_7        ), //i
    .port_state_in_13_1_0  (port_state_in_13_1_0        ), //i
    .port_state_in_13_1_1  (port_state_in_13_1_1        ), //i
    .port_state_in_13_1_2  (port_state_in_13_1_2        ), //i
    .port_state_in_13_1_3  (port_state_in_13_1_3        ), //i
    .port_state_in_13_1_4  (port_state_in_13_1_4        ), //i
    .port_state_in_13_1_5  (port_state_in_13_1_5        ), //i
    .port_state_in_13_1_6  (port_state_in_13_1_6        ), //i
    .port_state_in_13_1_7  (port_state_in_13_1_7        ), //i
    .port_state_in_14_0_0  (port_state_in_14_0_0        ), //i
    .port_state_in_14_0_1  (port_state_in_14_0_1        ), //i
    .port_state_in_14_0_2  (port_state_in_14_0_2        ), //i
    .port_state_in_14_0_3  (port_state_in_14_0_3        ), //i
    .port_state_in_14_0_4  (port_state_in_14_0_4        ), //i
    .port_state_in_14_0_5  (port_state_in_14_0_5        ), //i
    .port_state_in_14_0_6  (port_state_in_14_0_6        ), //i
    .port_state_in_14_0_7  (port_state_in_14_0_7        ), //i
    .port_state_in_14_1_0  (port_state_in_14_1_0        ), //i
    .port_state_in_14_1_1  (port_state_in_14_1_1        ), //i
    .port_state_in_14_1_2  (port_state_in_14_1_2        ), //i
    .port_state_in_14_1_3  (port_state_in_14_1_3        ), //i
    .port_state_in_14_1_4  (port_state_in_14_1_4        ), //i
    .port_state_in_14_1_5  (port_state_in_14_1_5        ), //i
    .port_state_in_14_1_6  (port_state_in_14_1_6        ), //i
    .port_state_in_14_1_7  (port_state_in_14_1_7        ), //i
    .port_state_in_15_0_0  (port_state_in_15_0_0        ), //i
    .port_state_in_15_0_1  (port_state_in_15_0_1        ), //i
    .port_state_in_15_0_2  (port_state_in_15_0_2        ), //i
    .port_state_in_15_0_3  (port_state_in_15_0_3        ), //i
    .port_state_in_15_0_4  (port_state_in_15_0_4        ), //i
    .port_state_in_15_0_5  (port_state_in_15_0_5        ), //i
    .port_state_in_15_0_6  (port_state_in_15_0_6        ), //i
    .port_state_in_15_0_7  (port_state_in_15_0_7        ), //i
    .port_state_in_15_1_0  (port_state_in_15_1_0        ), //i
    .port_state_in_15_1_1  (port_state_in_15_1_1        ), //i
    .port_state_in_15_1_2  (port_state_in_15_1_2        ), //i
    .port_state_in_15_1_3  (port_state_in_15_1_3        ), //i
    .port_state_in_15_1_4  (port_state_in_15_1_4        ), //i
    .port_state_in_15_1_5  (port_state_in_15_1_5        ), //i
    .port_state_in_15_1_6  (port_state_in_15_1_6        ), //i
    .port_state_in_15_1_7  (port_state_in_15_1_7        ), //i
    .port_key_0_0_0        (port_key_0_0_0              ), //i
    .port_key_0_0_1        (port_key_0_0_1              ), //i
    .port_key_0_0_2        (port_key_0_0_2              ), //i
    .port_key_0_0_3        (port_key_0_0_3              ), //i
    .port_key_0_0_4        (port_key_0_0_4              ), //i
    .port_key_0_0_5        (port_key_0_0_5              ), //i
    .port_key_0_0_6        (port_key_0_0_6              ), //i
    .port_key_0_0_7        (port_key_0_0_7              ), //i
    .port_key_0_1_0        (port_key_0_1_0              ), //i
    .port_key_0_1_1        (port_key_0_1_1              ), //i
    .port_key_0_1_2        (port_key_0_1_2              ), //i
    .port_key_0_1_3        (port_key_0_1_3              ), //i
    .port_key_0_1_4        (port_key_0_1_4              ), //i
    .port_key_0_1_5        (port_key_0_1_5              ), //i
    .port_key_0_1_6        (port_key_0_1_6              ), //i
    .port_key_0_1_7        (port_key_0_1_7              ), //i
    .port_key_1_0_0        (port_key_1_0_0              ), //i
    .port_key_1_0_1        (port_key_1_0_1              ), //i
    .port_key_1_0_2        (port_key_1_0_2              ), //i
    .port_key_1_0_3        (port_key_1_0_3              ), //i
    .port_key_1_0_4        (port_key_1_0_4              ), //i
    .port_key_1_0_5        (port_key_1_0_5              ), //i
    .port_key_1_0_6        (port_key_1_0_6              ), //i
    .port_key_1_0_7        (port_key_1_0_7              ), //i
    .port_key_1_1_0        (port_key_1_1_0              ), //i
    .port_key_1_1_1        (port_key_1_1_1              ), //i
    .port_key_1_1_2        (port_key_1_1_2              ), //i
    .port_key_1_1_3        (port_key_1_1_3              ), //i
    .port_key_1_1_4        (port_key_1_1_4              ), //i
    .port_key_1_1_5        (port_key_1_1_5              ), //i
    .port_key_1_1_6        (port_key_1_1_6              ), //i
    .port_key_1_1_7        (port_key_1_1_7              ), //i
    .port_key_2_0_0        (port_key_2_0_0              ), //i
    .port_key_2_0_1        (port_key_2_0_1              ), //i
    .port_key_2_0_2        (port_key_2_0_2              ), //i
    .port_key_2_0_3        (port_key_2_0_3              ), //i
    .port_key_2_0_4        (port_key_2_0_4              ), //i
    .port_key_2_0_5        (port_key_2_0_5              ), //i
    .port_key_2_0_6        (port_key_2_0_6              ), //i
    .port_key_2_0_7        (port_key_2_0_7              ), //i
    .port_key_2_1_0        (port_key_2_1_0              ), //i
    .port_key_2_1_1        (port_key_2_1_1              ), //i
    .port_key_2_1_2        (port_key_2_1_2              ), //i
    .port_key_2_1_3        (port_key_2_1_3              ), //i
    .port_key_2_1_4        (port_key_2_1_4              ), //i
    .port_key_2_1_5        (port_key_2_1_5              ), //i
    .port_key_2_1_6        (port_key_2_1_6              ), //i
    .port_key_2_1_7        (port_key_2_1_7              ), //i
    .port_key_3_0_0        (port_key_3_0_0              ), //i
    .port_key_3_0_1        (port_key_3_0_1              ), //i
    .port_key_3_0_2        (port_key_3_0_2              ), //i
    .port_key_3_0_3        (port_key_3_0_3              ), //i
    .port_key_3_0_4        (port_key_3_0_4              ), //i
    .port_key_3_0_5        (port_key_3_0_5              ), //i
    .port_key_3_0_6        (port_key_3_0_6              ), //i
    .port_key_3_0_7        (port_key_3_0_7              ), //i
    .port_key_3_1_0        (port_key_3_1_0              ), //i
    .port_key_3_1_1        (port_key_3_1_1              ), //i
    .port_key_3_1_2        (port_key_3_1_2              ), //i
    .port_key_3_1_3        (port_key_3_1_3              ), //i
    .port_key_3_1_4        (port_key_3_1_4              ), //i
    .port_key_3_1_5        (port_key_3_1_5              ), //i
    .port_key_3_1_6        (port_key_3_1_6              ), //i
    .port_key_3_1_7        (port_key_3_1_7              ), //i
    .port_key_4_0_0        (port_key_4_0_0              ), //i
    .port_key_4_0_1        (port_key_4_0_1              ), //i
    .port_key_4_0_2        (port_key_4_0_2              ), //i
    .port_key_4_0_3        (port_key_4_0_3              ), //i
    .port_key_4_0_4        (port_key_4_0_4              ), //i
    .port_key_4_0_5        (port_key_4_0_5              ), //i
    .port_key_4_0_6        (port_key_4_0_6              ), //i
    .port_key_4_0_7        (port_key_4_0_7              ), //i
    .port_key_4_1_0        (port_key_4_1_0              ), //i
    .port_key_4_1_1        (port_key_4_1_1              ), //i
    .port_key_4_1_2        (port_key_4_1_2              ), //i
    .port_key_4_1_3        (port_key_4_1_3              ), //i
    .port_key_4_1_4        (port_key_4_1_4              ), //i
    .port_key_4_1_5        (port_key_4_1_5              ), //i
    .port_key_4_1_6        (port_key_4_1_6              ), //i
    .port_key_4_1_7        (port_key_4_1_7              ), //i
    .port_key_5_0_0        (port_key_5_0_0              ), //i
    .port_key_5_0_1        (port_key_5_0_1              ), //i
    .port_key_5_0_2        (port_key_5_0_2              ), //i
    .port_key_5_0_3        (port_key_5_0_3              ), //i
    .port_key_5_0_4        (port_key_5_0_4              ), //i
    .port_key_5_0_5        (port_key_5_0_5              ), //i
    .port_key_5_0_6        (port_key_5_0_6              ), //i
    .port_key_5_0_7        (port_key_5_0_7              ), //i
    .port_key_5_1_0        (port_key_5_1_0              ), //i
    .port_key_5_1_1        (port_key_5_1_1              ), //i
    .port_key_5_1_2        (port_key_5_1_2              ), //i
    .port_key_5_1_3        (port_key_5_1_3              ), //i
    .port_key_5_1_4        (port_key_5_1_4              ), //i
    .port_key_5_1_5        (port_key_5_1_5              ), //i
    .port_key_5_1_6        (port_key_5_1_6              ), //i
    .port_key_5_1_7        (port_key_5_1_7              ), //i
    .port_key_6_0_0        (port_key_6_0_0              ), //i
    .port_key_6_0_1        (port_key_6_0_1              ), //i
    .port_key_6_0_2        (port_key_6_0_2              ), //i
    .port_key_6_0_3        (port_key_6_0_3              ), //i
    .port_key_6_0_4        (port_key_6_0_4              ), //i
    .port_key_6_0_5        (port_key_6_0_5              ), //i
    .port_key_6_0_6        (port_key_6_0_6              ), //i
    .port_key_6_0_7        (port_key_6_0_7              ), //i
    .port_key_6_1_0        (port_key_6_1_0              ), //i
    .port_key_6_1_1        (port_key_6_1_1              ), //i
    .port_key_6_1_2        (port_key_6_1_2              ), //i
    .port_key_6_1_3        (port_key_6_1_3              ), //i
    .port_key_6_1_4        (port_key_6_1_4              ), //i
    .port_key_6_1_5        (port_key_6_1_5              ), //i
    .port_key_6_1_6        (port_key_6_1_6              ), //i
    .port_key_6_1_7        (port_key_6_1_7              ), //i
    .port_key_7_0_0        (port_key_7_0_0              ), //i
    .port_key_7_0_1        (port_key_7_0_1              ), //i
    .port_key_7_0_2        (port_key_7_0_2              ), //i
    .port_key_7_0_3        (port_key_7_0_3              ), //i
    .port_key_7_0_4        (port_key_7_0_4              ), //i
    .port_key_7_0_5        (port_key_7_0_5              ), //i
    .port_key_7_0_6        (port_key_7_0_6              ), //i
    .port_key_7_0_7        (port_key_7_0_7              ), //i
    .port_key_7_1_0        (port_key_7_1_0              ), //i
    .port_key_7_1_1        (port_key_7_1_1              ), //i
    .port_key_7_1_2        (port_key_7_1_2              ), //i
    .port_key_7_1_3        (port_key_7_1_3              ), //i
    .port_key_7_1_4        (port_key_7_1_4              ), //i
    .port_key_7_1_5        (port_key_7_1_5              ), //i
    .port_key_7_1_6        (port_key_7_1_6              ), //i
    .port_key_7_1_7        (port_key_7_1_7              ), //i
    .port_key_8_0_0        (port_key_8_0_0              ), //i
    .port_key_8_0_1        (port_key_8_0_1              ), //i
    .port_key_8_0_2        (port_key_8_0_2              ), //i
    .port_key_8_0_3        (port_key_8_0_3              ), //i
    .port_key_8_0_4        (port_key_8_0_4              ), //i
    .port_key_8_0_5        (port_key_8_0_5              ), //i
    .port_key_8_0_6        (port_key_8_0_6              ), //i
    .port_key_8_0_7        (port_key_8_0_7              ), //i
    .port_key_8_1_0        (port_key_8_1_0              ), //i
    .port_key_8_1_1        (port_key_8_1_1              ), //i
    .port_key_8_1_2        (port_key_8_1_2              ), //i
    .port_key_8_1_3        (port_key_8_1_3              ), //i
    .port_key_8_1_4        (port_key_8_1_4              ), //i
    .port_key_8_1_5        (port_key_8_1_5              ), //i
    .port_key_8_1_6        (port_key_8_1_6              ), //i
    .port_key_8_1_7        (port_key_8_1_7              ), //i
    .port_key_9_0_0        (port_key_9_0_0              ), //i
    .port_key_9_0_1        (port_key_9_0_1              ), //i
    .port_key_9_0_2        (port_key_9_0_2              ), //i
    .port_key_9_0_3        (port_key_9_0_3              ), //i
    .port_key_9_0_4        (port_key_9_0_4              ), //i
    .port_key_9_0_5        (port_key_9_0_5              ), //i
    .port_key_9_0_6        (port_key_9_0_6              ), //i
    .port_key_9_0_7        (port_key_9_0_7              ), //i
    .port_key_9_1_0        (port_key_9_1_0              ), //i
    .port_key_9_1_1        (port_key_9_1_1              ), //i
    .port_key_9_1_2        (port_key_9_1_2              ), //i
    .port_key_9_1_3        (port_key_9_1_3              ), //i
    .port_key_9_1_4        (port_key_9_1_4              ), //i
    .port_key_9_1_5        (port_key_9_1_5              ), //i
    .port_key_9_1_6        (port_key_9_1_6              ), //i
    .port_key_9_1_7        (port_key_9_1_7              ), //i
    .port_key_10_0_0       (port_key_10_0_0             ), //i
    .port_key_10_0_1       (port_key_10_0_1             ), //i
    .port_key_10_0_2       (port_key_10_0_2             ), //i
    .port_key_10_0_3       (port_key_10_0_3             ), //i
    .port_key_10_0_4       (port_key_10_0_4             ), //i
    .port_key_10_0_5       (port_key_10_0_5             ), //i
    .port_key_10_0_6       (port_key_10_0_6             ), //i
    .port_key_10_0_7       (port_key_10_0_7             ), //i
    .port_key_10_1_0       (port_key_10_1_0             ), //i
    .port_key_10_1_1       (port_key_10_1_1             ), //i
    .port_key_10_1_2       (port_key_10_1_2             ), //i
    .port_key_10_1_3       (port_key_10_1_3             ), //i
    .port_key_10_1_4       (port_key_10_1_4             ), //i
    .port_key_10_1_5       (port_key_10_1_5             ), //i
    .port_key_10_1_6       (port_key_10_1_6             ), //i
    .port_key_10_1_7       (port_key_10_1_7             ), //i
    .port_key_11_0_0       (port_key_11_0_0             ), //i
    .port_key_11_0_1       (port_key_11_0_1             ), //i
    .port_key_11_0_2       (port_key_11_0_2             ), //i
    .port_key_11_0_3       (port_key_11_0_3             ), //i
    .port_key_11_0_4       (port_key_11_0_4             ), //i
    .port_key_11_0_5       (port_key_11_0_5             ), //i
    .port_key_11_0_6       (port_key_11_0_6             ), //i
    .port_key_11_0_7       (port_key_11_0_7             ), //i
    .port_key_11_1_0       (port_key_11_1_0             ), //i
    .port_key_11_1_1       (port_key_11_1_1             ), //i
    .port_key_11_1_2       (port_key_11_1_2             ), //i
    .port_key_11_1_3       (port_key_11_1_3             ), //i
    .port_key_11_1_4       (port_key_11_1_4             ), //i
    .port_key_11_1_5       (port_key_11_1_5             ), //i
    .port_key_11_1_6       (port_key_11_1_6             ), //i
    .port_key_11_1_7       (port_key_11_1_7             ), //i
    .port_key_12_0_0       (port_key_12_0_0             ), //i
    .port_key_12_0_1       (port_key_12_0_1             ), //i
    .port_key_12_0_2       (port_key_12_0_2             ), //i
    .port_key_12_0_3       (port_key_12_0_3             ), //i
    .port_key_12_0_4       (port_key_12_0_4             ), //i
    .port_key_12_0_5       (port_key_12_0_5             ), //i
    .port_key_12_0_6       (port_key_12_0_6             ), //i
    .port_key_12_0_7       (port_key_12_0_7             ), //i
    .port_key_12_1_0       (port_key_12_1_0             ), //i
    .port_key_12_1_1       (port_key_12_1_1             ), //i
    .port_key_12_1_2       (port_key_12_1_2             ), //i
    .port_key_12_1_3       (port_key_12_1_3             ), //i
    .port_key_12_1_4       (port_key_12_1_4             ), //i
    .port_key_12_1_5       (port_key_12_1_5             ), //i
    .port_key_12_1_6       (port_key_12_1_6             ), //i
    .port_key_12_1_7       (port_key_12_1_7             ), //i
    .port_key_13_0_0       (port_key_13_0_0             ), //i
    .port_key_13_0_1       (port_key_13_0_1             ), //i
    .port_key_13_0_2       (port_key_13_0_2             ), //i
    .port_key_13_0_3       (port_key_13_0_3             ), //i
    .port_key_13_0_4       (port_key_13_0_4             ), //i
    .port_key_13_0_5       (port_key_13_0_5             ), //i
    .port_key_13_0_6       (port_key_13_0_6             ), //i
    .port_key_13_0_7       (port_key_13_0_7             ), //i
    .port_key_13_1_0       (port_key_13_1_0             ), //i
    .port_key_13_1_1       (port_key_13_1_1             ), //i
    .port_key_13_1_2       (port_key_13_1_2             ), //i
    .port_key_13_1_3       (port_key_13_1_3             ), //i
    .port_key_13_1_4       (port_key_13_1_4             ), //i
    .port_key_13_1_5       (port_key_13_1_5             ), //i
    .port_key_13_1_6       (port_key_13_1_6             ), //i
    .port_key_13_1_7       (port_key_13_1_7             ), //i
    .port_key_14_0_0       (port_key_14_0_0             ), //i
    .port_key_14_0_1       (port_key_14_0_1             ), //i
    .port_key_14_0_2       (port_key_14_0_2             ), //i
    .port_key_14_0_3       (port_key_14_0_3             ), //i
    .port_key_14_0_4       (port_key_14_0_4             ), //i
    .port_key_14_0_5       (port_key_14_0_5             ), //i
    .port_key_14_0_6       (port_key_14_0_6             ), //i
    .port_key_14_0_7       (port_key_14_0_7             ), //i
    .port_key_14_1_0       (port_key_14_1_0             ), //i
    .port_key_14_1_1       (port_key_14_1_1             ), //i
    .port_key_14_1_2       (port_key_14_1_2             ), //i
    .port_key_14_1_3       (port_key_14_1_3             ), //i
    .port_key_14_1_4       (port_key_14_1_4             ), //i
    .port_key_14_1_5       (port_key_14_1_5             ), //i
    .port_key_14_1_6       (port_key_14_1_6             ), //i
    .port_key_14_1_7       (port_key_14_1_7             ), //i
    .port_key_15_0_0       (port_key_15_0_0             ), //i
    .port_key_15_0_1       (port_key_15_0_1             ), //i
    .port_key_15_0_2       (port_key_15_0_2             ), //i
    .port_key_15_0_3       (port_key_15_0_3             ), //i
    .port_key_15_0_4       (port_key_15_0_4             ), //i
    .port_key_15_0_5       (port_key_15_0_5             ), //i
    .port_key_15_0_6       (port_key_15_0_6             ), //i
    .port_key_15_0_7       (port_key_15_0_7             ), //i
    .port_key_15_1_0       (port_key_15_1_0             ), //i
    .port_key_15_1_1       (port_key_15_1_1             ), //i
    .port_key_15_1_2       (port_key_15_1_2             ), //i
    .port_key_15_1_3       (port_key_15_1_3             ), //i
    .port_key_15_1_4       (port_key_15_1_4             ), //i
    .port_key_15_1_5       (port_key_15_1_5             ), //i
    .port_key_15_1_6       (port_key_15_1_6             ), //i
    .port_key_15_1_7       (port_key_15_1_7             ), //i
    .port_state_out_0_0_0  (keyAdd_port_state_out_0_0_0 ), //o
    .port_state_out_0_0_1  (keyAdd_port_state_out_0_0_1 ), //o
    .port_state_out_0_0_2  (keyAdd_port_state_out_0_0_2 ), //o
    .port_state_out_0_0_3  (keyAdd_port_state_out_0_0_3 ), //o
    .port_state_out_0_0_4  (keyAdd_port_state_out_0_0_4 ), //o
    .port_state_out_0_0_5  (keyAdd_port_state_out_0_0_5 ), //o
    .port_state_out_0_0_6  (keyAdd_port_state_out_0_0_6 ), //o
    .port_state_out_0_0_7  (keyAdd_port_state_out_0_0_7 ), //o
    .port_state_out_0_1_0  (keyAdd_port_state_out_0_1_0 ), //o
    .port_state_out_0_1_1  (keyAdd_port_state_out_0_1_1 ), //o
    .port_state_out_0_1_2  (keyAdd_port_state_out_0_1_2 ), //o
    .port_state_out_0_1_3  (keyAdd_port_state_out_0_1_3 ), //o
    .port_state_out_0_1_4  (keyAdd_port_state_out_0_1_4 ), //o
    .port_state_out_0_1_5  (keyAdd_port_state_out_0_1_5 ), //o
    .port_state_out_0_1_6  (keyAdd_port_state_out_0_1_6 ), //o
    .port_state_out_0_1_7  (keyAdd_port_state_out_0_1_7 ), //o
    .port_state_out_1_0_0  (keyAdd_port_state_out_1_0_0 ), //o
    .port_state_out_1_0_1  (keyAdd_port_state_out_1_0_1 ), //o
    .port_state_out_1_0_2  (keyAdd_port_state_out_1_0_2 ), //o
    .port_state_out_1_0_3  (keyAdd_port_state_out_1_0_3 ), //o
    .port_state_out_1_0_4  (keyAdd_port_state_out_1_0_4 ), //o
    .port_state_out_1_0_5  (keyAdd_port_state_out_1_0_5 ), //o
    .port_state_out_1_0_6  (keyAdd_port_state_out_1_0_6 ), //o
    .port_state_out_1_0_7  (keyAdd_port_state_out_1_0_7 ), //o
    .port_state_out_1_1_0  (keyAdd_port_state_out_1_1_0 ), //o
    .port_state_out_1_1_1  (keyAdd_port_state_out_1_1_1 ), //o
    .port_state_out_1_1_2  (keyAdd_port_state_out_1_1_2 ), //o
    .port_state_out_1_1_3  (keyAdd_port_state_out_1_1_3 ), //o
    .port_state_out_1_1_4  (keyAdd_port_state_out_1_1_4 ), //o
    .port_state_out_1_1_5  (keyAdd_port_state_out_1_1_5 ), //o
    .port_state_out_1_1_6  (keyAdd_port_state_out_1_1_6 ), //o
    .port_state_out_1_1_7  (keyAdd_port_state_out_1_1_7 ), //o
    .port_state_out_2_0_0  (keyAdd_port_state_out_2_0_0 ), //o
    .port_state_out_2_0_1  (keyAdd_port_state_out_2_0_1 ), //o
    .port_state_out_2_0_2  (keyAdd_port_state_out_2_0_2 ), //o
    .port_state_out_2_0_3  (keyAdd_port_state_out_2_0_3 ), //o
    .port_state_out_2_0_4  (keyAdd_port_state_out_2_0_4 ), //o
    .port_state_out_2_0_5  (keyAdd_port_state_out_2_0_5 ), //o
    .port_state_out_2_0_6  (keyAdd_port_state_out_2_0_6 ), //o
    .port_state_out_2_0_7  (keyAdd_port_state_out_2_0_7 ), //o
    .port_state_out_2_1_0  (keyAdd_port_state_out_2_1_0 ), //o
    .port_state_out_2_1_1  (keyAdd_port_state_out_2_1_1 ), //o
    .port_state_out_2_1_2  (keyAdd_port_state_out_2_1_2 ), //o
    .port_state_out_2_1_3  (keyAdd_port_state_out_2_1_3 ), //o
    .port_state_out_2_1_4  (keyAdd_port_state_out_2_1_4 ), //o
    .port_state_out_2_1_5  (keyAdd_port_state_out_2_1_5 ), //o
    .port_state_out_2_1_6  (keyAdd_port_state_out_2_1_6 ), //o
    .port_state_out_2_1_7  (keyAdd_port_state_out_2_1_7 ), //o
    .port_state_out_3_0_0  (keyAdd_port_state_out_3_0_0 ), //o
    .port_state_out_3_0_1  (keyAdd_port_state_out_3_0_1 ), //o
    .port_state_out_3_0_2  (keyAdd_port_state_out_3_0_2 ), //o
    .port_state_out_3_0_3  (keyAdd_port_state_out_3_0_3 ), //o
    .port_state_out_3_0_4  (keyAdd_port_state_out_3_0_4 ), //o
    .port_state_out_3_0_5  (keyAdd_port_state_out_3_0_5 ), //o
    .port_state_out_3_0_6  (keyAdd_port_state_out_3_0_6 ), //o
    .port_state_out_3_0_7  (keyAdd_port_state_out_3_0_7 ), //o
    .port_state_out_3_1_0  (keyAdd_port_state_out_3_1_0 ), //o
    .port_state_out_3_1_1  (keyAdd_port_state_out_3_1_1 ), //o
    .port_state_out_3_1_2  (keyAdd_port_state_out_3_1_2 ), //o
    .port_state_out_3_1_3  (keyAdd_port_state_out_3_1_3 ), //o
    .port_state_out_3_1_4  (keyAdd_port_state_out_3_1_4 ), //o
    .port_state_out_3_1_5  (keyAdd_port_state_out_3_1_5 ), //o
    .port_state_out_3_1_6  (keyAdd_port_state_out_3_1_6 ), //o
    .port_state_out_3_1_7  (keyAdd_port_state_out_3_1_7 ), //o
    .port_state_out_4_0_0  (keyAdd_port_state_out_4_0_0 ), //o
    .port_state_out_4_0_1  (keyAdd_port_state_out_4_0_1 ), //o
    .port_state_out_4_0_2  (keyAdd_port_state_out_4_0_2 ), //o
    .port_state_out_4_0_3  (keyAdd_port_state_out_4_0_3 ), //o
    .port_state_out_4_0_4  (keyAdd_port_state_out_4_0_4 ), //o
    .port_state_out_4_0_5  (keyAdd_port_state_out_4_0_5 ), //o
    .port_state_out_4_0_6  (keyAdd_port_state_out_4_0_6 ), //o
    .port_state_out_4_0_7  (keyAdd_port_state_out_4_0_7 ), //o
    .port_state_out_4_1_0  (keyAdd_port_state_out_4_1_0 ), //o
    .port_state_out_4_1_1  (keyAdd_port_state_out_4_1_1 ), //o
    .port_state_out_4_1_2  (keyAdd_port_state_out_4_1_2 ), //o
    .port_state_out_4_1_3  (keyAdd_port_state_out_4_1_3 ), //o
    .port_state_out_4_1_4  (keyAdd_port_state_out_4_1_4 ), //o
    .port_state_out_4_1_5  (keyAdd_port_state_out_4_1_5 ), //o
    .port_state_out_4_1_6  (keyAdd_port_state_out_4_1_6 ), //o
    .port_state_out_4_1_7  (keyAdd_port_state_out_4_1_7 ), //o
    .port_state_out_5_0_0  (keyAdd_port_state_out_5_0_0 ), //o
    .port_state_out_5_0_1  (keyAdd_port_state_out_5_0_1 ), //o
    .port_state_out_5_0_2  (keyAdd_port_state_out_5_0_2 ), //o
    .port_state_out_5_0_3  (keyAdd_port_state_out_5_0_3 ), //o
    .port_state_out_5_0_4  (keyAdd_port_state_out_5_0_4 ), //o
    .port_state_out_5_0_5  (keyAdd_port_state_out_5_0_5 ), //o
    .port_state_out_5_0_6  (keyAdd_port_state_out_5_0_6 ), //o
    .port_state_out_5_0_7  (keyAdd_port_state_out_5_0_7 ), //o
    .port_state_out_5_1_0  (keyAdd_port_state_out_5_1_0 ), //o
    .port_state_out_5_1_1  (keyAdd_port_state_out_5_1_1 ), //o
    .port_state_out_5_1_2  (keyAdd_port_state_out_5_1_2 ), //o
    .port_state_out_5_1_3  (keyAdd_port_state_out_5_1_3 ), //o
    .port_state_out_5_1_4  (keyAdd_port_state_out_5_1_4 ), //o
    .port_state_out_5_1_5  (keyAdd_port_state_out_5_1_5 ), //o
    .port_state_out_5_1_6  (keyAdd_port_state_out_5_1_6 ), //o
    .port_state_out_5_1_7  (keyAdd_port_state_out_5_1_7 ), //o
    .port_state_out_6_0_0  (keyAdd_port_state_out_6_0_0 ), //o
    .port_state_out_6_0_1  (keyAdd_port_state_out_6_0_1 ), //o
    .port_state_out_6_0_2  (keyAdd_port_state_out_6_0_2 ), //o
    .port_state_out_6_0_3  (keyAdd_port_state_out_6_0_3 ), //o
    .port_state_out_6_0_4  (keyAdd_port_state_out_6_0_4 ), //o
    .port_state_out_6_0_5  (keyAdd_port_state_out_6_0_5 ), //o
    .port_state_out_6_0_6  (keyAdd_port_state_out_6_0_6 ), //o
    .port_state_out_6_0_7  (keyAdd_port_state_out_6_0_7 ), //o
    .port_state_out_6_1_0  (keyAdd_port_state_out_6_1_0 ), //o
    .port_state_out_6_1_1  (keyAdd_port_state_out_6_1_1 ), //o
    .port_state_out_6_1_2  (keyAdd_port_state_out_6_1_2 ), //o
    .port_state_out_6_1_3  (keyAdd_port_state_out_6_1_3 ), //o
    .port_state_out_6_1_4  (keyAdd_port_state_out_6_1_4 ), //o
    .port_state_out_6_1_5  (keyAdd_port_state_out_6_1_5 ), //o
    .port_state_out_6_1_6  (keyAdd_port_state_out_6_1_6 ), //o
    .port_state_out_6_1_7  (keyAdd_port_state_out_6_1_7 ), //o
    .port_state_out_7_0_0  (keyAdd_port_state_out_7_0_0 ), //o
    .port_state_out_7_0_1  (keyAdd_port_state_out_7_0_1 ), //o
    .port_state_out_7_0_2  (keyAdd_port_state_out_7_0_2 ), //o
    .port_state_out_7_0_3  (keyAdd_port_state_out_7_0_3 ), //o
    .port_state_out_7_0_4  (keyAdd_port_state_out_7_0_4 ), //o
    .port_state_out_7_0_5  (keyAdd_port_state_out_7_0_5 ), //o
    .port_state_out_7_0_6  (keyAdd_port_state_out_7_0_6 ), //o
    .port_state_out_7_0_7  (keyAdd_port_state_out_7_0_7 ), //o
    .port_state_out_7_1_0  (keyAdd_port_state_out_7_1_0 ), //o
    .port_state_out_7_1_1  (keyAdd_port_state_out_7_1_1 ), //o
    .port_state_out_7_1_2  (keyAdd_port_state_out_7_1_2 ), //o
    .port_state_out_7_1_3  (keyAdd_port_state_out_7_1_3 ), //o
    .port_state_out_7_1_4  (keyAdd_port_state_out_7_1_4 ), //o
    .port_state_out_7_1_5  (keyAdd_port_state_out_7_1_5 ), //o
    .port_state_out_7_1_6  (keyAdd_port_state_out_7_1_6 ), //o
    .port_state_out_7_1_7  (keyAdd_port_state_out_7_1_7 ), //o
    .port_state_out_8_0_0  (keyAdd_port_state_out_8_0_0 ), //o
    .port_state_out_8_0_1  (keyAdd_port_state_out_8_0_1 ), //o
    .port_state_out_8_0_2  (keyAdd_port_state_out_8_0_2 ), //o
    .port_state_out_8_0_3  (keyAdd_port_state_out_8_0_3 ), //o
    .port_state_out_8_0_4  (keyAdd_port_state_out_8_0_4 ), //o
    .port_state_out_8_0_5  (keyAdd_port_state_out_8_0_5 ), //o
    .port_state_out_8_0_6  (keyAdd_port_state_out_8_0_6 ), //o
    .port_state_out_8_0_7  (keyAdd_port_state_out_8_0_7 ), //o
    .port_state_out_8_1_0  (keyAdd_port_state_out_8_1_0 ), //o
    .port_state_out_8_1_1  (keyAdd_port_state_out_8_1_1 ), //o
    .port_state_out_8_1_2  (keyAdd_port_state_out_8_1_2 ), //o
    .port_state_out_8_1_3  (keyAdd_port_state_out_8_1_3 ), //o
    .port_state_out_8_1_4  (keyAdd_port_state_out_8_1_4 ), //o
    .port_state_out_8_1_5  (keyAdd_port_state_out_8_1_5 ), //o
    .port_state_out_8_1_6  (keyAdd_port_state_out_8_1_6 ), //o
    .port_state_out_8_1_7  (keyAdd_port_state_out_8_1_7 ), //o
    .port_state_out_9_0_0  (keyAdd_port_state_out_9_0_0 ), //o
    .port_state_out_9_0_1  (keyAdd_port_state_out_9_0_1 ), //o
    .port_state_out_9_0_2  (keyAdd_port_state_out_9_0_2 ), //o
    .port_state_out_9_0_3  (keyAdd_port_state_out_9_0_3 ), //o
    .port_state_out_9_0_4  (keyAdd_port_state_out_9_0_4 ), //o
    .port_state_out_9_0_5  (keyAdd_port_state_out_9_0_5 ), //o
    .port_state_out_9_0_6  (keyAdd_port_state_out_9_0_6 ), //o
    .port_state_out_9_0_7  (keyAdd_port_state_out_9_0_7 ), //o
    .port_state_out_9_1_0  (keyAdd_port_state_out_9_1_0 ), //o
    .port_state_out_9_1_1  (keyAdd_port_state_out_9_1_1 ), //o
    .port_state_out_9_1_2  (keyAdd_port_state_out_9_1_2 ), //o
    .port_state_out_9_1_3  (keyAdd_port_state_out_9_1_3 ), //o
    .port_state_out_9_1_4  (keyAdd_port_state_out_9_1_4 ), //o
    .port_state_out_9_1_5  (keyAdd_port_state_out_9_1_5 ), //o
    .port_state_out_9_1_6  (keyAdd_port_state_out_9_1_6 ), //o
    .port_state_out_9_1_7  (keyAdd_port_state_out_9_1_7 ), //o
    .port_state_out_10_0_0 (keyAdd_port_state_out_10_0_0), //o
    .port_state_out_10_0_1 (keyAdd_port_state_out_10_0_1), //o
    .port_state_out_10_0_2 (keyAdd_port_state_out_10_0_2), //o
    .port_state_out_10_0_3 (keyAdd_port_state_out_10_0_3), //o
    .port_state_out_10_0_4 (keyAdd_port_state_out_10_0_4), //o
    .port_state_out_10_0_5 (keyAdd_port_state_out_10_0_5), //o
    .port_state_out_10_0_6 (keyAdd_port_state_out_10_0_6), //o
    .port_state_out_10_0_7 (keyAdd_port_state_out_10_0_7), //o
    .port_state_out_10_1_0 (keyAdd_port_state_out_10_1_0), //o
    .port_state_out_10_1_1 (keyAdd_port_state_out_10_1_1), //o
    .port_state_out_10_1_2 (keyAdd_port_state_out_10_1_2), //o
    .port_state_out_10_1_3 (keyAdd_port_state_out_10_1_3), //o
    .port_state_out_10_1_4 (keyAdd_port_state_out_10_1_4), //o
    .port_state_out_10_1_5 (keyAdd_port_state_out_10_1_5), //o
    .port_state_out_10_1_6 (keyAdd_port_state_out_10_1_6), //o
    .port_state_out_10_1_7 (keyAdd_port_state_out_10_1_7), //o
    .port_state_out_11_0_0 (keyAdd_port_state_out_11_0_0), //o
    .port_state_out_11_0_1 (keyAdd_port_state_out_11_0_1), //o
    .port_state_out_11_0_2 (keyAdd_port_state_out_11_0_2), //o
    .port_state_out_11_0_3 (keyAdd_port_state_out_11_0_3), //o
    .port_state_out_11_0_4 (keyAdd_port_state_out_11_0_4), //o
    .port_state_out_11_0_5 (keyAdd_port_state_out_11_0_5), //o
    .port_state_out_11_0_6 (keyAdd_port_state_out_11_0_6), //o
    .port_state_out_11_0_7 (keyAdd_port_state_out_11_0_7), //o
    .port_state_out_11_1_0 (keyAdd_port_state_out_11_1_0), //o
    .port_state_out_11_1_1 (keyAdd_port_state_out_11_1_1), //o
    .port_state_out_11_1_2 (keyAdd_port_state_out_11_1_2), //o
    .port_state_out_11_1_3 (keyAdd_port_state_out_11_1_3), //o
    .port_state_out_11_1_4 (keyAdd_port_state_out_11_1_4), //o
    .port_state_out_11_1_5 (keyAdd_port_state_out_11_1_5), //o
    .port_state_out_11_1_6 (keyAdd_port_state_out_11_1_6), //o
    .port_state_out_11_1_7 (keyAdd_port_state_out_11_1_7), //o
    .port_state_out_12_0_0 (keyAdd_port_state_out_12_0_0), //o
    .port_state_out_12_0_1 (keyAdd_port_state_out_12_0_1), //o
    .port_state_out_12_0_2 (keyAdd_port_state_out_12_0_2), //o
    .port_state_out_12_0_3 (keyAdd_port_state_out_12_0_3), //o
    .port_state_out_12_0_4 (keyAdd_port_state_out_12_0_4), //o
    .port_state_out_12_0_5 (keyAdd_port_state_out_12_0_5), //o
    .port_state_out_12_0_6 (keyAdd_port_state_out_12_0_6), //o
    .port_state_out_12_0_7 (keyAdd_port_state_out_12_0_7), //o
    .port_state_out_12_1_0 (keyAdd_port_state_out_12_1_0), //o
    .port_state_out_12_1_1 (keyAdd_port_state_out_12_1_1), //o
    .port_state_out_12_1_2 (keyAdd_port_state_out_12_1_2), //o
    .port_state_out_12_1_3 (keyAdd_port_state_out_12_1_3), //o
    .port_state_out_12_1_4 (keyAdd_port_state_out_12_1_4), //o
    .port_state_out_12_1_5 (keyAdd_port_state_out_12_1_5), //o
    .port_state_out_12_1_6 (keyAdd_port_state_out_12_1_6), //o
    .port_state_out_12_1_7 (keyAdd_port_state_out_12_1_7), //o
    .port_state_out_13_0_0 (keyAdd_port_state_out_13_0_0), //o
    .port_state_out_13_0_1 (keyAdd_port_state_out_13_0_1), //o
    .port_state_out_13_0_2 (keyAdd_port_state_out_13_0_2), //o
    .port_state_out_13_0_3 (keyAdd_port_state_out_13_0_3), //o
    .port_state_out_13_0_4 (keyAdd_port_state_out_13_0_4), //o
    .port_state_out_13_0_5 (keyAdd_port_state_out_13_0_5), //o
    .port_state_out_13_0_6 (keyAdd_port_state_out_13_0_6), //o
    .port_state_out_13_0_7 (keyAdd_port_state_out_13_0_7), //o
    .port_state_out_13_1_0 (keyAdd_port_state_out_13_1_0), //o
    .port_state_out_13_1_1 (keyAdd_port_state_out_13_1_1), //o
    .port_state_out_13_1_2 (keyAdd_port_state_out_13_1_2), //o
    .port_state_out_13_1_3 (keyAdd_port_state_out_13_1_3), //o
    .port_state_out_13_1_4 (keyAdd_port_state_out_13_1_4), //o
    .port_state_out_13_1_5 (keyAdd_port_state_out_13_1_5), //o
    .port_state_out_13_1_6 (keyAdd_port_state_out_13_1_6), //o
    .port_state_out_13_1_7 (keyAdd_port_state_out_13_1_7), //o
    .port_state_out_14_0_0 (keyAdd_port_state_out_14_0_0), //o
    .port_state_out_14_0_1 (keyAdd_port_state_out_14_0_1), //o
    .port_state_out_14_0_2 (keyAdd_port_state_out_14_0_2), //o
    .port_state_out_14_0_3 (keyAdd_port_state_out_14_0_3), //o
    .port_state_out_14_0_4 (keyAdd_port_state_out_14_0_4), //o
    .port_state_out_14_0_5 (keyAdd_port_state_out_14_0_5), //o
    .port_state_out_14_0_6 (keyAdd_port_state_out_14_0_6), //o
    .port_state_out_14_0_7 (keyAdd_port_state_out_14_0_7), //o
    .port_state_out_14_1_0 (keyAdd_port_state_out_14_1_0), //o
    .port_state_out_14_1_1 (keyAdd_port_state_out_14_1_1), //o
    .port_state_out_14_1_2 (keyAdd_port_state_out_14_1_2), //o
    .port_state_out_14_1_3 (keyAdd_port_state_out_14_1_3), //o
    .port_state_out_14_1_4 (keyAdd_port_state_out_14_1_4), //o
    .port_state_out_14_1_5 (keyAdd_port_state_out_14_1_5), //o
    .port_state_out_14_1_6 (keyAdd_port_state_out_14_1_6), //o
    .port_state_out_14_1_7 (keyAdd_port_state_out_14_1_7), //o
    .port_state_out_15_0_0 (keyAdd_port_state_out_15_0_0), //o
    .port_state_out_15_0_1 (keyAdd_port_state_out_15_0_1), //o
    .port_state_out_15_0_2 (keyAdd_port_state_out_15_0_2), //o
    .port_state_out_15_0_3 (keyAdd_port_state_out_15_0_3), //o
    .port_state_out_15_0_4 (keyAdd_port_state_out_15_0_4), //o
    .port_state_out_15_0_5 (keyAdd_port_state_out_15_0_5), //o
    .port_state_out_15_0_6 (keyAdd_port_state_out_15_0_6), //o
    .port_state_out_15_0_7 (keyAdd_port_state_out_15_0_7), //o
    .port_state_out_15_1_0 (keyAdd_port_state_out_15_1_0), //o
    .port_state_out_15_1_1 (keyAdd_port_state_out_15_1_1), //o
    .port_state_out_15_1_2 (keyAdd_port_state_out_15_1_2), //o
    .port_state_out_15_1_3 (keyAdd_port_state_out_15_1_3), //o
    .port_state_out_15_1_4 (keyAdd_port_state_out_15_1_4), //o
    .port_state_out_15_1_5 (keyAdd_port_state_out_15_1_5), //o
    .port_state_out_15_1_6 (keyAdd_port_state_out_15_1_6), //o
    .port_state_out_15_1_7 (keyAdd_port_state_out_15_1_7)  //o
  );
  Sbox_AES_Canright_CMS_2shares sbox_AES_Canright_CMS_2shares_16 (
    .port_i_0_0 (keyAdd_port_state_out_0_0_0                ), //i
    .port_i_0_1 (keyAdd_port_state_out_0_0_1                ), //i
    .port_i_0_2 (keyAdd_port_state_out_0_0_2                ), //i
    .port_i_0_3 (keyAdd_port_state_out_0_0_3                ), //i
    .port_i_0_4 (keyAdd_port_state_out_0_0_4                ), //i
    .port_i_0_5 (keyAdd_port_state_out_0_0_5                ), //i
    .port_i_0_6 (keyAdd_port_state_out_0_0_6                ), //i
    .port_i_0_7 (keyAdd_port_state_out_0_0_7                ), //i
    .port_i_1_0 (keyAdd_port_state_out_0_1_0                ), //i
    .port_i_1_1 (keyAdd_port_state_out_0_1_1                ), //i
    .port_i_1_2 (keyAdd_port_state_out_0_1_2                ), //i
    .port_i_1_3 (keyAdd_port_state_out_0_1_3                ), //i
    .port_i_1_4 (keyAdd_port_state_out_0_1_4                ), //i
    .port_i_1_5 (keyAdd_port_state_out_0_1_5                ), //i
    .port_i_1_6 (keyAdd_port_state_out_0_1_6                ), //i
    .port_i_1_7 (keyAdd_port_state_out_0_1_7                ), //i
    .port_r_0   (port_rand_0_0                              ), //i
    .port_r_1   (port_rand_0_1                              ), //i
    .port_r_2   (port_rand_0_2                              ), //i
    .port_r_3   (port_rand_0_3                              ), //i
    .port_r_4   (port_rand_0_4                              ), //i
    .port_r_5   (port_rand_0_5                              ), //i
    .port_r_6   (port_rand_0_6                              ), //i
    .port_r_7   (port_rand_0_7                              ), //i
    .port_r_8   (port_rand_0_8                              ), //i
    .port_r_9   (port_rand_0_9                              ), //i
    .port_r_10  (port_rand_0_10                             ), //i
    .port_r_11  (port_rand_0_11                             ), //i
    .port_r_12  (port_rand_0_12                             ), //i
    .port_r_13  (port_rand_0_13                             ), //i
    .port_r_14  (port_rand_0_14                             ), //i
    .port_r_15  (port_rand_0_15                             ), //i
    .port_r_16  (port_rand_0_16                             ), //i
    .port_r_17  (port_rand_0_17                             ), //i
    .port_r_18  (port_rand_0_18                             ), //i
    .port_r_19  (port_rand_0_19                             ), //i
    .port_r_20  (port_rand_0_20                             ), //i
    .port_r_21  (port_rand_0_21                             ), //i
    .port_r_22  (port_rand_0_22                             ), //i
    .port_r_23  (port_rand_0_23                             ), //i
    .port_r_24  (port_rand_0_24                             ), //i
    .port_r_25  (port_rand_0_25                             ), //i
    .port_r_26  (port_rand_0_26                             ), //i
    .port_r_27  (port_rand_0_27                             ), //i
    .port_r_28  (port_rand_0_28                             ), //i
    .port_r_29  (port_rand_0_29                             ), //i
    .port_r_30  (port_rand_0_30                             ), //i
    .port_r_31  (port_rand_0_31                             ), //i
    .port_r_32  (port_rand_0_32                             ), //i
    .port_r_33  (port_rand_0_33                             ), //i
    .port_r_34  (port_rand_0_34                             ), //i
    .port_r_35  (port_rand_0_35                             ), //i
    .port_r_36  (port_rand_0_36                             ), //i
    .port_r_37  (port_rand_0_37                             ), //i
    .port_r_38  (port_rand_0_38                             ), //i
    .port_r_39  (port_rand_0_39                             ), //i
    .port_r_40  (port_rand_0_40                             ), //i
    .port_r_41  (port_rand_0_41                             ), //i
    .port_r_42  (port_rand_0_42                             ), //i
    .port_r_43  (port_rand_0_43                             ), //i
    .port_r_44  (port_rand_0_44                             ), //i
    .port_r_45  (port_rand_0_45                             ), //i
    .port_r_46  (port_rand_0_46                             ), //i
    .port_r_47  (port_rand_0_47                             ), //i
    .port_r_48  (port_rand_0_48                             ), //i
    .port_r_49  (port_rand_0_49                             ), //i
    .port_r_50  (port_rand_0_50                             ), //i
    .port_r_51  (port_rand_0_51                             ), //i
    .port_r_52  (port_rand_0_52                             ), //i
    .port_r_53  (port_rand_0_53                             ), //i
    .port_o_0_0 (sbox_AES_Canright_CMS_2shares_16_port_o_0_0), //o
    .port_o_0_1 (sbox_AES_Canright_CMS_2shares_16_port_o_0_1), //o
    .port_o_0_2 (sbox_AES_Canright_CMS_2shares_16_port_o_0_2), //o
    .port_o_0_3 (sbox_AES_Canright_CMS_2shares_16_port_o_0_3), //o
    .port_o_0_4 (sbox_AES_Canright_CMS_2shares_16_port_o_0_4), //o
    .port_o_0_5 (sbox_AES_Canright_CMS_2shares_16_port_o_0_5), //o
    .port_o_0_6 (sbox_AES_Canright_CMS_2shares_16_port_o_0_6), //o
    .port_o_0_7 (sbox_AES_Canright_CMS_2shares_16_port_o_0_7), //o
    .port_o_1_0 (sbox_AES_Canright_CMS_2shares_16_port_o_1_0), //o
    .port_o_1_1 (sbox_AES_Canright_CMS_2shares_16_port_o_1_1), //o
    .port_o_1_2 (sbox_AES_Canright_CMS_2shares_16_port_o_1_2), //o
    .port_o_1_3 (sbox_AES_Canright_CMS_2shares_16_port_o_1_3), //o
    .port_o_1_4 (sbox_AES_Canright_CMS_2shares_16_port_o_1_4), //o
    .port_o_1_5 (sbox_AES_Canright_CMS_2shares_16_port_o_1_5), //o
    .port_o_1_6 (sbox_AES_Canright_CMS_2shares_16_port_o_1_6), //o
    .port_o_1_7 (sbox_AES_Canright_CMS_2shares_16_port_o_1_7), //o
    .clk        (clk                                        ), //i
    .reset      (reset                                      )  //i
  );
  Sbox_AES_Canright_CMS_2shares sbox_AES_Canright_CMS_2shares_17 (
    .port_i_0_0 (keyAdd_port_state_out_1_0_0                ), //i
    .port_i_0_1 (keyAdd_port_state_out_1_0_1                ), //i
    .port_i_0_2 (keyAdd_port_state_out_1_0_2                ), //i
    .port_i_0_3 (keyAdd_port_state_out_1_0_3                ), //i
    .port_i_0_4 (keyAdd_port_state_out_1_0_4                ), //i
    .port_i_0_5 (keyAdd_port_state_out_1_0_5                ), //i
    .port_i_0_6 (keyAdd_port_state_out_1_0_6                ), //i
    .port_i_0_7 (keyAdd_port_state_out_1_0_7                ), //i
    .port_i_1_0 (keyAdd_port_state_out_1_1_0                ), //i
    .port_i_1_1 (keyAdd_port_state_out_1_1_1                ), //i
    .port_i_1_2 (keyAdd_port_state_out_1_1_2                ), //i
    .port_i_1_3 (keyAdd_port_state_out_1_1_3                ), //i
    .port_i_1_4 (keyAdd_port_state_out_1_1_4                ), //i
    .port_i_1_5 (keyAdd_port_state_out_1_1_5                ), //i
    .port_i_1_6 (keyAdd_port_state_out_1_1_6                ), //i
    .port_i_1_7 (keyAdd_port_state_out_1_1_7                ), //i
    .port_r_0   (port_rand_1_0                              ), //i
    .port_r_1   (port_rand_1_1                              ), //i
    .port_r_2   (port_rand_1_2                              ), //i
    .port_r_3   (port_rand_1_3                              ), //i
    .port_r_4   (port_rand_1_4                              ), //i
    .port_r_5   (port_rand_1_5                              ), //i
    .port_r_6   (port_rand_1_6                              ), //i
    .port_r_7   (port_rand_1_7                              ), //i
    .port_r_8   (port_rand_1_8                              ), //i
    .port_r_9   (port_rand_1_9                              ), //i
    .port_r_10  (port_rand_1_10                             ), //i
    .port_r_11  (port_rand_1_11                             ), //i
    .port_r_12  (port_rand_1_12                             ), //i
    .port_r_13  (port_rand_1_13                             ), //i
    .port_r_14  (port_rand_1_14                             ), //i
    .port_r_15  (port_rand_1_15                             ), //i
    .port_r_16  (port_rand_1_16                             ), //i
    .port_r_17  (port_rand_1_17                             ), //i
    .port_r_18  (port_rand_1_18                             ), //i
    .port_r_19  (port_rand_1_19                             ), //i
    .port_r_20  (port_rand_1_20                             ), //i
    .port_r_21  (port_rand_1_21                             ), //i
    .port_r_22  (port_rand_1_22                             ), //i
    .port_r_23  (port_rand_1_23                             ), //i
    .port_r_24  (port_rand_1_24                             ), //i
    .port_r_25  (port_rand_1_25                             ), //i
    .port_r_26  (port_rand_1_26                             ), //i
    .port_r_27  (port_rand_1_27                             ), //i
    .port_r_28  (port_rand_1_28                             ), //i
    .port_r_29  (port_rand_1_29                             ), //i
    .port_r_30  (port_rand_1_30                             ), //i
    .port_r_31  (port_rand_1_31                             ), //i
    .port_r_32  (port_rand_1_32                             ), //i
    .port_r_33  (port_rand_1_33                             ), //i
    .port_r_34  (port_rand_1_34                             ), //i
    .port_r_35  (port_rand_1_35                             ), //i
    .port_r_36  (port_rand_1_36                             ), //i
    .port_r_37  (port_rand_1_37                             ), //i
    .port_r_38  (port_rand_1_38                             ), //i
    .port_r_39  (port_rand_1_39                             ), //i
    .port_r_40  (port_rand_1_40                             ), //i
    .port_r_41  (port_rand_1_41                             ), //i
    .port_r_42  (port_rand_1_42                             ), //i
    .port_r_43  (port_rand_1_43                             ), //i
    .port_r_44  (port_rand_1_44                             ), //i
    .port_r_45  (port_rand_1_45                             ), //i
    .port_r_46  (port_rand_1_46                             ), //i
    .port_r_47  (port_rand_1_47                             ), //i
    .port_r_48  (port_rand_1_48                             ), //i
    .port_r_49  (port_rand_1_49                             ), //i
    .port_r_50  (port_rand_1_50                             ), //i
    .port_r_51  (port_rand_1_51                             ), //i
    .port_r_52  (port_rand_1_52                             ), //i
    .port_r_53  (port_rand_1_53                             ), //i
    .port_o_0_0 (sbox_AES_Canright_CMS_2shares_17_port_o_0_0), //o
    .port_o_0_1 (sbox_AES_Canright_CMS_2shares_17_port_o_0_1), //o
    .port_o_0_2 (sbox_AES_Canright_CMS_2shares_17_port_o_0_2), //o
    .port_o_0_3 (sbox_AES_Canright_CMS_2shares_17_port_o_0_3), //o
    .port_o_0_4 (sbox_AES_Canright_CMS_2shares_17_port_o_0_4), //o
    .port_o_0_5 (sbox_AES_Canright_CMS_2shares_17_port_o_0_5), //o
    .port_o_0_6 (sbox_AES_Canright_CMS_2shares_17_port_o_0_6), //o
    .port_o_0_7 (sbox_AES_Canright_CMS_2shares_17_port_o_0_7), //o
    .port_o_1_0 (sbox_AES_Canright_CMS_2shares_17_port_o_1_0), //o
    .port_o_1_1 (sbox_AES_Canright_CMS_2shares_17_port_o_1_1), //o
    .port_o_1_2 (sbox_AES_Canright_CMS_2shares_17_port_o_1_2), //o
    .port_o_1_3 (sbox_AES_Canright_CMS_2shares_17_port_o_1_3), //o
    .port_o_1_4 (sbox_AES_Canright_CMS_2shares_17_port_o_1_4), //o
    .port_o_1_5 (sbox_AES_Canright_CMS_2shares_17_port_o_1_5), //o
    .port_o_1_6 (sbox_AES_Canright_CMS_2shares_17_port_o_1_6), //o
    .port_o_1_7 (sbox_AES_Canright_CMS_2shares_17_port_o_1_7), //o
    .clk        (clk                                        ), //i
    .reset      (reset                                      )  //i
  );
  Sbox_AES_Canright_CMS_2shares sbox_AES_Canright_CMS_2shares_18 (
    .port_i_0_0 (keyAdd_port_state_out_2_0_0                ), //i
    .port_i_0_1 (keyAdd_port_state_out_2_0_1                ), //i
    .port_i_0_2 (keyAdd_port_state_out_2_0_2                ), //i
    .port_i_0_3 (keyAdd_port_state_out_2_0_3                ), //i
    .port_i_0_4 (keyAdd_port_state_out_2_0_4                ), //i
    .port_i_0_5 (keyAdd_port_state_out_2_0_5                ), //i
    .port_i_0_6 (keyAdd_port_state_out_2_0_6                ), //i
    .port_i_0_7 (keyAdd_port_state_out_2_0_7                ), //i
    .port_i_1_0 (keyAdd_port_state_out_2_1_0                ), //i
    .port_i_1_1 (keyAdd_port_state_out_2_1_1                ), //i
    .port_i_1_2 (keyAdd_port_state_out_2_1_2                ), //i
    .port_i_1_3 (keyAdd_port_state_out_2_1_3                ), //i
    .port_i_1_4 (keyAdd_port_state_out_2_1_4                ), //i
    .port_i_1_5 (keyAdd_port_state_out_2_1_5                ), //i
    .port_i_1_6 (keyAdd_port_state_out_2_1_6                ), //i
    .port_i_1_7 (keyAdd_port_state_out_2_1_7                ), //i
    .port_r_0   (port_rand_2_0                              ), //i
    .port_r_1   (port_rand_2_1                              ), //i
    .port_r_2   (port_rand_2_2                              ), //i
    .port_r_3   (port_rand_2_3                              ), //i
    .port_r_4   (port_rand_2_4                              ), //i
    .port_r_5   (port_rand_2_5                              ), //i
    .port_r_6   (port_rand_2_6                              ), //i
    .port_r_7   (port_rand_2_7                              ), //i
    .port_r_8   (port_rand_2_8                              ), //i
    .port_r_9   (port_rand_2_9                              ), //i
    .port_r_10  (port_rand_2_10                             ), //i
    .port_r_11  (port_rand_2_11                             ), //i
    .port_r_12  (port_rand_2_12                             ), //i
    .port_r_13  (port_rand_2_13                             ), //i
    .port_r_14  (port_rand_2_14                             ), //i
    .port_r_15  (port_rand_2_15                             ), //i
    .port_r_16  (port_rand_2_16                             ), //i
    .port_r_17  (port_rand_2_17                             ), //i
    .port_r_18  (port_rand_2_18                             ), //i
    .port_r_19  (port_rand_2_19                             ), //i
    .port_r_20  (port_rand_2_20                             ), //i
    .port_r_21  (port_rand_2_21                             ), //i
    .port_r_22  (port_rand_2_22                             ), //i
    .port_r_23  (port_rand_2_23                             ), //i
    .port_r_24  (port_rand_2_24                             ), //i
    .port_r_25  (port_rand_2_25                             ), //i
    .port_r_26  (port_rand_2_26                             ), //i
    .port_r_27  (port_rand_2_27                             ), //i
    .port_r_28  (port_rand_2_28                             ), //i
    .port_r_29  (port_rand_2_29                             ), //i
    .port_r_30  (port_rand_2_30                             ), //i
    .port_r_31  (port_rand_2_31                             ), //i
    .port_r_32  (port_rand_2_32                             ), //i
    .port_r_33  (port_rand_2_33                             ), //i
    .port_r_34  (port_rand_2_34                             ), //i
    .port_r_35  (port_rand_2_35                             ), //i
    .port_r_36  (port_rand_2_36                             ), //i
    .port_r_37  (port_rand_2_37                             ), //i
    .port_r_38  (port_rand_2_38                             ), //i
    .port_r_39  (port_rand_2_39                             ), //i
    .port_r_40  (port_rand_2_40                             ), //i
    .port_r_41  (port_rand_2_41                             ), //i
    .port_r_42  (port_rand_2_42                             ), //i
    .port_r_43  (port_rand_2_43                             ), //i
    .port_r_44  (port_rand_2_44                             ), //i
    .port_r_45  (port_rand_2_45                             ), //i
    .port_r_46  (port_rand_2_46                             ), //i
    .port_r_47  (port_rand_2_47                             ), //i
    .port_r_48  (port_rand_2_48                             ), //i
    .port_r_49  (port_rand_2_49                             ), //i
    .port_r_50  (port_rand_2_50                             ), //i
    .port_r_51  (port_rand_2_51                             ), //i
    .port_r_52  (port_rand_2_52                             ), //i
    .port_r_53  (port_rand_2_53                             ), //i
    .port_o_0_0 (sbox_AES_Canright_CMS_2shares_18_port_o_0_0), //o
    .port_o_0_1 (sbox_AES_Canright_CMS_2shares_18_port_o_0_1), //o
    .port_o_0_2 (sbox_AES_Canright_CMS_2shares_18_port_o_0_2), //o
    .port_o_0_3 (sbox_AES_Canright_CMS_2shares_18_port_o_0_3), //o
    .port_o_0_4 (sbox_AES_Canright_CMS_2shares_18_port_o_0_4), //o
    .port_o_0_5 (sbox_AES_Canright_CMS_2shares_18_port_o_0_5), //o
    .port_o_0_6 (sbox_AES_Canright_CMS_2shares_18_port_o_0_6), //o
    .port_o_0_7 (sbox_AES_Canright_CMS_2shares_18_port_o_0_7), //o
    .port_o_1_0 (sbox_AES_Canright_CMS_2shares_18_port_o_1_0), //o
    .port_o_1_1 (sbox_AES_Canright_CMS_2shares_18_port_o_1_1), //o
    .port_o_1_2 (sbox_AES_Canright_CMS_2shares_18_port_o_1_2), //o
    .port_o_1_3 (sbox_AES_Canright_CMS_2shares_18_port_o_1_3), //o
    .port_o_1_4 (sbox_AES_Canright_CMS_2shares_18_port_o_1_4), //o
    .port_o_1_5 (sbox_AES_Canright_CMS_2shares_18_port_o_1_5), //o
    .port_o_1_6 (sbox_AES_Canright_CMS_2shares_18_port_o_1_6), //o
    .port_o_1_7 (sbox_AES_Canright_CMS_2shares_18_port_o_1_7), //o
    .clk        (clk                                        ), //i
    .reset      (reset                                      )  //i
  );
  Sbox_AES_Canright_CMS_2shares sbox_AES_Canright_CMS_2shares_19 (
    .port_i_0_0 (keyAdd_port_state_out_3_0_0                ), //i
    .port_i_0_1 (keyAdd_port_state_out_3_0_1                ), //i
    .port_i_0_2 (keyAdd_port_state_out_3_0_2                ), //i
    .port_i_0_3 (keyAdd_port_state_out_3_0_3                ), //i
    .port_i_0_4 (keyAdd_port_state_out_3_0_4                ), //i
    .port_i_0_5 (keyAdd_port_state_out_3_0_5                ), //i
    .port_i_0_6 (keyAdd_port_state_out_3_0_6                ), //i
    .port_i_0_7 (keyAdd_port_state_out_3_0_7                ), //i
    .port_i_1_0 (keyAdd_port_state_out_3_1_0                ), //i
    .port_i_1_1 (keyAdd_port_state_out_3_1_1                ), //i
    .port_i_1_2 (keyAdd_port_state_out_3_1_2                ), //i
    .port_i_1_3 (keyAdd_port_state_out_3_1_3                ), //i
    .port_i_1_4 (keyAdd_port_state_out_3_1_4                ), //i
    .port_i_1_5 (keyAdd_port_state_out_3_1_5                ), //i
    .port_i_1_6 (keyAdd_port_state_out_3_1_6                ), //i
    .port_i_1_7 (keyAdd_port_state_out_3_1_7                ), //i
    .port_r_0   (port_rand_3_0                              ), //i
    .port_r_1   (port_rand_3_1                              ), //i
    .port_r_2   (port_rand_3_2                              ), //i
    .port_r_3   (port_rand_3_3                              ), //i
    .port_r_4   (port_rand_3_4                              ), //i
    .port_r_5   (port_rand_3_5                              ), //i
    .port_r_6   (port_rand_3_6                              ), //i
    .port_r_7   (port_rand_3_7                              ), //i
    .port_r_8   (port_rand_3_8                              ), //i
    .port_r_9   (port_rand_3_9                              ), //i
    .port_r_10  (port_rand_3_10                             ), //i
    .port_r_11  (port_rand_3_11                             ), //i
    .port_r_12  (port_rand_3_12                             ), //i
    .port_r_13  (port_rand_3_13                             ), //i
    .port_r_14  (port_rand_3_14                             ), //i
    .port_r_15  (port_rand_3_15                             ), //i
    .port_r_16  (port_rand_3_16                             ), //i
    .port_r_17  (port_rand_3_17                             ), //i
    .port_r_18  (port_rand_3_18                             ), //i
    .port_r_19  (port_rand_3_19                             ), //i
    .port_r_20  (port_rand_3_20                             ), //i
    .port_r_21  (port_rand_3_21                             ), //i
    .port_r_22  (port_rand_3_22                             ), //i
    .port_r_23  (port_rand_3_23                             ), //i
    .port_r_24  (port_rand_3_24                             ), //i
    .port_r_25  (port_rand_3_25                             ), //i
    .port_r_26  (port_rand_3_26                             ), //i
    .port_r_27  (port_rand_3_27                             ), //i
    .port_r_28  (port_rand_3_28                             ), //i
    .port_r_29  (port_rand_3_29                             ), //i
    .port_r_30  (port_rand_3_30                             ), //i
    .port_r_31  (port_rand_3_31                             ), //i
    .port_r_32  (port_rand_3_32                             ), //i
    .port_r_33  (port_rand_3_33                             ), //i
    .port_r_34  (port_rand_3_34                             ), //i
    .port_r_35  (port_rand_3_35                             ), //i
    .port_r_36  (port_rand_3_36                             ), //i
    .port_r_37  (port_rand_3_37                             ), //i
    .port_r_38  (port_rand_3_38                             ), //i
    .port_r_39  (port_rand_3_39                             ), //i
    .port_r_40  (port_rand_3_40                             ), //i
    .port_r_41  (port_rand_3_41                             ), //i
    .port_r_42  (port_rand_3_42                             ), //i
    .port_r_43  (port_rand_3_43                             ), //i
    .port_r_44  (port_rand_3_44                             ), //i
    .port_r_45  (port_rand_3_45                             ), //i
    .port_r_46  (port_rand_3_46                             ), //i
    .port_r_47  (port_rand_3_47                             ), //i
    .port_r_48  (port_rand_3_48                             ), //i
    .port_r_49  (port_rand_3_49                             ), //i
    .port_r_50  (port_rand_3_50                             ), //i
    .port_r_51  (port_rand_3_51                             ), //i
    .port_r_52  (port_rand_3_52                             ), //i
    .port_r_53  (port_rand_3_53                             ), //i
    .port_o_0_0 (sbox_AES_Canright_CMS_2shares_19_port_o_0_0), //o
    .port_o_0_1 (sbox_AES_Canright_CMS_2shares_19_port_o_0_1), //o
    .port_o_0_2 (sbox_AES_Canright_CMS_2shares_19_port_o_0_2), //o
    .port_o_0_3 (sbox_AES_Canright_CMS_2shares_19_port_o_0_3), //o
    .port_o_0_4 (sbox_AES_Canright_CMS_2shares_19_port_o_0_4), //o
    .port_o_0_5 (sbox_AES_Canright_CMS_2shares_19_port_o_0_5), //o
    .port_o_0_6 (sbox_AES_Canright_CMS_2shares_19_port_o_0_6), //o
    .port_o_0_7 (sbox_AES_Canright_CMS_2shares_19_port_o_0_7), //o
    .port_o_1_0 (sbox_AES_Canright_CMS_2shares_19_port_o_1_0), //o
    .port_o_1_1 (sbox_AES_Canright_CMS_2shares_19_port_o_1_1), //o
    .port_o_1_2 (sbox_AES_Canright_CMS_2shares_19_port_o_1_2), //o
    .port_o_1_3 (sbox_AES_Canright_CMS_2shares_19_port_o_1_3), //o
    .port_o_1_4 (sbox_AES_Canright_CMS_2shares_19_port_o_1_4), //o
    .port_o_1_5 (sbox_AES_Canright_CMS_2shares_19_port_o_1_5), //o
    .port_o_1_6 (sbox_AES_Canright_CMS_2shares_19_port_o_1_6), //o
    .port_o_1_7 (sbox_AES_Canright_CMS_2shares_19_port_o_1_7), //o
    .clk        (clk                                        ), //i
    .reset      (reset                                      )  //i
  );
  Sbox_AES_Canright_CMS_2shares sbox_AES_Canright_CMS_2shares_20 (
    .port_i_0_0 (keyAdd_port_state_out_4_0_0                ), //i
    .port_i_0_1 (keyAdd_port_state_out_4_0_1                ), //i
    .port_i_0_2 (keyAdd_port_state_out_4_0_2                ), //i
    .port_i_0_3 (keyAdd_port_state_out_4_0_3                ), //i
    .port_i_0_4 (keyAdd_port_state_out_4_0_4                ), //i
    .port_i_0_5 (keyAdd_port_state_out_4_0_5                ), //i
    .port_i_0_6 (keyAdd_port_state_out_4_0_6                ), //i
    .port_i_0_7 (keyAdd_port_state_out_4_0_7                ), //i
    .port_i_1_0 (keyAdd_port_state_out_4_1_0                ), //i
    .port_i_1_1 (keyAdd_port_state_out_4_1_1                ), //i
    .port_i_1_2 (keyAdd_port_state_out_4_1_2                ), //i
    .port_i_1_3 (keyAdd_port_state_out_4_1_3                ), //i
    .port_i_1_4 (keyAdd_port_state_out_4_1_4                ), //i
    .port_i_1_5 (keyAdd_port_state_out_4_1_5                ), //i
    .port_i_1_6 (keyAdd_port_state_out_4_1_6                ), //i
    .port_i_1_7 (keyAdd_port_state_out_4_1_7                ), //i
    .port_r_0   (port_rand_4_0                              ), //i
    .port_r_1   (port_rand_4_1                              ), //i
    .port_r_2   (port_rand_4_2                              ), //i
    .port_r_3   (port_rand_4_3                              ), //i
    .port_r_4   (port_rand_4_4                              ), //i
    .port_r_5   (port_rand_4_5                              ), //i
    .port_r_6   (port_rand_4_6                              ), //i
    .port_r_7   (port_rand_4_7                              ), //i
    .port_r_8   (port_rand_4_8                              ), //i
    .port_r_9   (port_rand_4_9                              ), //i
    .port_r_10  (port_rand_4_10                             ), //i
    .port_r_11  (port_rand_4_11                             ), //i
    .port_r_12  (port_rand_4_12                             ), //i
    .port_r_13  (port_rand_4_13                             ), //i
    .port_r_14  (port_rand_4_14                             ), //i
    .port_r_15  (port_rand_4_15                             ), //i
    .port_r_16  (port_rand_4_16                             ), //i
    .port_r_17  (port_rand_4_17                             ), //i
    .port_r_18  (port_rand_4_18                             ), //i
    .port_r_19  (port_rand_4_19                             ), //i
    .port_r_20  (port_rand_4_20                             ), //i
    .port_r_21  (port_rand_4_21                             ), //i
    .port_r_22  (port_rand_4_22                             ), //i
    .port_r_23  (port_rand_4_23                             ), //i
    .port_r_24  (port_rand_4_24                             ), //i
    .port_r_25  (port_rand_4_25                             ), //i
    .port_r_26  (port_rand_4_26                             ), //i
    .port_r_27  (port_rand_4_27                             ), //i
    .port_r_28  (port_rand_4_28                             ), //i
    .port_r_29  (port_rand_4_29                             ), //i
    .port_r_30  (port_rand_4_30                             ), //i
    .port_r_31  (port_rand_4_31                             ), //i
    .port_r_32  (port_rand_4_32                             ), //i
    .port_r_33  (port_rand_4_33                             ), //i
    .port_r_34  (port_rand_4_34                             ), //i
    .port_r_35  (port_rand_4_35                             ), //i
    .port_r_36  (port_rand_4_36                             ), //i
    .port_r_37  (port_rand_4_37                             ), //i
    .port_r_38  (port_rand_4_38                             ), //i
    .port_r_39  (port_rand_4_39                             ), //i
    .port_r_40  (port_rand_4_40                             ), //i
    .port_r_41  (port_rand_4_41                             ), //i
    .port_r_42  (port_rand_4_42                             ), //i
    .port_r_43  (port_rand_4_43                             ), //i
    .port_r_44  (port_rand_4_44                             ), //i
    .port_r_45  (port_rand_4_45                             ), //i
    .port_r_46  (port_rand_4_46                             ), //i
    .port_r_47  (port_rand_4_47                             ), //i
    .port_r_48  (port_rand_4_48                             ), //i
    .port_r_49  (port_rand_4_49                             ), //i
    .port_r_50  (port_rand_4_50                             ), //i
    .port_r_51  (port_rand_4_51                             ), //i
    .port_r_52  (port_rand_4_52                             ), //i
    .port_r_53  (port_rand_4_53                             ), //i
    .port_o_0_0 (sbox_AES_Canright_CMS_2shares_20_port_o_0_0), //o
    .port_o_0_1 (sbox_AES_Canright_CMS_2shares_20_port_o_0_1), //o
    .port_o_0_2 (sbox_AES_Canright_CMS_2shares_20_port_o_0_2), //o
    .port_o_0_3 (sbox_AES_Canright_CMS_2shares_20_port_o_0_3), //o
    .port_o_0_4 (sbox_AES_Canright_CMS_2shares_20_port_o_0_4), //o
    .port_o_0_5 (sbox_AES_Canright_CMS_2shares_20_port_o_0_5), //o
    .port_o_0_6 (sbox_AES_Canright_CMS_2shares_20_port_o_0_6), //o
    .port_o_0_7 (sbox_AES_Canright_CMS_2shares_20_port_o_0_7), //o
    .port_o_1_0 (sbox_AES_Canright_CMS_2shares_20_port_o_1_0), //o
    .port_o_1_1 (sbox_AES_Canright_CMS_2shares_20_port_o_1_1), //o
    .port_o_1_2 (sbox_AES_Canright_CMS_2shares_20_port_o_1_2), //o
    .port_o_1_3 (sbox_AES_Canright_CMS_2shares_20_port_o_1_3), //o
    .port_o_1_4 (sbox_AES_Canright_CMS_2shares_20_port_o_1_4), //o
    .port_o_1_5 (sbox_AES_Canright_CMS_2shares_20_port_o_1_5), //o
    .port_o_1_6 (sbox_AES_Canright_CMS_2shares_20_port_o_1_6), //o
    .port_o_1_7 (sbox_AES_Canright_CMS_2shares_20_port_o_1_7), //o
    .clk        (clk                                        ), //i
    .reset      (reset                                      )  //i
  );
  Sbox_AES_Canright_CMS_2shares sbox_AES_Canright_CMS_2shares_21 (
    .port_i_0_0 (keyAdd_port_state_out_5_0_0                ), //i
    .port_i_0_1 (keyAdd_port_state_out_5_0_1                ), //i
    .port_i_0_2 (keyAdd_port_state_out_5_0_2                ), //i
    .port_i_0_3 (keyAdd_port_state_out_5_0_3                ), //i
    .port_i_0_4 (keyAdd_port_state_out_5_0_4                ), //i
    .port_i_0_5 (keyAdd_port_state_out_5_0_5                ), //i
    .port_i_0_6 (keyAdd_port_state_out_5_0_6                ), //i
    .port_i_0_7 (keyAdd_port_state_out_5_0_7                ), //i
    .port_i_1_0 (keyAdd_port_state_out_5_1_0                ), //i
    .port_i_1_1 (keyAdd_port_state_out_5_1_1                ), //i
    .port_i_1_2 (keyAdd_port_state_out_5_1_2                ), //i
    .port_i_1_3 (keyAdd_port_state_out_5_1_3                ), //i
    .port_i_1_4 (keyAdd_port_state_out_5_1_4                ), //i
    .port_i_1_5 (keyAdd_port_state_out_5_1_5                ), //i
    .port_i_1_6 (keyAdd_port_state_out_5_1_6                ), //i
    .port_i_1_7 (keyAdd_port_state_out_5_1_7                ), //i
    .port_r_0   (port_rand_5_0                              ), //i
    .port_r_1   (port_rand_5_1                              ), //i
    .port_r_2   (port_rand_5_2                              ), //i
    .port_r_3   (port_rand_5_3                              ), //i
    .port_r_4   (port_rand_5_4                              ), //i
    .port_r_5   (port_rand_5_5                              ), //i
    .port_r_6   (port_rand_5_6                              ), //i
    .port_r_7   (port_rand_5_7                              ), //i
    .port_r_8   (port_rand_5_8                              ), //i
    .port_r_9   (port_rand_5_9                              ), //i
    .port_r_10  (port_rand_5_10                             ), //i
    .port_r_11  (port_rand_5_11                             ), //i
    .port_r_12  (port_rand_5_12                             ), //i
    .port_r_13  (port_rand_5_13                             ), //i
    .port_r_14  (port_rand_5_14                             ), //i
    .port_r_15  (port_rand_5_15                             ), //i
    .port_r_16  (port_rand_5_16                             ), //i
    .port_r_17  (port_rand_5_17                             ), //i
    .port_r_18  (port_rand_5_18                             ), //i
    .port_r_19  (port_rand_5_19                             ), //i
    .port_r_20  (port_rand_5_20                             ), //i
    .port_r_21  (port_rand_5_21                             ), //i
    .port_r_22  (port_rand_5_22                             ), //i
    .port_r_23  (port_rand_5_23                             ), //i
    .port_r_24  (port_rand_5_24                             ), //i
    .port_r_25  (port_rand_5_25                             ), //i
    .port_r_26  (port_rand_5_26                             ), //i
    .port_r_27  (port_rand_5_27                             ), //i
    .port_r_28  (port_rand_5_28                             ), //i
    .port_r_29  (port_rand_5_29                             ), //i
    .port_r_30  (port_rand_5_30                             ), //i
    .port_r_31  (port_rand_5_31                             ), //i
    .port_r_32  (port_rand_5_32                             ), //i
    .port_r_33  (port_rand_5_33                             ), //i
    .port_r_34  (port_rand_5_34                             ), //i
    .port_r_35  (port_rand_5_35                             ), //i
    .port_r_36  (port_rand_5_36                             ), //i
    .port_r_37  (port_rand_5_37                             ), //i
    .port_r_38  (port_rand_5_38                             ), //i
    .port_r_39  (port_rand_5_39                             ), //i
    .port_r_40  (port_rand_5_40                             ), //i
    .port_r_41  (port_rand_5_41                             ), //i
    .port_r_42  (port_rand_5_42                             ), //i
    .port_r_43  (port_rand_5_43                             ), //i
    .port_r_44  (port_rand_5_44                             ), //i
    .port_r_45  (port_rand_5_45                             ), //i
    .port_r_46  (port_rand_5_46                             ), //i
    .port_r_47  (port_rand_5_47                             ), //i
    .port_r_48  (port_rand_5_48                             ), //i
    .port_r_49  (port_rand_5_49                             ), //i
    .port_r_50  (port_rand_5_50                             ), //i
    .port_r_51  (port_rand_5_51                             ), //i
    .port_r_52  (port_rand_5_52                             ), //i
    .port_r_53  (port_rand_5_53                             ), //i
    .port_o_0_0 (sbox_AES_Canright_CMS_2shares_21_port_o_0_0), //o
    .port_o_0_1 (sbox_AES_Canright_CMS_2shares_21_port_o_0_1), //o
    .port_o_0_2 (sbox_AES_Canright_CMS_2shares_21_port_o_0_2), //o
    .port_o_0_3 (sbox_AES_Canright_CMS_2shares_21_port_o_0_3), //o
    .port_o_0_4 (sbox_AES_Canright_CMS_2shares_21_port_o_0_4), //o
    .port_o_0_5 (sbox_AES_Canright_CMS_2shares_21_port_o_0_5), //o
    .port_o_0_6 (sbox_AES_Canright_CMS_2shares_21_port_o_0_6), //o
    .port_o_0_7 (sbox_AES_Canright_CMS_2shares_21_port_o_0_7), //o
    .port_o_1_0 (sbox_AES_Canright_CMS_2shares_21_port_o_1_0), //o
    .port_o_1_1 (sbox_AES_Canright_CMS_2shares_21_port_o_1_1), //o
    .port_o_1_2 (sbox_AES_Canright_CMS_2shares_21_port_o_1_2), //o
    .port_o_1_3 (sbox_AES_Canright_CMS_2shares_21_port_o_1_3), //o
    .port_o_1_4 (sbox_AES_Canright_CMS_2shares_21_port_o_1_4), //o
    .port_o_1_5 (sbox_AES_Canright_CMS_2shares_21_port_o_1_5), //o
    .port_o_1_6 (sbox_AES_Canright_CMS_2shares_21_port_o_1_6), //o
    .port_o_1_7 (sbox_AES_Canright_CMS_2shares_21_port_o_1_7), //o
    .clk        (clk                                        ), //i
    .reset      (reset                                      )  //i
  );
  Sbox_AES_Canright_CMS_2shares sbox_AES_Canright_CMS_2shares_22 (
    .port_i_0_0 (keyAdd_port_state_out_6_0_0                ), //i
    .port_i_0_1 (keyAdd_port_state_out_6_0_1                ), //i
    .port_i_0_2 (keyAdd_port_state_out_6_0_2                ), //i
    .port_i_0_3 (keyAdd_port_state_out_6_0_3                ), //i
    .port_i_0_4 (keyAdd_port_state_out_6_0_4                ), //i
    .port_i_0_5 (keyAdd_port_state_out_6_0_5                ), //i
    .port_i_0_6 (keyAdd_port_state_out_6_0_6                ), //i
    .port_i_0_7 (keyAdd_port_state_out_6_0_7                ), //i
    .port_i_1_0 (keyAdd_port_state_out_6_1_0                ), //i
    .port_i_1_1 (keyAdd_port_state_out_6_1_1                ), //i
    .port_i_1_2 (keyAdd_port_state_out_6_1_2                ), //i
    .port_i_1_3 (keyAdd_port_state_out_6_1_3                ), //i
    .port_i_1_4 (keyAdd_port_state_out_6_1_4                ), //i
    .port_i_1_5 (keyAdd_port_state_out_6_1_5                ), //i
    .port_i_1_6 (keyAdd_port_state_out_6_1_6                ), //i
    .port_i_1_7 (keyAdd_port_state_out_6_1_7                ), //i
    .port_r_0   (port_rand_6_0                              ), //i
    .port_r_1   (port_rand_6_1                              ), //i
    .port_r_2   (port_rand_6_2                              ), //i
    .port_r_3   (port_rand_6_3                              ), //i
    .port_r_4   (port_rand_6_4                              ), //i
    .port_r_5   (port_rand_6_5                              ), //i
    .port_r_6   (port_rand_6_6                              ), //i
    .port_r_7   (port_rand_6_7                              ), //i
    .port_r_8   (port_rand_6_8                              ), //i
    .port_r_9   (port_rand_6_9                              ), //i
    .port_r_10  (port_rand_6_10                             ), //i
    .port_r_11  (port_rand_6_11                             ), //i
    .port_r_12  (port_rand_6_12                             ), //i
    .port_r_13  (port_rand_6_13                             ), //i
    .port_r_14  (port_rand_6_14                             ), //i
    .port_r_15  (port_rand_6_15                             ), //i
    .port_r_16  (port_rand_6_16                             ), //i
    .port_r_17  (port_rand_6_17                             ), //i
    .port_r_18  (port_rand_6_18                             ), //i
    .port_r_19  (port_rand_6_19                             ), //i
    .port_r_20  (port_rand_6_20                             ), //i
    .port_r_21  (port_rand_6_21                             ), //i
    .port_r_22  (port_rand_6_22                             ), //i
    .port_r_23  (port_rand_6_23                             ), //i
    .port_r_24  (port_rand_6_24                             ), //i
    .port_r_25  (port_rand_6_25                             ), //i
    .port_r_26  (port_rand_6_26                             ), //i
    .port_r_27  (port_rand_6_27                             ), //i
    .port_r_28  (port_rand_6_28                             ), //i
    .port_r_29  (port_rand_6_29                             ), //i
    .port_r_30  (port_rand_6_30                             ), //i
    .port_r_31  (port_rand_6_31                             ), //i
    .port_r_32  (port_rand_6_32                             ), //i
    .port_r_33  (port_rand_6_33                             ), //i
    .port_r_34  (port_rand_6_34                             ), //i
    .port_r_35  (port_rand_6_35                             ), //i
    .port_r_36  (port_rand_6_36                             ), //i
    .port_r_37  (port_rand_6_37                             ), //i
    .port_r_38  (port_rand_6_38                             ), //i
    .port_r_39  (port_rand_6_39                             ), //i
    .port_r_40  (port_rand_6_40                             ), //i
    .port_r_41  (port_rand_6_41                             ), //i
    .port_r_42  (port_rand_6_42                             ), //i
    .port_r_43  (port_rand_6_43                             ), //i
    .port_r_44  (port_rand_6_44                             ), //i
    .port_r_45  (port_rand_6_45                             ), //i
    .port_r_46  (port_rand_6_46                             ), //i
    .port_r_47  (port_rand_6_47                             ), //i
    .port_r_48  (port_rand_6_48                             ), //i
    .port_r_49  (port_rand_6_49                             ), //i
    .port_r_50  (port_rand_6_50                             ), //i
    .port_r_51  (port_rand_6_51                             ), //i
    .port_r_52  (port_rand_6_52                             ), //i
    .port_r_53  (port_rand_6_53                             ), //i
    .port_o_0_0 (sbox_AES_Canright_CMS_2shares_22_port_o_0_0), //o
    .port_o_0_1 (sbox_AES_Canright_CMS_2shares_22_port_o_0_1), //o
    .port_o_0_2 (sbox_AES_Canright_CMS_2shares_22_port_o_0_2), //o
    .port_o_0_3 (sbox_AES_Canright_CMS_2shares_22_port_o_0_3), //o
    .port_o_0_4 (sbox_AES_Canright_CMS_2shares_22_port_o_0_4), //o
    .port_o_0_5 (sbox_AES_Canright_CMS_2shares_22_port_o_0_5), //o
    .port_o_0_6 (sbox_AES_Canright_CMS_2shares_22_port_o_0_6), //o
    .port_o_0_7 (sbox_AES_Canright_CMS_2shares_22_port_o_0_7), //o
    .port_o_1_0 (sbox_AES_Canright_CMS_2shares_22_port_o_1_0), //o
    .port_o_1_1 (sbox_AES_Canright_CMS_2shares_22_port_o_1_1), //o
    .port_o_1_2 (sbox_AES_Canright_CMS_2shares_22_port_o_1_2), //o
    .port_o_1_3 (sbox_AES_Canright_CMS_2shares_22_port_o_1_3), //o
    .port_o_1_4 (sbox_AES_Canright_CMS_2shares_22_port_o_1_4), //o
    .port_o_1_5 (sbox_AES_Canright_CMS_2shares_22_port_o_1_5), //o
    .port_o_1_6 (sbox_AES_Canright_CMS_2shares_22_port_o_1_6), //o
    .port_o_1_7 (sbox_AES_Canright_CMS_2shares_22_port_o_1_7), //o
    .clk        (clk                                        ), //i
    .reset      (reset                                      )  //i
  );
  Sbox_AES_Canright_CMS_2shares sbox_AES_Canright_CMS_2shares_23 (
    .port_i_0_0 (keyAdd_port_state_out_7_0_0                ), //i
    .port_i_0_1 (keyAdd_port_state_out_7_0_1                ), //i
    .port_i_0_2 (keyAdd_port_state_out_7_0_2                ), //i
    .port_i_0_3 (keyAdd_port_state_out_7_0_3                ), //i
    .port_i_0_4 (keyAdd_port_state_out_7_0_4                ), //i
    .port_i_0_5 (keyAdd_port_state_out_7_0_5                ), //i
    .port_i_0_6 (keyAdd_port_state_out_7_0_6                ), //i
    .port_i_0_7 (keyAdd_port_state_out_7_0_7                ), //i
    .port_i_1_0 (keyAdd_port_state_out_7_1_0                ), //i
    .port_i_1_1 (keyAdd_port_state_out_7_1_1                ), //i
    .port_i_1_2 (keyAdd_port_state_out_7_1_2                ), //i
    .port_i_1_3 (keyAdd_port_state_out_7_1_3                ), //i
    .port_i_1_4 (keyAdd_port_state_out_7_1_4                ), //i
    .port_i_1_5 (keyAdd_port_state_out_7_1_5                ), //i
    .port_i_1_6 (keyAdd_port_state_out_7_1_6                ), //i
    .port_i_1_7 (keyAdd_port_state_out_7_1_7                ), //i
    .port_r_0   (port_rand_7_0                              ), //i
    .port_r_1   (port_rand_7_1                              ), //i
    .port_r_2   (port_rand_7_2                              ), //i
    .port_r_3   (port_rand_7_3                              ), //i
    .port_r_4   (port_rand_7_4                              ), //i
    .port_r_5   (port_rand_7_5                              ), //i
    .port_r_6   (port_rand_7_6                              ), //i
    .port_r_7   (port_rand_7_7                              ), //i
    .port_r_8   (port_rand_7_8                              ), //i
    .port_r_9   (port_rand_7_9                              ), //i
    .port_r_10  (port_rand_7_10                             ), //i
    .port_r_11  (port_rand_7_11                             ), //i
    .port_r_12  (port_rand_7_12                             ), //i
    .port_r_13  (port_rand_7_13                             ), //i
    .port_r_14  (port_rand_7_14                             ), //i
    .port_r_15  (port_rand_7_15                             ), //i
    .port_r_16  (port_rand_7_16                             ), //i
    .port_r_17  (port_rand_7_17                             ), //i
    .port_r_18  (port_rand_7_18                             ), //i
    .port_r_19  (port_rand_7_19                             ), //i
    .port_r_20  (port_rand_7_20                             ), //i
    .port_r_21  (port_rand_7_21                             ), //i
    .port_r_22  (port_rand_7_22                             ), //i
    .port_r_23  (port_rand_7_23                             ), //i
    .port_r_24  (port_rand_7_24                             ), //i
    .port_r_25  (port_rand_7_25                             ), //i
    .port_r_26  (port_rand_7_26                             ), //i
    .port_r_27  (port_rand_7_27                             ), //i
    .port_r_28  (port_rand_7_28                             ), //i
    .port_r_29  (port_rand_7_29                             ), //i
    .port_r_30  (port_rand_7_30                             ), //i
    .port_r_31  (port_rand_7_31                             ), //i
    .port_r_32  (port_rand_7_32                             ), //i
    .port_r_33  (port_rand_7_33                             ), //i
    .port_r_34  (port_rand_7_34                             ), //i
    .port_r_35  (port_rand_7_35                             ), //i
    .port_r_36  (port_rand_7_36                             ), //i
    .port_r_37  (port_rand_7_37                             ), //i
    .port_r_38  (port_rand_7_38                             ), //i
    .port_r_39  (port_rand_7_39                             ), //i
    .port_r_40  (port_rand_7_40                             ), //i
    .port_r_41  (port_rand_7_41                             ), //i
    .port_r_42  (port_rand_7_42                             ), //i
    .port_r_43  (port_rand_7_43                             ), //i
    .port_r_44  (port_rand_7_44                             ), //i
    .port_r_45  (port_rand_7_45                             ), //i
    .port_r_46  (port_rand_7_46                             ), //i
    .port_r_47  (port_rand_7_47                             ), //i
    .port_r_48  (port_rand_7_48                             ), //i
    .port_r_49  (port_rand_7_49                             ), //i
    .port_r_50  (port_rand_7_50                             ), //i
    .port_r_51  (port_rand_7_51                             ), //i
    .port_r_52  (port_rand_7_52                             ), //i
    .port_r_53  (port_rand_7_53                             ), //i
    .port_o_0_0 (sbox_AES_Canright_CMS_2shares_23_port_o_0_0), //o
    .port_o_0_1 (sbox_AES_Canright_CMS_2shares_23_port_o_0_1), //o
    .port_o_0_2 (sbox_AES_Canright_CMS_2shares_23_port_o_0_2), //o
    .port_o_0_3 (sbox_AES_Canright_CMS_2shares_23_port_o_0_3), //o
    .port_o_0_4 (sbox_AES_Canright_CMS_2shares_23_port_o_0_4), //o
    .port_o_0_5 (sbox_AES_Canright_CMS_2shares_23_port_o_0_5), //o
    .port_o_0_6 (sbox_AES_Canright_CMS_2shares_23_port_o_0_6), //o
    .port_o_0_7 (sbox_AES_Canright_CMS_2shares_23_port_o_0_7), //o
    .port_o_1_0 (sbox_AES_Canright_CMS_2shares_23_port_o_1_0), //o
    .port_o_1_1 (sbox_AES_Canright_CMS_2shares_23_port_o_1_1), //o
    .port_o_1_2 (sbox_AES_Canright_CMS_2shares_23_port_o_1_2), //o
    .port_o_1_3 (sbox_AES_Canright_CMS_2shares_23_port_o_1_3), //o
    .port_o_1_4 (sbox_AES_Canright_CMS_2shares_23_port_o_1_4), //o
    .port_o_1_5 (sbox_AES_Canright_CMS_2shares_23_port_o_1_5), //o
    .port_o_1_6 (sbox_AES_Canright_CMS_2shares_23_port_o_1_6), //o
    .port_o_1_7 (sbox_AES_Canright_CMS_2shares_23_port_o_1_7), //o
    .clk        (clk                                        ), //i
    .reset      (reset                                      )  //i
  );
  Sbox_AES_Canright_CMS_2shares sbox_AES_Canright_CMS_2shares_24 (
    .port_i_0_0 (keyAdd_port_state_out_8_0_0                ), //i
    .port_i_0_1 (keyAdd_port_state_out_8_0_1                ), //i
    .port_i_0_2 (keyAdd_port_state_out_8_0_2                ), //i
    .port_i_0_3 (keyAdd_port_state_out_8_0_3                ), //i
    .port_i_0_4 (keyAdd_port_state_out_8_0_4                ), //i
    .port_i_0_5 (keyAdd_port_state_out_8_0_5                ), //i
    .port_i_0_6 (keyAdd_port_state_out_8_0_6                ), //i
    .port_i_0_7 (keyAdd_port_state_out_8_0_7                ), //i
    .port_i_1_0 (keyAdd_port_state_out_8_1_0                ), //i
    .port_i_1_1 (keyAdd_port_state_out_8_1_1                ), //i
    .port_i_1_2 (keyAdd_port_state_out_8_1_2                ), //i
    .port_i_1_3 (keyAdd_port_state_out_8_1_3                ), //i
    .port_i_1_4 (keyAdd_port_state_out_8_1_4                ), //i
    .port_i_1_5 (keyAdd_port_state_out_8_1_5                ), //i
    .port_i_1_6 (keyAdd_port_state_out_8_1_6                ), //i
    .port_i_1_7 (keyAdd_port_state_out_8_1_7                ), //i
    .port_r_0   (port_rand_8_0                              ), //i
    .port_r_1   (port_rand_8_1                              ), //i
    .port_r_2   (port_rand_8_2                              ), //i
    .port_r_3   (port_rand_8_3                              ), //i
    .port_r_4   (port_rand_8_4                              ), //i
    .port_r_5   (port_rand_8_5                              ), //i
    .port_r_6   (port_rand_8_6                              ), //i
    .port_r_7   (port_rand_8_7                              ), //i
    .port_r_8   (port_rand_8_8                              ), //i
    .port_r_9   (port_rand_8_9                              ), //i
    .port_r_10  (port_rand_8_10                             ), //i
    .port_r_11  (port_rand_8_11                             ), //i
    .port_r_12  (port_rand_8_12                             ), //i
    .port_r_13  (port_rand_8_13                             ), //i
    .port_r_14  (port_rand_8_14                             ), //i
    .port_r_15  (port_rand_8_15                             ), //i
    .port_r_16  (port_rand_8_16                             ), //i
    .port_r_17  (port_rand_8_17                             ), //i
    .port_r_18  (port_rand_8_18                             ), //i
    .port_r_19  (port_rand_8_19                             ), //i
    .port_r_20  (port_rand_8_20                             ), //i
    .port_r_21  (port_rand_8_21                             ), //i
    .port_r_22  (port_rand_8_22                             ), //i
    .port_r_23  (port_rand_8_23                             ), //i
    .port_r_24  (port_rand_8_24                             ), //i
    .port_r_25  (port_rand_8_25                             ), //i
    .port_r_26  (port_rand_8_26                             ), //i
    .port_r_27  (port_rand_8_27                             ), //i
    .port_r_28  (port_rand_8_28                             ), //i
    .port_r_29  (port_rand_8_29                             ), //i
    .port_r_30  (port_rand_8_30                             ), //i
    .port_r_31  (port_rand_8_31                             ), //i
    .port_r_32  (port_rand_8_32                             ), //i
    .port_r_33  (port_rand_8_33                             ), //i
    .port_r_34  (port_rand_8_34                             ), //i
    .port_r_35  (port_rand_8_35                             ), //i
    .port_r_36  (port_rand_8_36                             ), //i
    .port_r_37  (port_rand_8_37                             ), //i
    .port_r_38  (port_rand_8_38                             ), //i
    .port_r_39  (port_rand_8_39                             ), //i
    .port_r_40  (port_rand_8_40                             ), //i
    .port_r_41  (port_rand_8_41                             ), //i
    .port_r_42  (port_rand_8_42                             ), //i
    .port_r_43  (port_rand_8_43                             ), //i
    .port_r_44  (port_rand_8_44                             ), //i
    .port_r_45  (port_rand_8_45                             ), //i
    .port_r_46  (port_rand_8_46                             ), //i
    .port_r_47  (port_rand_8_47                             ), //i
    .port_r_48  (port_rand_8_48                             ), //i
    .port_r_49  (port_rand_8_49                             ), //i
    .port_r_50  (port_rand_8_50                             ), //i
    .port_r_51  (port_rand_8_51                             ), //i
    .port_r_52  (port_rand_8_52                             ), //i
    .port_r_53  (port_rand_8_53                             ), //i
    .port_o_0_0 (sbox_AES_Canright_CMS_2shares_24_port_o_0_0), //o
    .port_o_0_1 (sbox_AES_Canright_CMS_2shares_24_port_o_0_1), //o
    .port_o_0_2 (sbox_AES_Canright_CMS_2shares_24_port_o_0_2), //o
    .port_o_0_3 (sbox_AES_Canright_CMS_2shares_24_port_o_0_3), //o
    .port_o_0_4 (sbox_AES_Canright_CMS_2shares_24_port_o_0_4), //o
    .port_o_0_5 (sbox_AES_Canright_CMS_2shares_24_port_o_0_5), //o
    .port_o_0_6 (sbox_AES_Canright_CMS_2shares_24_port_o_0_6), //o
    .port_o_0_7 (sbox_AES_Canright_CMS_2shares_24_port_o_0_7), //o
    .port_o_1_0 (sbox_AES_Canright_CMS_2shares_24_port_o_1_0), //o
    .port_o_1_1 (sbox_AES_Canright_CMS_2shares_24_port_o_1_1), //o
    .port_o_1_2 (sbox_AES_Canright_CMS_2shares_24_port_o_1_2), //o
    .port_o_1_3 (sbox_AES_Canright_CMS_2shares_24_port_o_1_3), //o
    .port_o_1_4 (sbox_AES_Canright_CMS_2shares_24_port_o_1_4), //o
    .port_o_1_5 (sbox_AES_Canright_CMS_2shares_24_port_o_1_5), //o
    .port_o_1_6 (sbox_AES_Canright_CMS_2shares_24_port_o_1_6), //o
    .port_o_1_7 (sbox_AES_Canright_CMS_2shares_24_port_o_1_7), //o
    .clk        (clk                                        ), //i
    .reset      (reset                                      )  //i
  );
  Sbox_AES_Canright_CMS_2shares sbox_AES_Canright_CMS_2shares_25 (
    .port_i_0_0 (keyAdd_port_state_out_9_0_0                ), //i
    .port_i_0_1 (keyAdd_port_state_out_9_0_1                ), //i
    .port_i_0_2 (keyAdd_port_state_out_9_0_2                ), //i
    .port_i_0_3 (keyAdd_port_state_out_9_0_3                ), //i
    .port_i_0_4 (keyAdd_port_state_out_9_0_4                ), //i
    .port_i_0_5 (keyAdd_port_state_out_9_0_5                ), //i
    .port_i_0_6 (keyAdd_port_state_out_9_0_6                ), //i
    .port_i_0_7 (keyAdd_port_state_out_9_0_7                ), //i
    .port_i_1_0 (keyAdd_port_state_out_9_1_0                ), //i
    .port_i_1_1 (keyAdd_port_state_out_9_1_1                ), //i
    .port_i_1_2 (keyAdd_port_state_out_9_1_2                ), //i
    .port_i_1_3 (keyAdd_port_state_out_9_1_3                ), //i
    .port_i_1_4 (keyAdd_port_state_out_9_1_4                ), //i
    .port_i_1_5 (keyAdd_port_state_out_9_1_5                ), //i
    .port_i_1_6 (keyAdd_port_state_out_9_1_6                ), //i
    .port_i_1_7 (keyAdd_port_state_out_9_1_7                ), //i
    .port_r_0   (port_rand_9_0                              ), //i
    .port_r_1   (port_rand_9_1                              ), //i
    .port_r_2   (port_rand_9_2                              ), //i
    .port_r_3   (port_rand_9_3                              ), //i
    .port_r_4   (port_rand_9_4                              ), //i
    .port_r_5   (port_rand_9_5                              ), //i
    .port_r_6   (port_rand_9_6                              ), //i
    .port_r_7   (port_rand_9_7                              ), //i
    .port_r_8   (port_rand_9_8                              ), //i
    .port_r_9   (port_rand_9_9                              ), //i
    .port_r_10  (port_rand_9_10                             ), //i
    .port_r_11  (port_rand_9_11                             ), //i
    .port_r_12  (port_rand_9_12                             ), //i
    .port_r_13  (port_rand_9_13                             ), //i
    .port_r_14  (port_rand_9_14                             ), //i
    .port_r_15  (port_rand_9_15                             ), //i
    .port_r_16  (port_rand_9_16                             ), //i
    .port_r_17  (port_rand_9_17                             ), //i
    .port_r_18  (port_rand_9_18                             ), //i
    .port_r_19  (port_rand_9_19                             ), //i
    .port_r_20  (port_rand_9_20                             ), //i
    .port_r_21  (port_rand_9_21                             ), //i
    .port_r_22  (port_rand_9_22                             ), //i
    .port_r_23  (port_rand_9_23                             ), //i
    .port_r_24  (port_rand_9_24                             ), //i
    .port_r_25  (port_rand_9_25                             ), //i
    .port_r_26  (port_rand_9_26                             ), //i
    .port_r_27  (port_rand_9_27                             ), //i
    .port_r_28  (port_rand_9_28                             ), //i
    .port_r_29  (port_rand_9_29                             ), //i
    .port_r_30  (port_rand_9_30                             ), //i
    .port_r_31  (port_rand_9_31                             ), //i
    .port_r_32  (port_rand_9_32                             ), //i
    .port_r_33  (port_rand_9_33                             ), //i
    .port_r_34  (port_rand_9_34                             ), //i
    .port_r_35  (port_rand_9_35                             ), //i
    .port_r_36  (port_rand_9_36                             ), //i
    .port_r_37  (port_rand_9_37                             ), //i
    .port_r_38  (port_rand_9_38                             ), //i
    .port_r_39  (port_rand_9_39                             ), //i
    .port_r_40  (port_rand_9_40                             ), //i
    .port_r_41  (port_rand_9_41                             ), //i
    .port_r_42  (port_rand_9_42                             ), //i
    .port_r_43  (port_rand_9_43                             ), //i
    .port_r_44  (port_rand_9_44                             ), //i
    .port_r_45  (port_rand_9_45                             ), //i
    .port_r_46  (port_rand_9_46                             ), //i
    .port_r_47  (port_rand_9_47                             ), //i
    .port_r_48  (port_rand_9_48                             ), //i
    .port_r_49  (port_rand_9_49                             ), //i
    .port_r_50  (port_rand_9_50                             ), //i
    .port_r_51  (port_rand_9_51                             ), //i
    .port_r_52  (port_rand_9_52                             ), //i
    .port_r_53  (port_rand_9_53                             ), //i
    .port_o_0_0 (sbox_AES_Canright_CMS_2shares_25_port_o_0_0), //o
    .port_o_0_1 (sbox_AES_Canright_CMS_2shares_25_port_o_0_1), //o
    .port_o_0_2 (sbox_AES_Canright_CMS_2shares_25_port_o_0_2), //o
    .port_o_0_3 (sbox_AES_Canright_CMS_2shares_25_port_o_0_3), //o
    .port_o_0_4 (sbox_AES_Canright_CMS_2shares_25_port_o_0_4), //o
    .port_o_0_5 (sbox_AES_Canright_CMS_2shares_25_port_o_0_5), //o
    .port_o_0_6 (sbox_AES_Canright_CMS_2shares_25_port_o_0_6), //o
    .port_o_0_7 (sbox_AES_Canright_CMS_2shares_25_port_o_0_7), //o
    .port_o_1_0 (sbox_AES_Canright_CMS_2shares_25_port_o_1_0), //o
    .port_o_1_1 (sbox_AES_Canright_CMS_2shares_25_port_o_1_1), //o
    .port_o_1_2 (sbox_AES_Canright_CMS_2shares_25_port_o_1_2), //o
    .port_o_1_3 (sbox_AES_Canright_CMS_2shares_25_port_o_1_3), //o
    .port_o_1_4 (sbox_AES_Canright_CMS_2shares_25_port_o_1_4), //o
    .port_o_1_5 (sbox_AES_Canright_CMS_2shares_25_port_o_1_5), //o
    .port_o_1_6 (sbox_AES_Canright_CMS_2shares_25_port_o_1_6), //o
    .port_o_1_7 (sbox_AES_Canright_CMS_2shares_25_port_o_1_7), //o
    .clk        (clk                                        ), //i
    .reset      (reset                                      )  //i
  );
  Sbox_AES_Canright_CMS_2shares sbox_AES_Canright_CMS_2shares_26 (
    .port_i_0_0 (keyAdd_port_state_out_10_0_0               ), //i
    .port_i_0_1 (keyAdd_port_state_out_10_0_1               ), //i
    .port_i_0_2 (keyAdd_port_state_out_10_0_2               ), //i
    .port_i_0_3 (keyAdd_port_state_out_10_0_3               ), //i
    .port_i_0_4 (keyAdd_port_state_out_10_0_4               ), //i
    .port_i_0_5 (keyAdd_port_state_out_10_0_5               ), //i
    .port_i_0_6 (keyAdd_port_state_out_10_0_6               ), //i
    .port_i_0_7 (keyAdd_port_state_out_10_0_7               ), //i
    .port_i_1_0 (keyAdd_port_state_out_10_1_0               ), //i
    .port_i_1_1 (keyAdd_port_state_out_10_1_1               ), //i
    .port_i_1_2 (keyAdd_port_state_out_10_1_2               ), //i
    .port_i_1_3 (keyAdd_port_state_out_10_1_3               ), //i
    .port_i_1_4 (keyAdd_port_state_out_10_1_4               ), //i
    .port_i_1_5 (keyAdd_port_state_out_10_1_5               ), //i
    .port_i_1_6 (keyAdd_port_state_out_10_1_6               ), //i
    .port_i_1_7 (keyAdd_port_state_out_10_1_7               ), //i
    .port_r_0   (port_rand_10_0                             ), //i
    .port_r_1   (port_rand_10_1                             ), //i
    .port_r_2   (port_rand_10_2                             ), //i
    .port_r_3   (port_rand_10_3                             ), //i
    .port_r_4   (port_rand_10_4                             ), //i
    .port_r_5   (port_rand_10_5                             ), //i
    .port_r_6   (port_rand_10_6                             ), //i
    .port_r_7   (port_rand_10_7                             ), //i
    .port_r_8   (port_rand_10_8                             ), //i
    .port_r_9   (port_rand_10_9                             ), //i
    .port_r_10  (port_rand_10_10                            ), //i
    .port_r_11  (port_rand_10_11                            ), //i
    .port_r_12  (port_rand_10_12                            ), //i
    .port_r_13  (port_rand_10_13                            ), //i
    .port_r_14  (port_rand_10_14                            ), //i
    .port_r_15  (port_rand_10_15                            ), //i
    .port_r_16  (port_rand_10_16                            ), //i
    .port_r_17  (port_rand_10_17                            ), //i
    .port_r_18  (port_rand_10_18                            ), //i
    .port_r_19  (port_rand_10_19                            ), //i
    .port_r_20  (port_rand_10_20                            ), //i
    .port_r_21  (port_rand_10_21                            ), //i
    .port_r_22  (port_rand_10_22                            ), //i
    .port_r_23  (port_rand_10_23                            ), //i
    .port_r_24  (port_rand_10_24                            ), //i
    .port_r_25  (port_rand_10_25                            ), //i
    .port_r_26  (port_rand_10_26                            ), //i
    .port_r_27  (port_rand_10_27                            ), //i
    .port_r_28  (port_rand_10_28                            ), //i
    .port_r_29  (port_rand_10_29                            ), //i
    .port_r_30  (port_rand_10_30                            ), //i
    .port_r_31  (port_rand_10_31                            ), //i
    .port_r_32  (port_rand_10_32                            ), //i
    .port_r_33  (port_rand_10_33                            ), //i
    .port_r_34  (port_rand_10_34                            ), //i
    .port_r_35  (port_rand_10_35                            ), //i
    .port_r_36  (port_rand_10_36                            ), //i
    .port_r_37  (port_rand_10_37                            ), //i
    .port_r_38  (port_rand_10_38                            ), //i
    .port_r_39  (port_rand_10_39                            ), //i
    .port_r_40  (port_rand_10_40                            ), //i
    .port_r_41  (port_rand_10_41                            ), //i
    .port_r_42  (port_rand_10_42                            ), //i
    .port_r_43  (port_rand_10_43                            ), //i
    .port_r_44  (port_rand_10_44                            ), //i
    .port_r_45  (port_rand_10_45                            ), //i
    .port_r_46  (port_rand_10_46                            ), //i
    .port_r_47  (port_rand_10_47                            ), //i
    .port_r_48  (port_rand_10_48                            ), //i
    .port_r_49  (port_rand_10_49                            ), //i
    .port_r_50  (port_rand_10_50                            ), //i
    .port_r_51  (port_rand_10_51                            ), //i
    .port_r_52  (port_rand_10_52                            ), //i
    .port_r_53  (port_rand_10_53                            ), //i
    .port_o_0_0 (sbox_AES_Canright_CMS_2shares_26_port_o_0_0), //o
    .port_o_0_1 (sbox_AES_Canright_CMS_2shares_26_port_o_0_1), //o
    .port_o_0_2 (sbox_AES_Canright_CMS_2shares_26_port_o_0_2), //o
    .port_o_0_3 (sbox_AES_Canright_CMS_2shares_26_port_o_0_3), //o
    .port_o_0_4 (sbox_AES_Canright_CMS_2shares_26_port_o_0_4), //o
    .port_o_0_5 (sbox_AES_Canright_CMS_2shares_26_port_o_0_5), //o
    .port_o_0_6 (sbox_AES_Canright_CMS_2shares_26_port_o_0_6), //o
    .port_o_0_7 (sbox_AES_Canright_CMS_2shares_26_port_o_0_7), //o
    .port_o_1_0 (sbox_AES_Canright_CMS_2shares_26_port_o_1_0), //o
    .port_o_1_1 (sbox_AES_Canright_CMS_2shares_26_port_o_1_1), //o
    .port_o_1_2 (sbox_AES_Canright_CMS_2shares_26_port_o_1_2), //o
    .port_o_1_3 (sbox_AES_Canright_CMS_2shares_26_port_o_1_3), //o
    .port_o_1_4 (sbox_AES_Canright_CMS_2shares_26_port_o_1_4), //o
    .port_o_1_5 (sbox_AES_Canright_CMS_2shares_26_port_o_1_5), //o
    .port_o_1_6 (sbox_AES_Canright_CMS_2shares_26_port_o_1_6), //o
    .port_o_1_7 (sbox_AES_Canright_CMS_2shares_26_port_o_1_7), //o
    .clk        (clk                                        ), //i
    .reset      (reset                                      )  //i
  );
  Sbox_AES_Canright_CMS_2shares sbox_AES_Canright_CMS_2shares_27 (
    .port_i_0_0 (keyAdd_port_state_out_11_0_0               ), //i
    .port_i_0_1 (keyAdd_port_state_out_11_0_1               ), //i
    .port_i_0_2 (keyAdd_port_state_out_11_0_2               ), //i
    .port_i_0_3 (keyAdd_port_state_out_11_0_3               ), //i
    .port_i_0_4 (keyAdd_port_state_out_11_0_4               ), //i
    .port_i_0_5 (keyAdd_port_state_out_11_0_5               ), //i
    .port_i_0_6 (keyAdd_port_state_out_11_0_6               ), //i
    .port_i_0_7 (keyAdd_port_state_out_11_0_7               ), //i
    .port_i_1_0 (keyAdd_port_state_out_11_1_0               ), //i
    .port_i_1_1 (keyAdd_port_state_out_11_1_1               ), //i
    .port_i_1_2 (keyAdd_port_state_out_11_1_2               ), //i
    .port_i_1_3 (keyAdd_port_state_out_11_1_3               ), //i
    .port_i_1_4 (keyAdd_port_state_out_11_1_4               ), //i
    .port_i_1_5 (keyAdd_port_state_out_11_1_5               ), //i
    .port_i_1_6 (keyAdd_port_state_out_11_1_6               ), //i
    .port_i_1_7 (keyAdd_port_state_out_11_1_7               ), //i
    .port_r_0   (port_rand_11_0                             ), //i
    .port_r_1   (port_rand_11_1                             ), //i
    .port_r_2   (port_rand_11_2                             ), //i
    .port_r_3   (port_rand_11_3                             ), //i
    .port_r_4   (port_rand_11_4                             ), //i
    .port_r_5   (port_rand_11_5                             ), //i
    .port_r_6   (port_rand_11_6                             ), //i
    .port_r_7   (port_rand_11_7                             ), //i
    .port_r_8   (port_rand_11_8                             ), //i
    .port_r_9   (port_rand_11_9                             ), //i
    .port_r_10  (port_rand_11_10                            ), //i
    .port_r_11  (port_rand_11_11                            ), //i
    .port_r_12  (port_rand_11_12                            ), //i
    .port_r_13  (port_rand_11_13                            ), //i
    .port_r_14  (port_rand_11_14                            ), //i
    .port_r_15  (port_rand_11_15                            ), //i
    .port_r_16  (port_rand_11_16                            ), //i
    .port_r_17  (port_rand_11_17                            ), //i
    .port_r_18  (port_rand_11_18                            ), //i
    .port_r_19  (port_rand_11_19                            ), //i
    .port_r_20  (port_rand_11_20                            ), //i
    .port_r_21  (port_rand_11_21                            ), //i
    .port_r_22  (port_rand_11_22                            ), //i
    .port_r_23  (port_rand_11_23                            ), //i
    .port_r_24  (port_rand_11_24                            ), //i
    .port_r_25  (port_rand_11_25                            ), //i
    .port_r_26  (port_rand_11_26                            ), //i
    .port_r_27  (port_rand_11_27                            ), //i
    .port_r_28  (port_rand_11_28                            ), //i
    .port_r_29  (port_rand_11_29                            ), //i
    .port_r_30  (port_rand_11_30                            ), //i
    .port_r_31  (port_rand_11_31                            ), //i
    .port_r_32  (port_rand_11_32                            ), //i
    .port_r_33  (port_rand_11_33                            ), //i
    .port_r_34  (port_rand_11_34                            ), //i
    .port_r_35  (port_rand_11_35                            ), //i
    .port_r_36  (port_rand_11_36                            ), //i
    .port_r_37  (port_rand_11_37                            ), //i
    .port_r_38  (port_rand_11_38                            ), //i
    .port_r_39  (port_rand_11_39                            ), //i
    .port_r_40  (port_rand_11_40                            ), //i
    .port_r_41  (port_rand_11_41                            ), //i
    .port_r_42  (port_rand_11_42                            ), //i
    .port_r_43  (port_rand_11_43                            ), //i
    .port_r_44  (port_rand_11_44                            ), //i
    .port_r_45  (port_rand_11_45                            ), //i
    .port_r_46  (port_rand_11_46                            ), //i
    .port_r_47  (port_rand_11_47                            ), //i
    .port_r_48  (port_rand_11_48                            ), //i
    .port_r_49  (port_rand_11_49                            ), //i
    .port_r_50  (port_rand_11_50                            ), //i
    .port_r_51  (port_rand_11_51                            ), //i
    .port_r_52  (port_rand_11_52                            ), //i
    .port_r_53  (port_rand_11_53                            ), //i
    .port_o_0_0 (sbox_AES_Canright_CMS_2shares_27_port_o_0_0), //o
    .port_o_0_1 (sbox_AES_Canright_CMS_2shares_27_port_o_0_1), //o
    .port_o_0_2 (sbox_AES_Canright_CMS_2shares_27_port_o_0_2), //o
    .port_o_0_3 (sbox_AES_Canright_CMS_2shares_27_port_o_0_3), //o
    .port_o_0_4 (sbox_AES_Canright_CMS_2shares_27_port_o_0_4), //o
    .port_o_0_5 (sbox_AES_Canright_CMS_2shares_27_port_o_0_5), //o
    .port_o_0_6 (sbox_AES_Canright_CMS_2shares_27_port_o_0_6), //o
    .port_o_0_7 (sbox_AES_Canright_CMS_2shares_27_port_o_0_7), //o
    .port_o_1_0 (sbox_AES_Canright_CMS_2shares_27_port_o_1_0), //o
    .port_o_1_1 (sbox_AES_Canright_CMS_2shares_27_port_o_1_1), //o
    .port_o_1_2 (sbox_AES_Canright_CMS_2shares_27_port_o_1_2), //o
    .port_o_1_3 (sbox_AES_Canright_CMS_2shares_27_port_o_1_3), //o
    .port_o_1_4 (sbox_AES_Canright_CMS_2shares_27_port_o_1_4), //o
    .port_o_1_5 (sbox_AES_Canright_CMS_2shares_27_port_o_1_5), //o
    .port_o_1_6 (sbox_AES_Canright_CMS_2shares_27_port_o_1_6), //o
    .port_o_1_7 (sbox_AES_Canright_CMS_2shares_27_port_o_1_7), //o
    .clk        (clk                                        ), //i
    .reset      (reset                                      )  //i
  );
  Sbox_AES_Canright_CMS_2shares sbox_AES_Canright_CMS_2shares_28 (
    .port_i_0_0 (keyAdd_port_state_out_12_0_0               ), //i
    .port_i_0_1 (keyAdd_port_state_out_12_0_1               ), //i
    .port_i_0_2 (keyAdd_port_state_out_12_0_2               ), //i
    .port_i_0_3 (keyAdd_port_state_out_12_0_3               ), //i
    .port_i_0_4 (keyAdd_port_state_out_12_0_4               ), //i
    .port_i_0_5 (keyAdd_port_state_out_12_0_5               ), //i
    .port_i_0_6 (keyAdd_port_state_out_12_0_6               ), //i
    .port_i_0_7 (keyAdd_port_state_out_12_0_7               ), //i
    .port_i_1_0 (keyAdd_port_state_out_12_1_0               ), //i
    .port_i_1_1 (keyAdd_port_state_out_12_1_1               ), //i
    .port_i_1_2 (keyAdd_port_state_out_12_1_2               ), //i
    .port_i_1_3 (keyAdd_port_state_out_12_1_3               ), //i
    .port_i_1_4 (keyAdd_port_state_out_12_1_4               ), //i
    .port_i_1_5 (keyAdd_port_state_out_12_1_5               ), //i
    .port_i_1_6 (keyAdd_port_state_out_12_1_6               ), //i
    .port_i_1_7 (keyAdd_port_state_out_12_1_7               ), //i
    .port_r_0   (port_rand_12_0                             ), //i
    .port_r_1   (port_rand_12_1                             ), //i
    .port_r_2   (port_rand_12_2                             ), //i
    .port_r_3   (port_rand_12_3                             ), //i
    .port_r_4   (port_rand_12_4                             ), //i
    .port_r_5   (port_rand_12_5                             ), //i
    .port_r_6   (port_rand_12_6                             ), //i
    .port_r_7   (port_rand_12_7                             ), //i
    .port_r_8   (port_rand_12_8                             ), //i
    .port_r_9   (port_rand_12_9                             ), //i
    .port_r_10  (port_rand_12_10                            ), //i
    .port_r_11  (port_rand_12_11                            ), //i
    .port_r_12  (port_rand_12_12                            ), //i
    .port_r_13  (port_rand_12_13                            ), //i
    .port_r_14  (port_rand_12_14                            ), //i
    .port_r_15  (port_rand_12_15                            ), //i
    .port_r_16  (port_rand_12_16                            ), //i
    .port_r_17  (port_rand_12_17                            ), //i
    .port_r_18  (port_rand_12_18                            ), //i
    .port_r_19  (port_rand_12_19                            ), //i
    .port_r_20  (port_rand_12_20                            ), //i
    .port_r_21  (port_rand_12_21                            ), //i
    .port_r_22  (port_rand_12_22                            ), //i
    .port_r_23  (port_rand_12_23                            ), //i
    .port_r_24  (port_rand_12_24                            ), //i
    .port_r_25  (port_rand_12_25                            ), //i
    .port_r_26  (port_rand_12_26                            ), //i
    .port_r_27  (port_rand_12_27                            ), //i
    .port_r_28  (port_rand_12_28                            ), //i
    .port_r_29  (port_rand_12_29                            ), //i
    .port_r_30  (port_rand_12_30                            ), //i
    .port_r_31  (port_rand_12_31                            ), //i
    .port_r_32  (port_rand_12_32                            ), //i
    .port_r_33  (port_rand_12_33                            ), //i
    .port_r_34  (port_rand_12_34                            ), //i
    .port_r_35  (port_rand_12_35                            ), //i
    .port_r_36  (port_rand_12_36                            ), //i
    .port_r_37  (port_rand_12_37                            ), //i
    .port_r_38  (port_rand_12_38                            ), //i
    .port_r_39  (port_rand_12_39                            ), //i
    .port_r_40  (port_rand_12_40                            ), //i
    .port_r_41  (port_rand_12_41                            ), //i
    .port_r_42  (port_rand_12_42                            ), //i
    .port_r_43  (port_rand_12_43                            ), //i
    .port_r_44  (port_rand_12_44                            ), //i
    .port_r_45  (port_rand_12_45                            ), //i
    .port_r_46  (port_rand_12_46                            ), //i
    .port_r_47  (port_rand_12_47                            ), //i
    .port_r_48  (port_rand_12_48                            ), //i
    .port_r_49  (port_rand_12_49                            ), //i
    .port_r_50  (port_rand_12_50                            ), //i
    .port_r_51  (port_rand_12_51                            ), //i
    .port_r_52  (port_rand_12_52                            ), //i
    .port_r_53  (port_rand_12_53                            ), //i
    .port_o_0_0 (sbox_AES_Canright_CMS_2shares_28_port_o_0_0), //o
    .port_o_0_1 (sbox_AES_Canright_CMS_2shares_28_port_o_0_1), //o
    .port_o_0_2 (sbox_AES_Canright_CMS_2shares_28_port_o_0_2), //o
    .port_o_0_3 (sbox_AES_Canright_CMS_2shares_28_port_o_0_3), //o
    .port_o_0_4 (sbox_AES_Canright_CMS_2shares_28_port_o_0_4), //o
    .port_o_0_5 (sbox_AES_Canright_CMS_2shares_28_port_o_0_5), //o
    .port_o_0_6 (sbox_AES_Canright_CMS_2shares_28_port_o_0_6), //o
    .port_o_0_7 (sbox_AES_Canright_CMS_2shares_28_port_o_0_7), //o
    .port_o_1_0 (sbox_AES_Canright_CMS_2shares_28_port_o_1_0), //o
    .port_o_1_1 (sbox_AES_Canright_CMS_2shares_28_port_o_1_1), //o
    .port_o_1_2 (sbox_AES_Canright_CMS_2shares_28_port_o_1_2), //o
    .port_o_1_3 (sbox_AES_Canright_CMS_2shares_28_port_o_1_3), //o
    .port_o_1_4 (sbox_AES_Canright_CMS_2shares_28_port_o_1_4), //o
    .port_o_1_5 (sbox_AES_Canright_CMS_2shares_28_port_o_1_5), //o
    .port_o_1_6 (sbox_AES_Canright_CMS_2shares_28_port_o_1_6), //o
    .port_o_1_7 (sbox_AES_Canright_CMS_2shares_28_port_o_1_7), //o
    .clk        (clk                                        ), //i
    .reset      (reset                                      )  //i
  );
  Sbox_AES_Canright_CMS_2shares sbox_AES_Canright_CMS_2shares_29 (
    .port_i_0_0 (keyAdd_port_state_out_13_0_0               ), //i
    .port_i_0_1 (keyAdd_port_state_out_13_0_1               ), //i
    .port_i_0_2 (keyAdd_port_state_out_13_0_2               ), //i
    .port_i_0_3 (keyAdd_port_state_out_13_0_3               ), //i
    .port_i_0_4 (keyAdd_port_state_out_13_0_4               ), //i
    .port_i_0_5 (keyAdd_port_state_out_13_0_5               ), //i
    .port_i_0_6 (keyAdd_port_state_out_13_0_6               ), //i
    .port_i_0_7 (keyAdd_port_state_out_13_0_7               ), //i
    .port_i_1_0 (keyAdd_port_state_out_13_1_0               ), //i
    .port_i_1_1 (keyAdd_port_state_out_13_1_1               ), //i
    .port_i_1_2 (keyAdd_port_state_out_13_1_2               ), //i
    .port_i_1_3 (keyAdd_port_state_out_13_1_3               ), //i
    .port_i_1_4 (keyAdd_port_state_out_13_1_4               ), //i
    .port_i_1_5 (keyAdd_port_state_out_13_1_5               ), //i
    .port_i_1_6 (keyAdd_port_state_out_13_1_6               ), //i
    .port_i_1_7 (keyAdd_port_state_out_13_1_7               ), //i
    .port_r_0   (port_rand_13_0                             ), //i
    .port_r_1   (port_rand_13_1                             ), //i
    .port_r_2   (port_rand_13_2                             ), //i
    .port_r_3   (port_rand_13_3                             ), //i
    .port_r_4   (port_rand_13_4                             ), //i
    .port_r_5   (port_rand_13_5                             ), //i
    .port_r_6   (port_rand_13_6                             ), //i
    .port_r_7   (port_rand_13_7                             ), //i
    .port_r_8   (port_rand_13_8                             ), //i
    .port_r_9   (port_rand_13_9                             ), //i
    .port_r_10  (port_rand_13_10                            ), //i
    .port_r_11  (port_rand_13_11                            ), //i
    .port_r_12  (port_rand_13_12                            ), //i
    .port_r_13  (port_rand_13_13                            ), //i
    .port_r_14  (port_rand_13_14                            ), //i
    .port_r_15  (port_rand_13_15                            ), //i
    .port_r_16  (port_rand_13_16                            ), //i
    .port_r_17  (port_rand_13_17                            ), //i
    .port_r_18  (port_rand_13_18                            ), //i
    .port_r_19  (port_rand_13_19                            ), //i
    .port_r_20  (port_rand_13_20                            ), //i
    .port_r_21  (port_rand_13_21                            ), //i
    .port_r_22  (port_rand_13_22                            ), //i
    .port_r_23  (port_rand_13_23                            ), //i
    .port_r_24  (port_rand_13_24                            ), //i
    .port_r_25  (port_rand_13_25                            ), //i
    .port_r_26  (port_rand_13_26                            ), //i
    .port_r_27  (port_rand_13_27                            ), //i
    .port_r_28  (port_rand_13_28                            ), //i
    .port_r_29  (port_rand_13_29                            ), //i
    .port_r_30  (port_rand_13_30                            ), //i
    .port_r_31  (port_rand_13_31                            ), //i
    .port_r_32  (port_rand_13_32                            ), //i
    .port_r_33  (port_rand_13_33                            ), //i
    .port_r_34  (port_rand_13_34                            ), //i
    .port_r_35  (port_rand_13_35                            ), //i
    .port_r_36  (port_rand_13_36                            ), //i
    .port_r_37  (port_rand_13_37                            ), //i
    .port_r_38  (port_rand_13_38                            ), //i
    .port_r_39  (port_rand_13_39                            ), //i
    .port_r_40  (port_rand_13_40                            ), //i
    .port_r_41  (port_rand_13_41                            ), //i
    .port_r_42  (port_rand_13_42                            ), //i
    .port_r_43  (port_rand_13_43                            ), //i
    .port_r_44  (port_rand_13_44                            ), //i
    .port_r_45  (port_rand_13_45                            ), //i
    .port_r_46  (port_rand_13_46                            ), //i
    .port_r_47  (port_rand_13_47                            ), //i
    .port_r_48  (port_rand_13_48                            ), //i
    .port_r_49  (port_rand_13_49                            ), //i
    .port_r_50  (port_rand_13_50                            ), //i
    .port_r_51  (port_rand_13_51                            ), //i
    .port_r_52  (port_rand_13_52                            ), //i
    .port_r_53  (port_rand_13_53                            ), //i
    .port_o_0_0 (sbox_AES_Canright_CMS_2shares_29_port_o_0_0), //o
    .port_o_0_1 (sbox_AES_Canright_CMS_2shares_29_port_o_0_1), //o
    .port_o_0_2 (sbox_AES_Canright_CMS_2shares_29_port_o_0_2), //o
    .port_o_0_3 (sbox_AES_Canright_CMS_2shares_29_port_o_0_3), //o
    .port_o_0_4 (sbox_AES_Canright_CMS_2shares_29_port_o_0_4), //o
    .port_o_0_5 (sbox_AES_Canright_CMS_2shares_29_port_o_0_5), //o
    .port_o_0_6 (sbox_AES_Canright_CMS_2shares_29_port_o_0_6), //o
    .port_o_0_7 (sbox_AES_Canright_CMS_2shares_29_port_o_0_7), //o
    .port_o_1_0 (sbox_AES_Canright_CMS_2shares_29_port_o_1_0), //o
    .port_o_1_1 (sbox_AES_Canright_CMS_2shares_29_port_o_1_1), //o
    .port_o_1_2 (sbox_AES_Canright_CMS_2shares_29_port_o_1_2), //o
    .port_o_1_3 (sbox_AES_Canright_CMS_2shares_29_port_o_1_3), //o
    .port_o_1_4 (sbox_AES_Canright_CMS_2shares_29_port_o_1_4), //o
    .port_o_1_5 (sbox_AES_Canright_CMS_2shares_29_port_o_1_5), //o
    .port_o_1_6 (sbox_AES_Canright_CMS_2shares_29_port_o_1_6), //o
    .port_o_1_7 (sbox_AES_Canright_CMS_2shares_29_port_o_1_7), //o
    .clk        (clk                                        ), //i
    .reset      (reset                                      )  //i
  );
  Sbox_AES_Canright_CMS_2shares sbox_AES_Canright_CMS_2shares_30 (
    .port_i_0_0 (keyAdd_port_state_out_14_0_0               ), //i
    .port_i_0_1 (keyAdd_port_state_out_14_0_1               ), //i
    .port_i_0_2 (keyAdd_port_state_out_14_0_2               ), //i
    .port_i_0_3 (keyAdd_port_state_out_14_0_3               ), //i
    .port_i_0_4 (keyAdd_port_state_out_14_0_4               ), //i
    .port_i_0_5 (keyAdd_port_state_out_14_0_5               ), //i
    .port_i_0_6 (keyAdd_port_state_out_14_0_6               ), //i
    .port_i_0_7 (keyAdd_port_state_out_14_0_7               ), //i
    .port_i_1_0 (keyAdd_port_state_out_14_1_0               ), //i
    .port_i_1_1 (keyAdd_port_state_out_14_1_1               ), //i
    .port_i_1_2 (keyAdd_port_state_out_14_1_2               ), //i
    .port_i_1_3 (keyAdd_port_state_out_14_1_3               ), //i
    .port_i_1_4 (keyAdd_port_state_out_14_1_4               ), //i
    .port_i_1_5 (keyAdd_port_state_out_14_1_5               ), //i
    .port_i_1_6 (keyAdd_port_state_out_14_1_6               ), //i
    .port_i_1_7 (keyAdd_port_state_out_14_1_7               ), //i
    .port_r_0   (port_rand_14_0                             ), //i
    .port_r_1   (port_rand_14_1                             ), //i
    .port_r_2   (port_rand_14_2                             ), //i
    .port_r_3   (port_rand_14_3                             ), //i
    .port_r_4   (port_rand_14_4                             ), //i
    .port_r_5   (port_rand_14_5                             ), //i
    .port_r_6   (port_rand_14_6                             ), //i
    .port_r_7   (port_rand_14_7                             ), //i
    .port_r_8   (port_rand_14_8                             ), //i
    .port_r_9   (port_rand_14_9                             ), //i
    .port_r_10  (port_rand_14_10                            ), //i
    .port_r_11  (port_rand_14_11                            ), //i
    .port_r_12  (port_rand_14_12                            ), //i
    .port_r_13  (port_rand_14_13                            ), //i
    .port_r_14  (port_rand_14_14                            ), //i
    .port_r_15  (port_rand_14_15                            ), //i
    .port_r_16  (port_rand_14_16                            ), //i
    .port_r_17  (port_rand_14_17                            ), //i
    .port_r_18  (port_rand_14_18                            ), //i
    .port_r_19  (port_rand_14_19                            ), //i
    .port_r_20  (port_rand_14_20                            ), //i
    .port_r_21  (port_rand_14_21                            ), //i
    .port_r_22  (port_rand_14_22                            ), //i
    .port_r_23  (port_rand_14_23                            ), //i
    .port_r_24  (port_rand_14_24                            ), //i
    .port_r_25  (port_rand_14_25                            ), //i
    .port_r_26  (port_rand_14_26                            ), //i
    .port_r_27  (port_rand_14_27                            ), //i
    .port_r_28  (port_rand_14_28                            ), //i
    .port_r_29  (port_rand_14_29                            ), //i
    .port_r_30  (port_rand_14_30                            ), //i
    .port_r_31  (port_rand_14_31                            ), //i
    .port_r_32  (port_rand_14_32                            ), //i
    .port_r_33  (port_rand_14_33                            ), //i
    .port_r_34  (port_rand_14_34                            ), //i
    .port_r_35  (port_rand_14_35                            ), //i
    .port_r_36  (port_rand_14_36                            ), //i
    .port_r_37  (port_rand_14_37                            ), //i
    .port_r_38  (port_rand_14_38                            ), //i
    .port_r_39  (port_rand_14_39                            ), //i
    .port_r_40  (port_rand_14_40                            ), //i
    .port_r_41  (port_rand_14_41                            ), //i
    .port_r_42  (port_rand_14_42                            ), //i
    .port_r_43  (port_rand_14_43                            ), //i
    .port_r_44  (port_rand_14_44                            ), //i
    .port_r_45  (port_rand_14_45                            ), //i
    .port_r_46  (port_rand_14_46                            ), //i
    .port_r_47  (port_rand_14_47                            ), //i
    .port_r_48  (port_rand_14_48                            ), //i
    .port_r_49  (port_rand_14_49                            ), //i
    .port_r_50  (port_rand_14_50                            ), //i
    .port_r_51  (port_rand_14_51                            ), //i
    .port_r_52  (port_rand_14_52                            ), //i
    .port_r_53  (port_rand_14_53                            ), //i
    .port_o_0_0 (sbox_AES_Canright_CMS_2shares_30_port_o_0_0), //o
    .port_o_0_1 (sbox_AES_Canright_CMS_2shares_30_port_o_0_1), //o
    .port_o_0_2 (sbox_AES_Canright_CMS_2shares_30_port_o_0_2), //o
    .port_o_0_3 (sbox_AES_Canright_CMS_2shares_30_port_o_0_3), //o
    .port_o_0_4 (sbox_AES_Canright_CMS_2shares_30_port_o_0_4), //o
    .port_o_0_5 (sbox_AES_Canright_CMS_2shares_30_port_o_0_5), //o
    .port_o_0_6 (sbox_AES_Canright_CMS_2shares_30_port_o_0_6), //o
    .port_o_0_7 (sbox_AES_Canright_CMS_2shares_30_port_o_0_7), //o
    .port_o_1_0 (sbox_AES_Canright_CMS_2shares_30_port_o_1_0), //o
    .port_o_1_1 (sbox_AES_Canright_CMS_2shares_30_port_o_1_1), //o
    .port_o_1_2 (sbox_AES_Canright_CMS_2shares_30_port_o_1_2), //o
    .port_o_1_3 (sbox_AES_Canright_CMS_2shares_30_port_o_1_3), //o
    .port_o_1_4 (sbox_AES_Canright_CMS_2shares_30_port_o_1_4), //o
    .port_o_1_5 (sbox_AES_Canright_CMS_2shares_30_port_o_1_5), //o
    .port_o_1_6 (sbox_AES_Canright_CMS_2shares_30_port_o_1_6), //o
    .port_o_1_7 (sbox_AES_Canright_CMS_2shares_30_port_o_1_7), //o
    .clk        (clk                                        ), //i
    .reset      (reset                                      )  //i
  );
  Sbox_AES_Canright_CMS_2shares sbox_AES_Canright_CMS_2shares_31 (
    .port_i_0_0 (keyAdd_port_state_out_15_0_0               ), //i
    .port_i_0_1 (keyAdd_port_state_out_15_0_1               ), //i
    .port_i_0_2 (keyAdd_port_state_out_15_0_2               ), //i
    .port_i_0_3 (keyAdd_port_state_out_15_0_3               ), //i
    .port_i_0_4 (keyAdd_port_state_out_15_0_4               ), //i
    .port_i_0_5 (keyAdd_port_state_out_15_0_5               ), //i
    .port_i_0_6 (keyAdd_port_state_out_15_0_6               ), //i
    .port_i_0_7 (keyAdd_port_state_out_15_0_7               ), //i
    .port_i_1_0 (keyAdd_port_state_out_15_1_0               ), //i
    .port_i_1_1 (keyAdd_port_state_out_15_1_1               ), //i
    .port_i_1_2 (keyAdd_port_state_out_15_1_2               ), //i
    .port_i_1_3 (keyAdd_port_state_out_15_1_3               ), //i
    .port_i_1_4 (keyAdd_port_state_out_15_1_4               ), //i
    .port_i_1_5 (keyAdd_port_state_out_15_1_5               ), //i
    .port_i_1_6 (keyAdd_port_state_out_15_1_6               ), //i
    .port_i_1_7 (keyAdd_port_state_out_15_1_7               ), //i
    .port_r_0   (port_rand_15_0                             ), //i
    .port_r_1   (port_rand_15_1                             ), //i
    .port_r_2   (port_rand_15_2                             ), //i
    .port_r_3   (port_rand_15_3                             ), //i
    .port_r_4   (port_rand_15_4                             ), //i
    .port_r_5   (port_rand_15_5                             ), //i
    .port_r_6   (port_rand_15_6                             ), //i
    .port_r_7   (port_rand_15_7                             ), //i
    .port_r_8   (port_rand_15_8                             ), //i
    .port_r_9   (port_rand_15_9                             ), //i
    .port_r_10  (port_rand_15_10                            ), //i
    .port_r_11  (port_rand_15_11                            ), //i
    .port_r_12  (port_rand_15_12                            ), //i
    .port_r_13  (port_rand_15_13                            ), //i
    .port_r_14  (port_rand_15_14                            ), //i
    .port_r_15  (port_rand_15_15                            ), //i
    .port_r_16  (port_rand_15_16                            ), //i
    .port_r_17  (port_rand_15_17                            ), //i
    .port_r_18  (port_rand_15_18                            ), //i
    .port_r_19  (port_rand_15_19                            ), //i
    .port_r_20  (port_rand_15_20                            ), //i
    .port_r_21  (port_rand_15_21                            ), //i
    .port_r_22  (port_rand_15_22                            ), //i
    .port_r_23  (port_rand_15_23                            ), //i
    .port_r_24  (port_rand_15_24                            ), //i
    .port_r_25  (port_rand_15_25                            ), //i
    .port_r_26  (port_rand_15_26                            ), //i
    .port_r_27  (port_rand_15_27                            ), //i
    .port_r_28  (port_rand_15_28                            ), //i
    .port_r_29  (port_rand_15_29                            ), //i
    .port_r_30  (port_rand_15_30                            ), //i
    .port_r_31  (port_rand_15_31                            ), //i
    .port_r_32  (port_rand_15_32                            ), //i
    .port_r_33  (port_rand_15_33                            ), //i
    .port_r_34  (port_rand_15_34                            ), //i
    .port_r_35  (port_rand_15_35                            ), //i
    .port_r_36  (port_rand_15_36                            ), //i
    .port_r_37  (port_rand_15_37                            ), //i
    .port_r_38  (port_rand_15_38                            ), //i
    .port_r_39  (port_rand_15_39                            ), //i
    .port_r_40  (port_rand_15_40                            ), //i
    .port_r_41  (port_rand_15_41                            ), //i
    .port_r_42  (port_rand_15_42                            ), //i
    .port_r_43  (port_rand_15_43                            ), //i
    .port_r_44  (port_rand_15_44                            ), //i
    .port_r_45  (port_rand_15_45                            ), //i
    .port_r_46  (port_rand_15_46                            ), //i
    .port_r_47  (port_rand_15_47                            ), //i
    .port_r_48  (port_rand_15_48                            ), //i
    .port_r_49  (port_rand_15_49                            ), //i
    .port_r_50  (port_rand_15_50                            ), //i
    .port_r_51  (port_rand_15_51                            ), //i
    .port_r_52  (port_rand_15_52                            ), //i
    .port_r_53  (port_rand_15_53                            ), //i
    .port_o_0_0 (sbox_AES_Canright_CMS_2shares_31_port_o_0_0), //o
    .port_o_0_1 (sbox_AES_Canright_CMS_2shares_31_port_o_0_1), //o
    .port_o_0_2 (sbox_AES_Canright_CMS_2shares_31_port_o_0_2), //o
    .port_o_0_3 (sbox_AES_Canright_CMS_2shares_31_port_o_0_3), //o
    .port_o_0_4 (sbox_AES_Canright_CMS_2shares_31_port_o_0_4), //o
    .port_o_0_5 (sbox_AES_Canright_CMS_2shares_31_port_o_0_5), //o
    .port_o_0_6 (sbox_AES_Canright_CMS_2shares_31_port_o_0_6), //o
    .port_o_0_7 (sbox_AES_Canright_CMS_2shares_31_port_o_0_7), //o
    .port_o_1_0 (sbox_AES_Canright_CMS_2shares_31_port_o_1_0), //o
    .port_o_1_1 (sbox_AES_Canright_CMS_2shares_31_port_o_1_1), //o
    .port_o_1_2 (sbox_AES_Canright_CMS_2shares_31_port_o_1_2), //o
    .port_o_1_3 (sbox_AES_Canright_CMS_2shares_31_port_o_1_3), //o
    .port_o_1_4 (sbox_AES_Canright_CMS_2shares_31_port_o_1_4), //o
    .port_o_1_5 (sbox_AES_Canright_CMS_2shares_31_port_o_1_5), //o
    .port_o_1_6 (sbox_AES_Canright_CMS_2shares_31_port_o_1_6), //o
    .port_o_1_7 (sbox_AES_Canright_CMS_2shares_31_port_o_1_7), //o
    .clk        (clk                                        ), //i
    .reset      (reset                                      )  //i
  );
  AES_ShiftRows shiftRows (
    .port_state_in_0_0_0   (subBytes_out_0_0_0             ), //i
    .port_state_in_0_0_1   (subBytes_out_0_0_1             ), //i
    .port_state_in_0_0_2   (subBytes_out_0_0_2             ), //i
    .port_state_in_0_0_3   (subBytes_out_0_0_3             ), //i
    .port_state_in_0_0_4   (subBytes_out_0_0_4             ), //i
    .port_state_in_0_0_5   (subBytes_out_0_0_5             ), //i
    .port_state_in_0_0_6   (subBytes_out_0_0_6             ), //i
    .port_state_in_0_0_7   (subBytes_out_0_0_7             ), //i
    .port_state_in_0_1_0   (subBytes_out_0_1_0             ), //i
    .port_state_in_0_1_1   (subBytes_out_0_1_1             ), //i
    .port_state_in_0_1_2   (subBytes_out_0_1_2             ), //i
    .port_state_in_0_1_3   (subBytes_out_0_1_3             ), //i
    .port_state_in_0_1_4   (subBytes_out_0_1_4             ), //i
    .port_state_in_0_1_5   (subBytes_out_0_1_5             ), //i
    .port_state_in_0_1_6   (subBytes_out_0_1_6             ), //i
    .port_state_in_0_1_7   (subBytes_out_0_1_7             ), //i
    .port_state_in_1_0_0   (subBytes_out_1_0_0             ), //i
    .port_state_in_1_0_1   (subBytes_out_1_0_1             ), //i
    .port_state_in_1_0_2   (subBytes_out_1_0_2             ), //i
    .port_state_in_1_0_3   (subBytes_out_1_0_3             ), //i
    .port_state_in_1_0_4   (subBytes_out_1_0_4             ), //i
    .port_state_in_1_0_5   (subBytes_out_1_0_5             ), //i
    .port_state_in_1_0_6   (subBytes_out_1_0_6             ), //i
    .port_state_in_1_0_7   (subBytes_out_1_0_7             ), //i
    .port_state_in_1_1_0   (subBytes_out_1_1_0             ), //i
    .port_state_in_1_1_1   (subBytes_out_1_1_1             ), //i
    .port_state_in_1_1_2   (subBytes_out_1_1_2             ), //i
    .port_state_in_1_1_3   (subBytes_out_1_1_3             ), //i
    .port_state_in_1_1_4   (subBytes_out_1_1_4             ), //i
    .port_state_in_1_1_5   (subBytes_out_1_1_5             ), //i
    .port_state_in_1_1_6   (subBytes_out_1_1_6             ), //i
    .port_state_in_1_1_7   (subBytes_out_1_1_7             ), //i
    .port_state_in_2_0_0   (subBytes_out_2_0_0             ), //i
    .port_state_in_2_0_1   (subBytes_out_2_0_1             ), //i
    .port_state_in_2_0_2   (subBytes_out_2_0_2             ), //i
    .port_state_in_2_0_3   (subBytes_out_2_0_3             ), //i
    .port_state_in_2_0_4   (subBytes_out_2_0_4             ), //i
    .port_state_in_2_0_5   (subBytes_out_2_0_5             ), //i
    .port_state_in_2_0_6   (subBytes_out_2_0_6             ), //i
    .port_state_in_2_0_7   (subBytes_out_2_0_7             ), //i
    .port_state_in_2_1_0   (subBytes_out_2_1_0             ), //i
    .port_state_in_2_1_1   (subBytes_out_2_1_1             ), //i
    .port_state_in_2_1_2   (subBytes_out_2_1_2             ), //i
    .port_state_in_2_1_3   (subBytes_out_2_1_3             ), //i
    .port_state_in_2_1_4   (subBytes_out_2_1_4             ), //i
    .port_state_in_2_1_5   (subBytes_out_2_1_5             ), //i
    .port_state_in_2_1_6   (subBytes_out_2_1_6             ), //i
    .port_state_in_2_1_7   (subBytes_out_2_1_7             ), //i
    .port_state_in_3_0_0   (subBytes_out_3_0_0             ), //i
    .port_state_in_3_0_1   (subBytes_out_3_0_1             ), //i
    .port_state_in_3_0_2   (subBytes_out_3_0_2             ), //i
    .port_state_in_3_0_3   (subBytes_out_3_0_3             ), //i
    .port_state_in_3_0_4   (subBytes_out_3_0_4             ), //i
    .port_state_in_3_0_5   (subBytes_out_3_0_5             ), //i
    .port_state_in_3_0_6   (subBytes_out_3_0_6             ), //i
    .port_state_in_3_0_7   (subBytes_out_3_0_7             ), //i
    .port_state_in_3_1_0   (subBytes_out_3_1_0             ), //i
    .port_state_in_3_1_1   (subBytes_out_3_1_1             ), //i
    .port_state_in_3_1_2   (subBytes_out_3_1_2             ), //i
    .port_state_in_3_1_3   (subBytes_out_3_1_3             ), //i
    .port_state_in_3_1_4   (subBytes_out_3_1_4             ), //i
    .port_state_in_3_1_5   (subBytes_out_3_1_5             ), //i
    .port_state_in_3_1_6   (subBytes_out_3_1_6             ), //i
    .port_state_in_3_1_7   (subBytes_out_3_1_7             ), //i
    .port_state_in_4_0_0   (subBytes_out_4_0_0             ), //i
    .port_state_in_4_0_1   (subBytes_out_4_0_1             ), //i
    .port_state_in_4_0_2   (subBytes_out_4_0_2             ), //i
    .port_state_in_4_0_3   (subBytes_out_4_0_3             ), //i
    .port_state_in_4_0_4   (subBytes_out_4_0_4             ), //i
    .port_state_in_4_0_5   (subBytes_out_4_0_5             ), //i
    .port_state_in_4_0_6   (subBytes_out_4_0_6             ), //i
    .port_state_in_4_0_7   (subBytes_out_4_0_7             ), //i
    .port_state_in_4_1_0   (subBytes_out_4_1_0             ), //i
    .port_state_in_4_1_1   (subBytes_out_4_1_1             ), //i
    .port_state_in_4_1_2   (subBytes_out_4_1_2             ), //i
    .port_state_in_4_1_3   (subBytes_out_4_1_3             ), //i
    .port_state_in_4_1_4   (subBytes_out_4_1_4             ), //i
    .port_state_in_4_1_5   (subBytes_out_4_1_5             ), //i
    .port_state_in_4_1_6   (subBytes_out_4_1_6             ), //i
    .port_state_in_4_1_7   (subBytes_out_4_1_7             ), //i
    .port_state_in_5_0_0   (subBytes_out_5_0_0             ), //i
    .port_state_in_5_0_1   (subBytes_out_5_0_1             ), //i
    .port_state_in_5_0_2   (subBytes_out_5_0_2             ), //i
    .port_state_in_5_0_3   (subBytes_out_5_0_3             ), //i
    .port_state_in_5_0_4   (subBytes_out_5_0_4             ), //i
    .port_state_in_5_0_5   (subBytes_out_5_0_5             ), //i
    .port_state_in_5_0_6   (subBytes_out_5_0_6             ), //i
    .port_state_in_5_0_7   (subBytes_out_5_0_7             ), //i
    .port_state_in_5_1_0   (subBytes_out_5_1_0             ), //i
    .port_state_in_5_1_1   (subBytes_out_5_1_1             ), //i
    .port_state_in_5_1_2   (subBytes_out_5_1_2             ), //i
    .port_state_in_5_1_3   (subBytes_out_5_1_3             ), //i
    .port_state_in_5_1_4   (subBytes_out_5_1_4             ), //i
    .port_state_in_5_1_5   (subBytes_out_5_1_5             ), //i
    .port_state_in_5_1_6   (subBytes_out_5_1_6             ), //i
    .port_state_in_5_1_7   (subBytes_out_5_1_7             ), //i
    .port_state_in_6_0_0   (subBytes_out_6_0_0             ), //i
    .port_state_in_6_0_1   (subBytes_out_6_0_1             ), //i
    .port_state_in_6_0_2   (subBytes_out_6_0_2             ), //i
    .port_state_in_6_0_3   (subBytes_out_6_0_3             ), //i
    .port_state_in_6_0_4   (subBytes_out_6_0_4             ), //i
    .port_state_in_6_0_5   (subBytes_out_6_0_5             ), //i
    .port_state_in_6_0_6   (subBytes_out_6_0_6             ), //i
    .port_state_in_6_0_7   (subBytes_out_6_0_7             ), //i
    .port_state_in_6_1_0   (subBytes_out_6_1_0             ), //i
    .port_state_in_6_1_1   (subBytes_out_6_1_1             ), //i
    .port_state_in_6_1_2   (subBytes_out_6_1_2             ), //i
    .port_state_in_6_1_3   (subBytes_out_6_1_3             ), //i
    .port_state_in_6_1_4   (subBytes_out_6_1_4             ), //i
    .port_state_in_6_1_5   (subBytes_out_6_1_5             ), //i
    .port_state_in_6_1_6   (subBytes_out_6_1_6             ), //i
    .port_state_in_6_1_7   (subBytes_out_6_1_7             ), //i
    .port_state_in_7_0_0   (subBytes_out_7_0_0             ), //i
    .port_state_in_7_0_1   (subBytes_out_7_0_1             ), //i
    .port_state_in_7_0_2   (subBytes_out_7_0_2             ), //i
    .port_state_in_7_0_3   (subBytes_out_7_0_3             ), //i
    .port_state_in_7_0_4   (subBytes_out_7_0_4             ), //i
    .port_state_in_7_0_5   (subBytes_out_7_0_5             ), //i
    .port_state_in_7_0_6   (subBytes_out_7_0_6             ), //i
    .port_state_in_7_0_7   (subBytes_out_7_0_7             ), //i
    .port_state_in_7_1_0   (subBytes_out_7_1_0             ), //i
    .port_state_in_7_1_1   (subBytes_out_7_1_1             ), //i
    .port_state_in_7_1_2   (subBytes_out_7_1_2             ), //i
    .port_state_in_7_1_3   (subBytes_out_7_1_3             ), //i
    .port_state_in_7_1_4   (subBytes_out_7_1_4             ), //i
    .port_state_in_7_1_5   (subBytes_out_7_1_5             ), //i
    .port_state_in_7_1_6   (subBytes_out_7_1_6             ), //i
    .port_state_in_7_1_7   (subBytes_out_7_1_7             ), //i
    .port_state_in_8_0_0   (subBytes_out_8_0_0             ), //i
    .port_state_in_8_0_1   (subBytes_out_8_0_1             ), //i
    .port_state_in_8_0_2   (subBytes_out_8_0_2             ), //i
    .port_state_in_8_0_3   (subBytes_out_8_0_3             ), //i
    .port_state_in_8_0_4   (subBytes_out_8_0_4             ), //i
    .port_state_in_8_0_5   (subBytes_out_8_0_5             ), //i
    .port_state_in_8_0_6   (subBytes_out_8_0_6             ), //i
    .port_state_in_8_0_7   (subBytes_out_8_0_7             ), //i
    .port_state_in_8_1_0   (subBytes_out_8_1_0             ), //i
    .port_state_in_8_1_1   (subBytes_out_8_1_1             ), //i
    .port_state_in_8_1_2   (subBytes_out_8_1_2             ), //i
    .port_state_in_8_1_3   (subBytes_out_8_1_3             ), //i
    .port_state_in_8_1_4   (subBytes_out_8_1_4             ), //i
    .port_state_in_8_1_5   (subBytes_out_8_1_5             ), //i
    .port_state_in_8_1_6   (subBytes_out_8_1_6             ), //i
    .port_state_in_8_1_7   (subBytes_out_8_1_7             ), //i
    .port_state_in_9_0_0   (subBytes_out_9_0_0             ), //i
    .port_state_in_9_0_1   (subBytes_out_9_0_1             ), //i
    .port_state_in_9_0_2   (subBytes_out_9_0_2             ), //i
    .port_state_in_9_0_3   (subBytes_out_9_0_3             ), //i
    .port_state_in_9_0_4   (subBytes_out_9_0_4             ), //i
    .port_state_in_9_0_5   (subBytes_out_9_0_5             ), //i
    .port_state_in_9_0_6   (subBytes_out_9_0_6             ), //i
    .port_state_in_9_0_7   (subBytes_out_9_0_7             ), //i
    .port_state_in_9_1_0   (subBytes_out_9_1_0             ), //i
    .port_state_in_9_1_1   (subBytes_out_9_1_1             ), //i
    .port_state_in_9_1_2   (subBytes_out_9_1_2             ), //i
    .port_state_in_9_1_3   (subBytes_out_9_1_3             ), //i
    .port_state_in_9_1_4   (subBytes_out_9_1_4             ), //i
    .port_state_in_9_1_5   (subBytes_out_9_1_5             ), //i
    .port_state_in_9_1_6   (subBytes_out_9_1_6             ), //i
    .port_state_in_9_1_7   (subBytes_out_9_1_7             ), //i
    .port_state_in_10_0_0  (subBytes_out_10_0_0            ), //i
    .port_state_in_10_0_1  (subBytes_out_10_0_1            ), //i
    .port_state_in_10_0_2  (subBytes_out_10_0_2            ), //i
    .port_state_in_10_0_3  (subBytes_out_10_0_3            ), //i
    .port_state_in_10_0_4  (subBytes_out_10_0_4            ), //i
    .port_state_in_10_0_5  (subBytes_out_10_0_5            ), //i
    .port_state_in_10_0_6  (subBytes_out_10_0_6            ), //i
    .port_state_in_10_0_7  (subBytes_out_10_0_7            ), //i
    .port_state_in_10_1_0  (subBytes_out_10_1_0            ), //i
    .port_state_in_10_1_1  (subBytes_out_10_1_1            ), //i
    .port_state_in_10_1_2  (subBytes_out_10_1_2            ), //i
    .port_state_in_10_1_3  (subBytes_out_10_1_3            ), //i
    .port_state_in_10_1_4  (subBytes_out_10_1_4            ), //i
    .port_state_in_10_1_5  (subBytes_out_10_1_5            ), //i
    .port_state_in_10_1_6  (subBytes_out_10_1_6            ), //i
    .port_state_in_10_1_7  (subBytes_out_10_1_7            ), //i
    .port_state_in_11_0_0  (subBytes_out_11_0_0            ), //i
    .port_state_in_11_0_1  (subBytes_out_11_0_1            ), //i
    .port_state_in_11_0_2  (subBytes_out_11_0_2            ), //i
    .port_state_in_11_0_3  (subBytes_out_11_0_3            ), //i
    .port_state_in_11_0_4  (subBytes_out_11_0_4            ), //i
    .port_state_in_11_0_5  (subBytes_out_11_0_5            ), //i
    .port_state_in_11_0_6  (subBytes_out_11_0_6            ), //i
    .port_state_in_11_0_7  (subBytes_out_11_0_7            ), //i
    .port_state_in_11_1_0  (subBytes_out_11_1_0            ), //i
    .port_state_in_11_1_1  (subBytes_out_11_1_1            ), //i
    .port_state_in_11_1_2  (subBytes_out_11_1_2            ), //i
    .port_state_in_11_1_3  (subBytes_out_11_1_3            ), //i
    .port_state_in_11_1_4  (subBytes_out_11_1_4            ), //i
    .port_state_in_11_1_5  (subBytes_out_11_1_5            ), //i
    .port_state_in_11_1_6  (subBytes_out_11_1_6            ), //i
    .port_state_in_11_1_7  (subBytes_out_11_1_7            ), //i
    .port_state_in_12_0_0  (subBytes_out_12_0_0            ), //i
    .port_state_in_12_0_1  (subBytes_out_12_0_1            ), //i
    .port_state_in_12_0_2  (subBytes_out_12_0_2            ), //i
    .port_state_in_12_0_3  (subBytes_out_12_0_3            ), //i
    .port_state_in_12_0_4  (subBytes_out_12_0_4            ), //i
    .port_state_in_12_0_5  (subBytes_out_12_0_5            ), //i
    .port_state_in_12_0_6  (subBytes_out_12_0_6            ), //i
    .port_state_in_12_0_7  (subBytes_out_12_0_7            ), //i
    .port_state_in_12_1_0  (subBytes_out_12_1_0            ), //i
    .port_state_in_12_1_1  (subBytes_out_12_1_1            ), //i
    .port_state_in_12_1_2  (subBytes_out_12_1_2            ), //i
    .port_state_in_12_1_3  (subBytes_out_12_1_3            ), //i
    .port_state_in_12_1_4  (subBytes_out_12_1_4            ), //i
    .port_state_in_12_1_5  (subBytes_out_12_1_5            ), //i
    .port_state_in_12_1_6  (subBytes_out_12_1_6            ), //i
    .port_state_in_12_1_7  (subBytes_out_12_1_7            ), //i
    .port_state_in_13_0_0  (subBytes_out_13_0_0            ), //i
    .port_state_in_13_0_1  (subBytes_out_13_0_1            ), //i
    .port_state_in_13_0_2  (subBytes_out_13_0_2            ), //i
    .port_state_in_13_0_3  (subBytes_out_13_0_3            ), //i
    .port_state_in_13_0_4  (subBytes_out_13_0_4            ), //i
    .port_state_in_13_0_5  (subBytes_out_13_0_5            ), //i
    .port_state_in_13_0_6  (subBytes_out_13_0_6            ), //i
    .port_state_in_13_0_7  (subBytes_out_13_0_7            ), //i
    .port_state_in_13_1_0  (subBytes_out_13_1_0            ), //i
    .port_state_in_13_1_1  (subBytes_out_13_1_1            ), //i
    .port_state_in_13_1_2  (subBytes_out_13_1_2            ), //i
    .port_state_in_13_1_3  (subBytes_out_13_1_3            ), //i
    .port_state_in_13_1_4  (subBytes_out_13_1_4            ), //i
    .port_state_in_13_1_5  (subBytes_out_13_1_5            ), //i
    .port_state_in_13_1_6  (subBytes_out_13_1_6            ), //i
    .port_state_in_13_1_7  (subBytes_out_13_1_7            ), //i
    .port_state_in_14_0_0  (subBytes_out_14_0_0            ), //i
    .port_state_in_14_0_1  (subBytes_out_14_0_1            ), //i
    .port_state_in_14_0_2  (subBytes_out_14_0_2            ), //i
    .port_state_in_14_0_3  (subBytes_out_14_0_3            ), //i
    .port_state_in_14_0_4  (subBytes_out_14_0_4            ), //i
    .port_state_in_14_0_5  (subBytes_out_14_0_5            ), //i
    .port_state_in_14_0_6  (subBytes_out_14_0_6            ), //i
    .port_state_in_14_0_7  (subBytes_out_14_0_7            ), //i
    .port_state_in_14_1_0  (subBytes_out_14_1_0            ), //i
    .port_state_in_14_1_1  (subBytes_out_14_1_1            ), //i
    .port_state_in_14_1_2  (subBytes_out_14_1_2            ), //i
    .port_state_in_14_1_3  (subBytes_out_14_1_3            ), //i
    .port_state_in_14_1_4  (subBytes_out_14_1_4            ), //i
    .port_state_in_14_1_5  (subBytes_out_14_1_5            ), //i
    .port_state_in_14_1_6  (subBytes_out_14_1_6            ), //i
    .port_state_in_14_1_7  (subBytes_out_14_1_7            ), //i
    .port_state_in_15_0_0  (subBytes_out_15_0_0            ), //i
    .port_state_in_15_0_1  (subBytes_out_15_0_1            ), //i
    .port_state_in_15_0_2  (subBytes_out_15_0_2            ), //i
    .port_state_in_15_0_3  (subBytes_out_15_0_3            ), //i
    .port_state_in_15_0_4  (subBytes_out_15_0_4            ), //i
    .port_state_in_15_0_5  (subBytes_out_15_0_5            ), //i
    .port_state_in_15_0_6  (subBytes_out_15_0_6            ), //i
    .port_state_in_15_0_7  (subBytes_out_15_0_7            ), //i
    .port_state_in_15_1_0  (subBytes_out_15_1_0            ), //i
    .port_state_in_15_1_1  (subBytes_out_15_1_1            ), //i
    .port_state_in_15_1_2  (subBytes_out_15_1_2            ), //i
    .port_state_in_15_1_3  (subBytes_out_15_1_3            ), //i
    .port_state_in_15_1_4  (subBytes_out_15_1_4            ), //i
    .port_state_in_15_1_5  (subBytes_out_15_1_5            ), //i
    .port_state_in_15_1_6  (subBytes_out_15_1_6            ), //i
    .port_state_in_15_1_7  (subBytes_out_15_1_7            ), //i
    .port_state_out_0_0_0  (shiftRows_port_state_out_0_0_0 ), //o
    .port_state_out_0_0_1  (shiftRows_port_state_out_0_0_1 ), //o
    .port_state_out_0_0_2  (shiftRows_port_state_out_0_0_2 ), //o
    .port_state_out_0_0_3  (shiftRows_port_state_out_0_0_3 ), //o
    .port_state_out_0_0_4  (shiftRows_port_state_out_0_0_4 ), //o
    .port_state_out_0_0_5  (shiftRows_port_state_out_0_0_5 ), //o
    .port_state_out_0_0_6  (shiftRows_port_state_out_0_0_6 ), //o
    .port_state_out_0_0_7  (shiftRows_port_state_out_0_0_7 ), //o
    .port_state_out_0_1_0  (shiftRows_port_state_out_0_1_0 ), //o
    .port_state_out_0_1_1  (shiftRows_port_state_out_0_1_1 ), //o
    .port_state_out_0_1_2  (shiftRows_port_state_out_0_1_2 ), //o
    .port_state_out_0_1_3  (shiftRows_port_state_out_0_1_3 ), //o
    .port_state_out_0_1_4  (shiftRows_port_state_out_0_1_4 ), //o
    .port_state_out_0_1_5  (shiftRows_port_state_out_0_1_5 ), //o
    .port_state_out_0_1_6  (shiftRows_port_state_out_0_1_6 ), //o
    .port_state_out_0_1_7  (shiftRows_port_state_out_0_1_7 ), //o
    .port_state_out_1_0_0  (shiftRows_port_state_out_1_0_0 ), //o
    .port_state_out_1_0_1  (shiftRows_port_state_out_1_0_1 ), //o
    .port_state_out_1_0_2  (shiftRows_port_state_out_1_0_2 ), //o
    .port_state_out_1_0_3  (shiftRows_port_state_out_1_0_3 ), //o
    .port_state_out_1_0_4  (shiftRows_port_state_out_1_0_4 ), //o
    .port_state_out_1_0_5  (shiftRows_port_state_out_1_0_5 ), //o
    .port_state_out_1_0_6  (shiftRows_port_state_out_1_0_6 ), //o
    .port_state_out_1_0_7  (shiftRows_port_state_out_1_0_7 ), //o
    .port_state_out_1_1_0  (shiftRows_port_state_out_1_1_0 ), //o
    .port_state_out_1_1_1  (shiftRows_port_state_out_1_1_1 ), //o
    .port_state_out_1_1_2  (shiftRows_port_state_out_1_1_2 ), //o
    .port_state_out_1_1_3  (shiftRows_port_state_out_1_1_3 ), //o
    .port_state_out_1_1_4  (shiftRows_port_state_out_1_1_4 ), //o
    .port_state_out_1_1_5  (shiftRows_port_state_out_1_1_5 ), //o
    .port_state_out_1_1_6  (shiftRows_port_state_out_1_1_6 ), //o
    .port_state_out_1_1_7  (shiftRows_port_state_out_1_1_7 ), //o
    .port_state_out_2_0_0  (shiftRows_port_state_out_2_0_0 ), //o
    .port_state_out_2_0_1  (shiftRows_port_state_out_2_0_1 ), //o
    .port_state_out_2_0_2  (shiftRows_port_state_out_2_0_2 ), //o
    .port_state_out_2_0_3  (shiftRows_port_state_out_2_0_3 ), //o
    .port_state_out_2_0_4  (shiftRows_port_state_out_2_0_4 ), //o
    .port_state_out_2_0_5  (shiftRows_port_state_out_2_0_5 ), //o
    .port_state_out_2_0_6  (shiftRows_port_state_out_2_0_6 ), //o
    .port_state_out_2_0_7  (shiftRows_port_state_out_2_0_7 ), //o
    .port_state_out_2_1_0  (shiftRows_port_state_out_2_1_0 ), //o
    .port_state_out_2_1_1  (shiftRows_port_state_out_2_1_1 ), //o
    .port_state_out_2_1_2  (shiftRows_port_state_out_2_1_2 ), //o
    .port_state_out_2_1_3  (shiftRows_port_state_out_2_1_3 ), //o
    .port_state_out_2_1_4  (shiftRows_port_state_out_2_1_4 ), //o
    .port_state_out_2_1_5  (shiftRows_port_state_out_2_1_5 ), //o
    .port_state_out_2_1_6  (shiftRows_port_state_out_2_1_6 ), //o
    .port_state_out_2_1_7  (shiftRows_port_state_out_2_1_7 ), //o
    .port_state_out_3_0_0  (shiftRows_port_state_out_3_0_0 ), //o
    .port_state_out_3_0_1  (shiftRows_port_state_out_3_0_1 ), //o
    .port_state_out_3_0_2  (shiftRows_port_state_out_3_0_2 ), //o
    .port_state_out_3_0_3  (shiftRows_port_state_out_3_0_3 ), //o
    .port_state_out_3_0_4  (shiftRows_port_state_out_3_0_4 ), //o
    .port_state_out_3_0_5  (shiftRows_port_state_out_3_0_5 ), //o
    .port_state_out_3_0_6  (shiftRows_port_state_out_3_0_6 ), //o
    .port_state_out_3_0_7  (shiftRows_port_state_out_3_0_7 ), //o
    .port_state_out_3_1_0  (shiftRows_port_state_out_3_1_0 ), //o
    .port_state_out_3_1_1  (shiftRows_port_state_out_3_1_1 ), //o
    .port_state_out_3_1_2  (shiftRows_port_state_out_3_1_2 ), //o
    .port_state_out_3_1_3  (shiftRows_port_state_out_3_1_3 ), //o
    .port_state_out_3_1_4  (shiftRows_port_state_out_3_1_4 ), //o
    .port_state_out_3_1_5  (shiftRows_port_state_out_3_1_5 ), //o
    .port_state_out_3_1_6  (shiftRows_port_state_out_3_1_6 ), //o
    .port_state_out_3_1_7  (shiftRows_port_state_out_3_1_7 ), //o
    .port_state_out_4_0_0  (shiftRows_port_state_out_4_0_0 ), //o
    .port_state_out_4_0_1  (shiftRows_port_state_out_4_0_1 ), //o
    .port_state_out_4_0_2  (shiftRows_port_state_out_4_0_2 ), //o
    .port_state_out_4_0_3  (shiftRows_port_state_out_4_0_3 ), //o
    .port_state_out_4_0_4  (shiftRows_port_state_out_4_0_4 ), //o
    .port_state_out_4_0_5  (shiftRows_port_state_out_4_0_5 ), //o
    .port_state_out_4_0_6  (shiftRows_port_state_out_4_0_6 ), //o
    .port_state_out_4_0_7  (shiftRows_port_state_out_4_0_7 ), //o
    .port_state_out_4_1_0  (shiftRows_port_state_out_4_1_0 ), //o
    .port_state_out_4_1_1  (shiftRows_port_state_out_4_1_1 ), //o
    .port_state_out_4_1_2  (shiftRows_port_state_out_4_1_2 ), //o
    .port_state_out_4_1_3  (shiftRows_port_state_out_4_1_3 ), //o
    .port_state_out_4_1_4  (shiftRows_port_state_out_4_1_4 ), //o
    .port_state_out_4_1_5  (shiftRows_port_state_out_4_1_5 ), //o
    .port_state_out_4_1_6  (shiftRows_port_state_out_4_1_6 ), //o
    .port_state_out_4_1_7  (shiftRows_port_state_out_4_1_7 ), //o
    .port_state_out_5_0_0  (shiftRows_port_state_out_5_0_0 ), //o
    .port_state_out_5_0_1  (shiftRows_port_state_out_5_0_1 ), //o
    .port_state_out_5_0_2  (shiftRows_port_state_out_5_0_2 ), //o
    .port_state_out_5_0_3  (shiftRows_port_state_out_5_0_3 ), //o
    .port_state_out_5_0_4  (shiftRows_port_state_out_5_0_4 ), //o
    .port_state_out_5_0_5  (shiftRows_port_state_out_5_0_5 ), //o
    .port_state_out_5_0_6  (shiftRows_port_state_out_5_0_6 ), //o
    .port_state_out_5_0_7  (shiftRows_port_state_out_5_0_7 ), //o
    .port_state_out_5_1_0  (shiftRows_port_state_out_5_1_0 ), //o
    .port_state_out_5_1_1  (shiftRows_port_state_out_5_1_1 ), //o
    .port_state_out_5_1_2  (shiftRows_port_state_out_5_1_2 ), //o
    .port_state_out_5_1_3  (shiftRows_port_state_out_5_1_3 ), //o
    .port_state_out_5_1_4  (shiftRows_port_state_out_5_1_4 ), //o
    .port_state_out_5_1_5  (shiftRows_port_state_out_5_1_5 ), //o
    .port_state_out_5_1_6  (shiftRows_port_state_out_5_1_6 ), //o
    .port_state_out_5_1_7  (shiftRows_port_state_out_5_1_7 ), //o
    .port_state_out_6_0_0  (shiftRows_port_state_out_6_0_0 ), //o
    .port_state_out_6_0_1  (shiftRows_port_state_out_6_0_1 ), //o
    .port_state_out_6_0_2  (shiftRows_port_state_out_6_0_2 ), //o
    .port_state_out_6_0_3  (shiftRows_port_state_out_6_0_3 ), //o
    .port_state_out_6_0_4  (shiftRows_port_state_out_6_0_4 ), //o
    .port_state_out_6_0_5  (shiftRows_port_state_out_6_0_5 ), //o
    .port_state_out_6_0_6  (shiftRows_port_state_out_6_0_6 ), //o
    .port_state_out_6_0_7  (shiftRows_port_state_out_6_0_7 ), //o
    .port_state_out_6_1_0  (shiftRows_port_state_out_6_1_0 ), //o
    .port_state_out_6_1_1  (shiftRows_port_state_out_6_1_1 ), //o
    .port_state_out_6_1_2  (shiftRows_port_state_out_6_1_2 ), //o
    .port_state_out_6_1_3  (shiftRows_port_state_out_6_1_3 ), //o
    .port_state_out_6_1_4  (shiftRows_port_state_out_6_1_4 ), //o
    .port_state_out_6_1_5  (shiftRows_port_state_out_6_1_5 ), //o
    .port_state_out_6_1_6  (shiftRows_port_state_out_6_1_6 ), //o
    .port_state_out_6_1_7  (shiftRows_port_state_out_6_1_7 ), //o
    .port_state_out_7_0_0  (shiftRows_port_state_out_7_0_0 ), //o
    .port_state_out_7_0_1  (shiftRows_port_state_out_7_0_1 ), //o
    .port_state_out_7_0_2  (shiftRows_port_state_out_7_0_2 ), //o
    .port_state_out_7_0_3  (shiftRows_port_state_out_7_0_3 ), //o
    .port_state_out_7_0_4  (shiftRows_port_state_out_7_0_4 ), //o
    .port_state_out_7_0_5  (shiftRows_port_state_out_7_0_5 ), //o
    .port_state_out_7_0_6  (shiftRows_port_state_out_7_0_6 ), //o
    .port_state_out_7_0_7  (shiftRows_port_state_out_7_0_7 ), //o
    .port_state_out_7_1_0  (shiftRows_port_state_out_7_1_0 ), //o
    .port_state_out_7_1_1  (shiftRows_port_state_out_7_1_1 ), //o
    .port_state_out_7_1_2  (shiftRows_port_state_out_7_1_2 ), //o
    .port_state_out_7_1_3  (shiftRows_port_state_out_7_1_3 ), //o
    .port_state_out_7_1_4  (shiftRows_port_state_out_7_1_4 ), //o
    .port_state_out_7_1_5  (shiftRows_port_state_out_7_1_5 ), //o
    .port_state_out_7_1_6  (shiftRows_port_state_out_7_1_6 ), //o
    .port_state_out_7_1_7  (shiftRows_port_state_out_7_1_7 ), //o
    .port_state_out_8_0_0  (shiftRows_port_state_out_8_0_0 ), //o
    .port_state_out_8_0_1  (shiftRows_port_state_out_8_0_1 ), //o
    .port_state_out_8_0_2  (shiftRows_port_state_out_8_0_2 ), //o
    .port_state_out_8_0_3  (shiftRows_port_state_out_8_0_3 ), //o
    .port_state_out_8_0_4  (shiftRows_port_state_out_8_0_4 ), //o
    .port_state_out_8_0_5  (shiftRows_port_state_out_8_0_5 ), //o
    .port_state_out_8_0_6  (shiftRows_port_state_out_8_0_6 ), //o
    .port_state_out_8_0_7  (shiftRows_port_state_out_8_0_7 ), //o
    .port_state_out_8_1_0  (shiftRows_port_state_out_8_1_0 ), //o
    .port_state_out_8_1_1  (shiftRows_port_state_out_8_1_1 ), //o
    .port_state_out_8_1_2  (shiftRows_port_state_out_8_1_2 ), //o
    .port_state_out_8_1_3  (shiftRows_port_state_out_8_1_3 ), //o
    .port_state_out_8_1_4  (shiftRows_port_state_out_8_1_4 ), //o
    .port_state_out_8_1_5  (shiftRows_port_state_out_8_1_5 ), //o
    .port_state_out_8_1_6  (shiftRows_port_state_out_8_1_6 ), //o
    .port_state_out_8_1_7  (shiftRows_port_state_out_8_1_7 ), //o
    .port_state_out_9_0_0  (shiftRows_port_state_out_9_0_0 ), //o
    .port_state_out_9_0_1  (shiftRows_port_state_out_9_0_1 ), //o
    .port_state_out_9_0_2  (shiftRows_port_state_out_9_0_2 ), //o
    .port_state_out_9_0_3  (shiftRows_port_state_out_9_0_3 ), //o
    .port_state_out_9_0_4  (shiftRows_port_state_out_9_0_4 ), //o
    .port_state_out_9_0_5  (shiftRows_port_state_out_9_0_5 ), //o
    .port_state_out_9_0_6  (shiftRows_port_state_out_9_0_6 ), //o
    .port_state_out_9_0_7  (shiftRows_port_state_out_9_0_7 ), //o
    .port_state_out_9_1_0  (shiftRows_port_state_out_9_1_0 ), //o
    .port_state_out_9_1_1  (shiftRows_port_state_out_9_1_1 ), //o
    .port_state_out_9_1_2  (shiftRows_port_state_out_9_1_2 ), //o
    .port_state_out_9_1_3  (shiftRows_port_state_out_9_1_3 ), //o
    .port_state_out_9_1_4  (shiftRows_port_state_out_9_1_4 ), //o
    .port_state_out_9_1_5  (shiftRows_port_state_out_9_1_5 ), //o
    .port_state_out_9_1_6  (shiftRows_port_state_out_9_1_6 ), //o
    .port_state_out_9_1_7  (shiftRows_port_state_out_9_1_7 ), //o
    .port_state_out_10_0_0 (shiftRows_port_state_out_10_0_0), //o
    .port_state_out_10_0_1 (shiftRows_port_state_out_10_0_1), //o
    .port_state_out_10_0_2 (shiftRows_port_state_out_10_0_2), //o
    .port_state_out_10_0_3 (shiftRows_port_state_out_10_0_3), //o
    .port_state_out_10_0_4 (shiftRows_port_state_out_10_0_4), //o
    .port_state_out_10_0_5 (shiftRows_port_state_out_10_0_5), //o
    .port_state_out_10_0_6 (shiftRows_port_state_out_10_0_6), //o
    .port_state_out_10_0_7 (shiftRows_port_state_out_10_0_7), //o
    .port_state_out_10_1_0 (shiftRows_port_state_out_10_1_0), //o
    .port_state_out_10_1_1 (shiftRows_port_state_out_10_1_1), //o
    .port_state_out_10_1_2 (shiftRows_port_state_out_10_1_2), //o
    .port_state_out_10_1_3 (shiftRows_port_state_out_10_1_3), //o
    .port_state_out_10_1_4 (shiftRows_port_state_out_10_1_4), //o
    .port_state_out_10_1_5 (shiftRows_port_state_out_10_1_5), //o
    .port_state_out_10_1_6 (shiftRows_port_state_out_10_1_6), //o
    .port_state_out_10_1_7 (shiftRows_port_state_out_10_1_7), //o
    .port_state_out_11_0_0 (shiftRows_port_state_out_11_0_0), //o
    .port_state_out_11_0_1 (shiftRows_port_state_out_11_0_1), //o
    .port_state_out_11_0_2 (shiftRows_port_state_out_11_0_2), //o
    .port_state_out_11_0_3 (shiftRows_port_state_out_11_0_3), //o
    .port_state_out_11_0_4 (shiftRows_port_state_out_11_0_4), //o
    .port_state_out_11_0_5 (shiftRows_port_state_out_11_0_5), //o
    .port_state_out_11_0_6 (shiftRows_port_state_out_11_0_6), //o
    .port_state_out_11_0_7 (shiftRows_port_state_out_11_0_7), //o
    .port_state_out_11_1_0 (shiftRows_port_state_out_11_1_0), //o
    .port_state_out_11_1_1 (shiftRows_port_state_out_11_1_1), //o
    .port_state_out_11_1_2 (shiftRows_port_state_out_11_1_2), //o
    .port_state_out_11_1_3 (shiftRows_port_state_out_11_1_3), //o
    .port_state_out_11_1_4 (shiftRows_port_state_out_11_1_4), //o
    .port_state_out_11_1_5 (shiftRows_port_state_out_11_1_5), //o
    .port_state_out_11_1_6 (shiftRows_port_state_out_11_1_6), //o
    .port_state_out_11_1_7 (shiftRows_port_state_out_11_1_7), //o
    .port_state_out_12_0_0 (shiftRows_port_state_out_12_0_0), //o
    .port_state_out_12_0_1 (shiftRows_port_state_out_12_0_1), //o
    .port_state_out_12_0_2 (shiftRows_port_state_out_12_0_2), //o
    .port_state_out_12_0_3 (shiftRows_port_state_out_12_0_3), //o
    .port_state_out_12_0_4 (shiftRows_port_state_out_12_0_4), //o
    .port_state_out_12_0_5 (shiftRows_port_state_out_12_0_5), //o
    .port_state_out_12_0_6 (shiftRows_port_state_out_12_0_6), //o
    .port_state_out_12_0_7 (shiftRows_port_state_out_12_0_7), //o
    .port_state_out_12_1_0 (shiftRows_port_state_out_12_1_0), //o
    .port_state_out_12_1_1 (shiftRows_port_state_out_12_1_1), //o
    .port_state_out_12_1_2 (shiftRows_port_state_out_12_1_2), //o
    .port_state_out_12_1_3 (shiftRows_port_state_out_12_1_3), //o
    .port_state_out_12_1_4 (shiftRows_port_state_out_12_1_4), //o
    .port_state_out_12_1_5 (shiftRows_port_state_out_12_1_5), //o
    .port_state_out_12_1_6 (shiftRows_port_state_out_12_1_6), //o
    .port_state_out_12_1_7 (shiftRows_port_state_out_12_1_7), //o
    .port_state_out_13_0_0 (shiftRows_port_state_out_13_0_0), //o
    .port_state_out_13_0_1 (shiftRows_port_state_out_13_0_1), //o
    .port_state_out_13_0_2 (shiftRows_port_state_out_13_0_2), //o
    .port_state_out_13_0_3 (shiftRows_port_state_out_13_0_3), //o
    .port_state_out_13_0_4 (shiftRows_port_state_out_13_0_4), //o
    .port_state_out_13_0_5 (shiftRows_port_state_out_13_0_5), //o
    .port_state_out_13_0_6 (shiftRows_port_state_out_13_0_6), //o
    .port_state_out_13_0_7 (shiftRows_port_state_out_13_0_7), //o
    .port_state_out_13_1_0 (shiftRows_port_state_out_13_1_0), //o
    .port_state_out_13_1_1 (shiftRows_port_state_out_13_1_1), //o
    .port_state_out_13_1_2 (shiftRows_port_state_out_13_1_2), //o
    .port_state_out_13_1_3 (shiftRows_port_state_out_13_1_3), //o
    .port_state_out_13_1_4 (shiftRows_port_state_out_13_1_4), //o
    .port_state_out_13_1_5 (shiftRows_port_state_out_13_1_5), //o
    .port_state_out_13_1_6 (shiftRows_port_state_out_13_1_6), //o
    .port_state_out_13_1_7 (shiftRows_port_state_out_13_1_7), //o
    .port_state_out_14_0_0 (shiftRows_port_state_out_14_0_0), //o
    .port_state_out_14_0_1 (shiftRows_port_state_out_14_0_1), //o
    .port_state_out_14_0_2 (shiftRows_port_state_out_14_0_2), //o
    .port_state_out_14_0_3 (shiftRows_port_state_out_14_0_3), //o
    .port_state_out_14_0_4 (shiftRows_port_state_out_14_0_4), //o
    .port_state_out_14_0_5 (shiftRows_port_state_out_14_0_5), //o
    .port_state_out_14_0_6 (shiftRows_port_state_out_14_0_6), //o
    .port_state_out_14_0_7 (shiftRows_port_state_out_14_0_7), //o
    .port_state_out_14_1_0 (shiftRows_port_state_out_14_1_0), //o
    .port_state_out_14_1_1 (shiftRows_port_state_out_14_1_1), //o
    .port_state_out_14_1_2 (shiftRows_port_state_out_14_1_2), //o
    .port_state_out_14_1_3 (shiftRows_port_state_out_14_1_3), //o
    .port_state_out_14_1_4 (shiftRows_port_state_out_14_1_4), //o
    .port_state_out_14_1_5 (shiftRows_port_state_out_14_1_5), //o
    .port_state_out_14_1_6 (shiftRows_port_state_out_14_1_6), //o
    .port_state_out_14_1_7 (shiftRows_port_state_out_14_1_7), //o
    .port_state_out_15_0_0 (shiftRows_port_state_out_15_0_0), //o
    .port_state_out_15_0_1 (shiftRows_port_state_out_15_0_1), //o
    .port_state_out_15_0_2 (shiftRows_port_state_out_15_0_2), //o
    .port_state_out_15_0_3 (shiftRows_port_state_out_15_0_3), //o
    .port_state_out_15_0_4 (shiftRows_port_state_out_15_0_4), //o
    .port_state_out_15_0_5 (shiftRows_port_state_out_15_0_5), //o
    .port_state_out_15_0_6 (shiftRows_port_state_out_15_0_6), //o
    .port_state_out_15_0_7 (shiftRows_port_state_out_15_0_7), //o
    .port_state_out_15_1_0 (shiftRows_port_state_out_15_1_0), //o
    .port_state_out_15_1_1 (shiftRows_port_state_out_15_1_1), //o
    .port_state_out_15_1_2 (shiftRows_port_state_out_15_1_2), //o
    .port_state_out_15_1_3 (shiftRows_port_state_out_15_1_3), //o
    .port_state_out_15_1_4 (shiftRows_port_state_out_15_1_4), //o
    .port_state_out_15_1_5 (shiftRows_port_state_out_15_1_5), //o
    .port_state_out_15_1_6 (shiftRows_port_state_out_15_1_6), //o
    .port_state_out_15_1_7 (shiftRows_port_state_out_15_1_7)  //o
  );
  Aes_MixColumn mixColumns (
    .port_state_in_0_0_0   (shiftRows_port_state_out_0_0_0  ), //i
    .port_state_in_0_0_1   (shiftRows_port_state_out_0_0_1  ), //i
    .port_state_in_0_0_2   (shiftRows_port_state_out_0_0_2  ), //i
    .port_state_in_0_0_3   (shiftRows_port_state_out_0_0_3  ), //i
    .port_state_in_0_0_4   (shiftRows_port_state_out_0_0_4  ), //i
    .port_state_in_0_0_5   (shiftRows_port_state_out_0_0_5  ), //i
    .port_state_in_0_0_6   (shiftRows_port_state_out_0_0_6  ), //i
    .port_state_in_0_0_7   (shiftRows_port_state_out_0_0_7  ), //i
    .port_state_in_0_1_0   (shiftRows_port_state_out_0_1_0  ), //i
    .port_state_in_0_1_1   (shiftRows_port_state_out_0_1_1  ), //i
    .port_state_in_0_1_2   (shiftRows_port_state_out_0_1_2  ), //i
    .port_state_in_0_1_3   (shiftRows_port_state_out_0_1_3  ), //i
    .port_state_in_0_1_4   (shiftRows_port_state_out_0_1_4  ), //i
    .port_state_in_0_1_5   (shiftRows_port_state_out_0_1_5  ), //i
    .port_state_in_0_1_6   (shiftRows_port_state_out_0_1_6  ), //i
    .port_state_in_0_1_7   (shiftRows_port_state_out_0_1_7  ), //i
    .port_state_in_1_0_0   (shiftRows_port_state_out_1_0_0  ), //i
    .port_state_in_1_0_1   (shiftRows_port_state_out_1_0_1  ), //i
    .port_state_in_1_0_2   (shiftRows_port_state_out_1_0_2  ), //i
    .port_state_in_1_0_3   (shiftRows_port_state_out_1_0_3  ), //i
    .port_state_in_1_0_4   (shiftRows_port_state_out_1_0_4  ), //i
    .port_state_in_1_0_5   (shiftRows_port_state_out_1_0_5  ), //i
    .port_state_in_1_0_6   (shiftRows_port_state_out_1_0_6  ), //i
    .port_state_in_1_0_7   (shiftRows_port_state_out_1_0_7  ), //i
    .port_state_in_1_1_0   (shiftRows_port_state_out_1_1_0  ), //i
    .port_state_in_1_1_1   (shiftRows_port_state_out_1_1_1  ), //i
    .port_state_in_1_1_2   (shiftRows_port_state_out_1_1_2  ), //i
    .port_state_in_1_1_3   (shiftRows_port_state_out_1_1_3  ), //i
    .port_state_in_1_1_4   (shiftRows_port_state_out_1_1_4  ), //i
    .port_state_in_1_1_5   (shiftRows_port_state_out_1_1_5  ), //i
    .port_state_in_1_1_6   (shiftRows_port_state_out_1_1_6  ), //i
    .port_state_in_1_1_7   (shiftRows_port_state_out_1_1_7  ), //i
    .port_state_in_2_0_0   (shiftRows_port_state_out_2_0_0  ), //i
    .port_state_in_2_0_1   (shiftRows_port_state_out_2_0_1  ), //i
    .port_state_in_2_0_2   (shiftRows_port_state_out_2_0_2  ), //i
    .port_state_in_2_0_3   (shiftRows_port_state_out_2_0_3  ), //i
    .port_state_in_2_0_4   (shiftRows_port_state_out_2_0_4  ), //i
    .port_state_in_2_0_5   (shiftRows_port_state_out_2_0_5  ), //i
    .port_state_in_2_0_6   (shiftRows_port_state_out_2_0_6  ), //i
    .port_state_in_2_0_7   (shiftRows_port_state_out_2_0_7  ), //i
    .port_state_in_2_1_0   (shiftRows_port_state_out_2_1_0  ), //i
    .port_state_in_2_1_1   (shiftRows_port_state_out_2_1_1  ), //i
    .port_state_in_2_1_2   (shiftRows_port_state_out_2_1_2  ), //i
    .port_state_in_2_1_3   (shiftRows_port_state_out_2_1_3  ), //i
    .port_state_in_2_1_4   (shiftRows_port_state_out_2_1_4  ), //i
    .port_state_in_2_1_5   (shiftRows_port_state_out_2_1_5  ), //i
    .port_state_in_2_1_6   (shiftRows_port_state_out_2_1_6  ), //i
    .port_state_in_2_1_7   (shiftRows_port_state_out_2_1_7  ), //i
    .port_state_in_3_0_0   (shiftRows_port_state_out_3_0_0  ), //i
    .port_state_in_3_0_1   (shiftRows_port_state_out_3_0_1  ), //i
    .port_state_in_3_0_2   (shiftRows_port_state_out_3_0_2  ), //i
    .port_state_in_3_0_3   (shiftRows_port_state_out_3_0_3  ), //i
    .port_state_in_3_0_4   (shiftRows_port_state_out_3_0_4  ), //i
    .port_state_in_3_0_5   (shiftRows_port_state_out_3_0_5  ), //i
    .port_state_in_3_0_6   (shiftRows_port_state_out_3_0_6  ), //i
    .port_state_in_3_0_7   (shiftRows_port_state_out_3_0_7  ), //i
    .port_state_in_3_1_0   (shiftRows_port_state_out_3_1_0  ), //i
    .port_state_in_3_1_1   (shiftRows_port_state_out_3_1_1  ), //i
    .port_state_in_3_1_2   (shiftRows_port_state_out_3_1_2  ), //i
    .port_state_in_3_1_3   (shiftRows_port_state_out_3_1_3  ), //i
    .port_state_in_3_1_4   (shiftRows_port_state_out_3_1_4  ), //i
    .port_state_in_3_1_5   (shiftRows_port_state_out_3_1_5  ), //i
    .port_state_in_3_1_6   (shiftRows_port_state_out_3_1_6  ), //i
    .port_state_in_3_1_7   (shiftRows_port_state_out_3_1_7  ), //i
    .port_state_in_4_0_0   (shiftRows_port_state_out_4_0_0  ), //i
    .port_state_in_4_0_1   (shiftRows_port_state_out_4_0_1  ), //i
    .port_state_in_4_0_2   (shiftRows_port_state_out_4_0_2  ), //i
    .port_state_in_4_0_3   (shiftRows_port_state_out_4_0_3  ), //i
    .port_state_in_4_0_4   (shiftRows_port_state_out_4_0_4  ), //i
    .port_state_in_4_0_5   (shiftRows_port_state_out_4_0_5  ), //i
    .port_state_in_4_0_6   (shiftRows_port_state_out_4_0_6  ), //i
    .port_state_in_4_0_7   (shiftRows_port_state_out_4_0_7  ), //i
    .port_state_in_4_1_0   (shiftRows_port_state_out_4_1_0  ), //i
    .port_state_in_4_1_1   (shiftRows_port_state_out_4_1_1  ), //i
    .port_state_in_4_1_2   (shiftRows_port_state_out_4_1_2  ), //i
    .port_state_in_4_1_3   (shiftRows_port_state_out_4_1_3  ), //i
    .port_state_in_4_1_4   (shiftRows_port_state_out_4_1_4  ), //i
    .port_state_in_4_1_5   (shiftRows_port_state_out_4_1_5  ), //i
    .port_state_in_4_1_6   (shiftRows_port_state_out_4_1_6  ), //i
    .port_state_in_4_1_7   (shiftRows_port_state_out_4_1_7  ), //i
    .port_state_in_5_0_0   (shiftRows_port_state_out_5_0_0  ), //i
    .port_state_in_5_0_1   (shiftRows_port_state_out_5_0_1  ), //i
    .port_state_in_5_0_2   (shiftRows_port_state_out_5_0_2  ), //i
    .port_state_in_5_0_3   (shiftRows_port_state_out_5_0_3  ), //i
    .port_state_in_5_0_4   (shiftRows_port_state_out_5_0_4  ), //i
    .port_state_in_5_0_5   (shiftRows_port_state_out_5_0_5  ), //i
    .port_state_in_5_0_6   (shiftRows_port_state_out_5_0_6  ), //i
    .port_state_in_5_0_7   (shiftRows_port_state_out_5_0_7  ), //i
    .port_state_in_5_1_0   (shiftRows_port_state_out_5_1_0  ), //i
    .port_state_in_5_1_1   (shiftRows_port_state_out_5_1_1  ), //i
    .port_state_in_5_1_2   (shiftRows_port_state_out_5_1_2  ), //i
    .port_state_in_5_1_3   (shiftRows_port_state_out_5_1_3  ), //i
    .port_state_in_5_1_4   (shiftRows_port_state_out_5_1_4  ), //i
    .port_state_in_5_1_5   (shiftRows_port_state_out_5_1_5  ), //i
    .port_state_in_5_1_6   (shiftRows_port_state_out_5_1_6  ), //i
    .port_state_in_5_1_7   (shiftRows_port_state_out_5_1_7  ), //i
    .port_state_in_6_0_0   (shiftRows_port_state_out_6_0_0  ), //i
    .port_state_in_6_0_1   (shiftRows_port_state_out_6_0_1  ), //i
    .port_state_in_6_0_2   (shiftRows_port_state_out_6_0_2  ), //i
    .port_state_in_6_0_3   (shiftRows_port_state_out_6_0_3  ), //i
    .port_state_in_6_0_4   (shiftRows_port_state_out_6_0_4  ), //i
    .port_state_in_6_0_5   (shiftRows_port_state_out_6_0_5  ), //i
    .port_state_in_6_0_6   (shiftRows_port_state_out_6_0_6  ), //i
    .port_state_in_6_0_7   (shiftRows_port_state_out_6_0_7  ), //i
    .port_state_in_6_1_0   (shiftRows_port_state_out_6_1_0  ), //i
    .port_state_in_6_1_1   (shiftRows_port_state_out_6_1_1  ), //i
    .port_state_in_6_1_2   (shiftRows_port_state_out_6_1_2  ), //i
    .port_state_in_6_1_3   (shiftRows_port_state_out_6_1_3  ), //i
    .port_state_in_6_1_4   (shiftRows_port_state_out_6_1_4  ), //i
    .port_state_in_6_1_5   (shiftRows_port_state_out_6_1_5  ), //i
    .port_state_in_6_1_6   (shiftRows_port_state_out_6_1_6  ), //i
    .port_state_in_6_1_7   (shiftRows_port_state_out_6_1_7  ), //i
    .port_state_in_7_0_0   (shiftRows_port_state_out_7_0_0  ), //i
    .port_state_in_7_0_1   (shiftRows_port_state_out_7_0_1  ), //i
    .port_state_in_7_0_2   (shiftRows_port_state_out_7_0_2  ), //i
    .port_state_in_7_0_3   (shiftRows_port_state_out_7_0_3  ), //i
    .port_state_in_7_0_4   (shiftRows_port_state_out_7_0_4  ), //i
    .port_state_in_7_0_5   (shiftRows_port_state_out_7_0_5  ), //i
    .port_state_in_7_0_6   (shiftRows_port_state_out_7_0_6  ), //i
    .port_state_in_7_0_7   (shiftRows_port_state_out_7_0_7  ), //i
    .port_state_in_7_1_0   (shiftRows_port_state_out_7_1_0  ), //i
    .port_state_in_7_1_1   (shiftRows_port_state_out_7_1_1  ), //i
    .port_state_in_7_1_2   (shiftRows_port_state_out_7_1_2  ), //i
    .port_state_in_7_1_3   (shiftRows_port_state_out_7_1_3  ), //i
    .port_state_in_7_1_4   (shiftRows_port_state_out_7_1_4  ), //i
    .port_state_in_7_1_5   (shiftRows_port_state_out_7_1_5  ), //i
    .port_state_in_7_1_6   (shiftRows_port_state_out_7_1_6  ), //i
    .port_state_in_7_1_7   (shiftRows_port_state_out_7_1_7  ), //i
    .port_state_in_8_0_0   (shiftRows_port_state_out_8_0_0  ), //i
    .port_state_in_8_0_1   (shiftRows_port_state_out_8_0_1  ), //i
    .port_state_in_8_0_2   (shiftRows_port_state_out_8_0_2  ), //i
    .port_state_in_8_0_3   (shiftRows_port_state_out_8_0_3  ), //i
    .port_state_in_8_0_4   (shiftRows_port_state_out_8_0_4  ), //i
    .port_state_in_8_0_5   (shiftRows_port_state_out_8_0_5  ), //i
    .port_state_in_8_0_6   (shiftRows_port_state_out_8_0_6  ), //i
    .port_state_in_8_0_7   (shiftRows_port_state_out_8_0_7  ), //i
    .port_state_in_8_1_0   (shiftRows_port_state_out_8_1_0  ), //i
    .port_state_in_8_1_1   (shiftRows_port_state_out_8_1_1  ), //i
    .port_state_in_8_1_2   (shiftRows_port_state_out_8_1_2  ), //i
    .port_state_in_8_1_3   (shiftRows_port_state_out_8_1_3  ), //i
    .port_state_in_8_1_4   (shiftRows_port_state_out_8_1_4  ), //i
    .port_state_in_8_1_5   (shiftRows_port_state_out_8_1_5  ), //i
    .port_state_in_8_1_6   (shiftRows_port_state_out_8_1_6  ), //i
    .port_state_in_8_1_7   (shiftRows_port_state_out_8_1_7  ), //i
    .port_state_in_9_0_0   (shiftRows_port_state_out_9_0_0  ), //i
    .port_state_in_9_0_1   (shiftRows_port_state_out_9_0_1  ), //i
    .port_state_in_9_0_2   (shiftRows_port_state_out_9_0_2  ), //i
    .port_state_in_9_0_3   (shiftRows_port_state_out_9_0_3  ), //i
    .port_state_in_9_0_4   (shiftRows_port_state_out_9_0_4  ), //i
    .port_state_in_9_0_5   (shiftRows_port_state_out_9_0_5  ), //i
    .port_state_in_9_0_6   (shiftRows_port_state_out_9_0_6  ), //i
    .port_state_in_9_0_7   (shiftRows_port_state_out_9_0_7  ), //i
    .port_state_in_9_1_0   (shiftRows_port_state_out_9_1_0  ), //i
    .port_state_in_9_1_1   (shiftRows_port_state_out_9_1_1  ), //i
    .port_state_in_9_1_2   (shiftRows_port_state_out_9_1_2  ), //i
    .port_state_in_9_1_3   (shiftRows_port_state_out_9_1_3  ), //i
    .port_state_in_9_1_4   (shiftRows_port_state_out_9_1_4  ), //i
    .port_state_in_9_1_5   (shiftRows_port_state_out_9_1_5  ), //i
    .port_state_in_9_1_6   (shiftRows_port_state_out_9_1_6  ), //i
    .port_state_in_9_1_7   (shiftRows_port_state_out_9_1_7  ), //i
    .port_state_in_10_0_0  (shiftRows_port_state_out_10_0_0 ), //i
    .port_state_in_10_0_1  (shiftRows_port_state_out_10_0_1 ), //i
    .port_state_in_10_0_2  (shiftRows_port_state_out_10_0_2 ), //i
    .port_state_in_10_0_3  (shiftRows_port_state_out_10_0_3 ), //i
    .port_state_in_10_0_4  (shiftRows_port_state_out_10_0_4 ), //i
    .port_state_in_10_0_5  (shiftRows_port_state_out_10_0_5 ), //i
    .port_state_in_10_0_6  (shiftRows_port_state_out_10_0_6 ), //i
    .port_state_in_10_0_7  (shiftRows_port_state_out_10_0_7 ), //i
    .port_state_in_10_1_0  (shiftRows_port_state_out_10_1_0 ), //i
    .port_state_in_10_1_1  (shiftRows_port_state_out_10_1_1 ), //i
    .port_state_in_10_1_2  (shiftRows_port_state_out_10_1_2 ), //i
    .port_state_in_10_1_3  (shiftRows_port_state_out_10_1_3 ), //i
    .port_state_in_10_1_4  (shiftRows_port_state_out_10_1_4 ), //i
    .port_state_in_10_1_5  (shiftRows_port_state_out_10_1_5 ), //i
    .port_state_in_10_1_6  (shiftRows_port_state_out_10_1_6 ), //i
    .port_state_in_10_1_7  (shiftRows_port_state_out_10_1_7 ), //i
    .port_state_in_11_0_0  (shiftRows_port_state_out_11_0_0 ), //i
    .port_state_in_11_0_1  (shiftRows_port_state_out_11_0_1 ), //i
    .port_state_in_11_0_2  (shiftRows_port_state_out_11_0_2 ), //i
    .port_state_in_11_0_3  (shiftRows_port_state_out_11_0_3 ), //i
    .port_state_in_11_0_4  (shiftRows_port_state_out_11_0_4 ), //i
    .port_state_in_11_0_5  (shiftRows_port_state_out_11_0_5 ), //i
    .port_state_in_11_0_6  (shiftRows_port_state_out_11_0_6 ), //i
    .port_state_in_11_0_7  (shiftRows_port_state_out_11_0_7 ), //i
    .port_state_in_11_1_0  (shiftRows_port_state_out_11_1_0 ), //i
    .port_state_in_11_1_1  (shiftRows_port_state_out_11_1_1 ), //i
    .port_state_in_11_1_2  (shiftRows_port_state_out_11_1_2 ), //i
    .port_state_in_11_1_3  (shiftRows_port_state_out_11_1_3 ), //i
    .port_state_in_11_1_4  (shiftRows_port_state_out_11_1_4 ), //i
    .port_state_in_11_1_5  (shiftRows_port_state_out_11_1_5 ), //i
    .port_state_in_11_1_6  (shiftRows_port_state_out_11_1_6 ), //i
    .port_state_in_11_1_7  (shiftRows_port_state_out_11_1_7 ), //i
    .port_state_in_12_0_0  (shiftRows_port_state_out_12_0_0 ), //i
    .port_state_in_12_0_1  (shiftRows_port_state_out_12_0_1 ), //i
    .port_state_in_12_0_2  (shiftRows_port_state_out_12_0_2 ), //i
    .port_state_in_12_0_3  (shiftRows_port_state_out_12_0_3 ), //i
    .port_state_in_12_0_4  (shiftRows_port_state_out_12_0_4 ), //i
    .port_state_in_12_0_5  (shiftRows_port_state_out_12_0_5 ), //i
    .port_state_in_12_0_6  (shiftRows_port_state_out_12_0_6 ), //i
    .port_state_in_12_0_7  (shiftRows_port_state_out_12_0_7 ), //i
    .port_state_in_12_1_0  (shiftRows_port_state_out_12_1_0 ), //i
    .port_state_in_12_1_1  (shiftRows_port_state_out_12_1_1 ), //i
    .port_state_in_12_1_2  (shiftRows_port_state_out_12_1_2 ), //i
    .port_state_in_12_1_3  (shiftRows_port_state_out_12_1_3 ), //i
    .port_state_in_12_1_4  (shiftRows_port_state_out_12_1_4 ), //i
    .port_state_in_12_1_5  (shiftRows_port_state_out_12_1_5 ), //i
    .port_state_in_12_1_6  (shiftRows_port_state_out_12_1_6 ), //i
    .port_state_in_12_1_7  (shiftRows_port_state_out_12_1_7 ), //i
    .port_state_in_13_0_0  (shiftRows_port_state_out_13_0_0 ), //i
    .port_state_in_13_0_1  (shiftRows_port_state_out_13_0_1 ), //i
    .port_state_in_13_0_2  (shiftRows_port_state_out_13_0_2 ), //i
    .port_state_in_13_0_3  (shiftRows_port_state_out_13_0_3 ), //i
    .port_state_in_13_0_4  (shiftRows_port_state_out_13_0_4 ), //i
    .port_state_in_13_0_5  (shiftRows_port_state_out_13_0_5 ), //i
    .port_state_in_13_0_6  (shiftRows_port_state_out_13_0_6 ), //i
    .port_state_in_13_0_7  (shiftRows_port_state_out_13_0_7 ), //i
    .port_state_in_13_1_0  (shiftRows_port_state_out_13_1_0 ), //i
    .port_state_in_13_1_1  (shiftRows_port_state_out_13_1_1 ), //i
    .port_state_in_13_1_2  (shiftRows_port_state_out_13_1_2 ), //i
    .port_state_in_13_1_3  (shiftRows_port_state_out_13_1_3 ), //i
    .port_state_in_13_1_4  (shiftRows_port_state_out_13_1_4 ), //i
    .port_state_in_13_1_5  (shiftRows_port_state_out_13_1_5 ), //i
    .port_state_in_13_1_6  (shiftRows_port_state_out_13_1_6 ), //i
    .port_state_in_13_1_7  (shiftRows_port_state_out_13_1_7 ), //i
    .port_state_in_14_0_0  (shiftRows_port_state_out_14_0_0 ), //i
    .port_state_in_14_0_1  (shiftRows_port_state_out_14_0_1 ), //i
    .port_state_in_14_0_2  (shiftRows_port_state_out_14_0_2 ), //i
    .port_state_in_14_0_3  (shiftRows_port_state_out_14_0_3 ), //i
    .port_state_in_14_0_4  (shiftRows_port_state_out_14_0_4 ), //i
    .port_state_in_14_0_5  (shiftRows_port_state_out_14_0_5 ), //i
    .port_state_in_14_0_6  (shiftRows_port_state_out_14_0_6 ), //i
    .port_state_in_14_0_7  (shiftRows_port_state_out_14_0_7 ), //i
    .port_state_in_14_1_0  (shiftRows_port_state_out_14_1_0 ), //i
    .port_state_in_14_1_1  (shiftRows_port_state_out_14_1_1 ), //i
    .port_state_in_14_1_2  (shiftRows_port_state_out_14_1_2 ), //i
    .port_state_in_14_1_3  (shiftRows_port_state_out_14_1_3 ), //i
    .port_state_in_14_1_4  (shiftRows_port_state_out_14_1_4 ), //i
    .port_state_in_14_1_5  (shiftRows_port_state_out_14_1_5 ), //i
    .port_state_in_14_1_6  (shiftRows_port_state_out_14_1_6 ), //i
    .port_state_in_14_1_7  (shiftRows_port_state_out_14_1_7 ), //i
    .port_state_in_15_0_0  (shiftRows_port_state_out_15_0_0 ), //i
    .port_state_in_15_0_1  (shiftRows_port_state_out_15_0_1 ), //i
    .port_state_in_15_0_2  (shiftRows_port_state_out_15_0_2 ), //i
    .port_state_in_15_0_3  (shiftRows_port_state_out_15_0_3 ), //i
    .port_state_in_15_0_4  (shiftRows_port_state_out_15_0_4 ), //i
    .port_state_in_15_0_5  (shiftRows_port_state_out_15_0_5 ), //i
    .port_state_in_15_0_6  (shiftRows_port_state_out_15_0_6 ), //i
    .port_state_in_15_0_7  (shiftRows_port_state_out_15_0_7 ), //i
    .port_state_in_15_1_0  (shiftRows_port_state_out_15_1_0 ), //i
    .port_state_in_15_1_1  (shiftRows_port_state_out_15_1_1 ), //i
    .port_state_in_15_1_2  (shiftRows_port_state_out_15_1_2 ), //i
    .port_state_in_15_1_3  (shiftRows_port_state_out_15_1_3 ), //i
    .port_state_in_15_1_4  (shiftRows_port_state_out_15_1_4 ), //i
    .port_state_in_15_1_5  (shiftRows_port_state_out_15_1_5 ), //i
    .port_state_in_15_1_6  (shiftRows_port_state_out_15_1_6 ), //i
    .port_state_in_15_1_7  (shiftRows_port_state_out_15_1_7 ), //i
    .port_state_out_0_0_0  (mixColumns_port_state_out_0_0_0 ), //o
    .port_state_out_0_0_1  (mixColumns_port_state_out_0_0_1 ), //o
    .port_state_out_0_0_2  (mixColumns_port_state_out_0_0_2 ), //o
    .port_state_out_0_0_3  (mixColumns_port_state_out_0_0_3 ), //o
    .port_state_out_0_0_4  (mixColumns_port_state_out_0_0_4 ), //o
    .port_state_out_0_0_5  (mixColumns_port_state_out_0_0_5 ), //o
    .port_state_out_0_0_6  (mixColumns_port_state_out_0_0_6 ), //o
    .port_state_out_0_0_7  (mixColumns_port_state_out_0_0_7 ), //o
    .port_state_out_0_1_0  (mixColumns_port_state_out_0_1_0 ), //o
    .port_state_out_0_1_1  (mixColumns_port_state_out_0_1_1 ), //o
    .port_state_out_0_1_2  (mixColumns_port_state_out_0_1_2 ), //o
    .port_state_out_0_1_3  (mixColumns_port_state_out_0_1_3 ), //o
    .port_state_out_0_1_4  (mixColumns_port_state_out_0_1_4 ), //o
    .port_state_out_0_1_5  (mixColumns_port_state_out_0_1_5 ), //o
    .port_state_out_0_1_6  (mixColumns_port_state_out_0_1_6 ), //o
    .port_state_out_0_1_7  (mixColumns_port_state_out_0_1_7 ), //o
    .port_state_out_1_0_0  (mixColumns_port_state_out_1_0_0 ), //o
    .port_state_out_1_0_1  (mixColumns_port_state_out_1_0_1 ), //o
    .port_state_out_1_0_2  (mixColumns_port_state_out_1_0_2 ), //o
    .port_state_out_1_0_3  (mixColumns_port_state_out_1_0_3 ), //o
    .port_state_out_1_0_4  (mixColumns_port_state_out_1_0_4 ), //o
    .port_state_out_1_0_5  (mixColumns_port_state_out_1_0_5 ), //o
    .port_state_out_1_0_6  (mixColumns_port_state_out_1_0_6 ), //o
    .port_state_out_1_0_7  (mixColumns_port_state_out_1_0_7 ), //o
    .port_state_out_1_1_0  (mixColumns_port_state_out_1_1_0 ), //o
    .port_state_out_1_1_1  (mixColumns_port_state_out_1_1_1 ), //o
    .port_state_out_1_1_2  (mixColumns_port_state_out_1_1_2 ), //o
    .port_state_out_1_1_3  (mixColumns_port_state_out_1_1_3 ), //o
    .port_state_out_1_1_4  (mixColumns_port_state_out_1_1_4 ), //o
    .port_state_out_1_1_5  (mixColumns_port_state_out_1_1_5 ), //o
    .port_state_out_1_1_6  (mixColumns_port_state_out_1_1_6 ), //o
    .port_state_out_1_1_7  (mixColumns_port_state_out_1_1_7 ), //o
    .port_state_out_2_0_0  (mixColumns_port_state_out_2_0_0 ), //o
    .port_state_out_2_0_1  (mixColumns_port_state_out_2_0_1 ), //o
    .port_state_out_2_0_2  (mixColumns_port_state_out_2_0_2 ), //o
    .port_state_out_2_0_3  (mixColumns_port_state_out_2_0_3 ), //o
    .port_state_out_2_0_4  (mixColumns_port_state_out_2_0_4 ), //o
    .port_state_out_2_0_5  (mixColumns_port_state_out_2_0_5 ), //o
    .port_state_out_2_0_6  (mixColumns_port_state_out_2_0_6 ), //o
    .port_state_out_2_0_7  (mixColumns_port_state_out_2_0_7 ), //o
    .port_state_out_2_1_0  (mixColumns_port_state_out_2_1_0 ), //o
    .port_state_out_2_1_1  (mixColumns_port_state_out_2_1_1 ), //o
    .port_state_out_2_1_2  (mixColumns_port_state_out_2_1_2 ), //o
    .port_state_out_2_1_3  (mixColumns_port_state_out_2_1_3 ), //o
    .port_state_out_2_1_4  (mixColumns_port_state_out_2_1_4 ), //o
    .port_state_out_2_1_5  (mixColumns_port_state_out_2_1_5 ), //o
    .port_state_out_2_1_6  (mixColumns_port_state_out_2_1_6 ), //o
    .port_state_out_2_1_7  (mixColumns_port_state_out_2_1_7 ), //o
    .port_state_out_3_0_0  (mixColumns_port_state_out_3_0_0 ), //o
    .port_state_out_3_0_1  (mixColumns_port_state_out_3_0_1 ), //o
    .port_state_out_3_0_2  (mixColumns_port_state_out_3_0_2 ), //o
    .port_state_out_3_0_3  (mixColumns_port_state_out_3_0_3 ), //o
    .port_state_out_3_0_4  (mixColumns_port_state_out_3_0_4 ), //o
    .port_state_out_3_0_5  (mixColumns_port_state_out_3_0_5 ), //o
    .port_state_out_3_0_6  (mixColumns_port_state_out_3_0_6 ), //o
    .port_state_out_3_0_7  (mixColumns_port_state_out_3_0_7 ), //o
    .port_state_out_3_1_0  (mixColumns_port_state_out_3_1_0 ), //o
    .port_state_out_3_1_1  (mixColumns_port_state_out_3_1_1 ), //o
    .port_state_out_3_1_2  (mixColumns_port_state_out_3_1_2 ), //o
    .port_state_out_3_1_3  (mixColumns_port_state_out_3_1_3 ), //o
    .port_state_out_3_1_4  (mixColumns_port_state_out_3_1_4 ), //o
    .port_state_out_3_1_5  (mixColumns_port_state_out_3_1_5 ), //o
    .port_state_out_3_1_6  (mixColumns_port_state_out_3_1_6 ), //o
    .port_state_out_3_1_7  (mixColumns_port_state_out_3_1_7 ), //o
    .port_state_out_4_0_0  (mixColumns_port_state_out_4_0_0 ), //o
    .port_state_out_4_0_1  (mixColumns_port_state_out_4_0_1 ), //o
    .port_state_out_4_0_2  (mixColumns_port_state_out_4_0_2 ), //o
    .port_state_out_4_0_3  (mixColumns_port_state_out_4_0_3 ), //o
    .port_state_out_4_0_4  (mixColumns_port_state_out_4_0_4 ), //o
    .port_state_out_4_0_5  (mixColumns_port_state_out_4_0_5 ), //o
    .port_state_out_4_0_6  (mixColumns_port_state_out_4_0_6 ), //o
    .port_state_out_4_0_7  (mixColumns_port_state_out_4_0_7 ), //o
    .port_state_out_4_1_0  (mixColumns_port_state_out_4_1_0 ), //o
    .port_state_out_4_1_1  (mixColumns_port_state_out_4_1_1 ), //o
    .port_state_out_4_1_2  (mixColumns_port_state_out_4_1_2 ), //o
    .port_state_out_4_1_3  (mixColumns_port_state_out_4_1_3 ), //o
    .port_state_out_4_1_4  (mixColumns_port_state_out_4_1_4 ), //o
    .port_state_out_4_1_5  (mixColumns_port_state_out_4_1_5 ), //o
    .port_state_out_4_1_6  (mixColumns_port_state_out_4_1_6 ), //o
    .port_state_out_4_1_7  (mixColumns_port_state_out_4_1_7 ), //o
    .port_state_out_5_0_0  (mixColumns_port_state_out_5_0_0 ), //o
    .port_state_out_5_0_1  (mixColumns_port_state_out_5_0_1 ), //o
    .port_state_out_5_0_2  (mixColumns_port_state_out_5_0_2 ), //o
    .port_state_out_5_0_3  (mixColumns_port_state_out_5_0_3 ), //o
    .port_state_out_5_0_4  (mixColumns_port_state_out_5_0_4 ), //o
    .port_state_out_5_0_5  (mixColumns_port_state_out_5_0_5 ), //o
    .port_state_out_5_0_6  (mixColumns_port_state_out_5_0_6 ), //o
    .port_state_out_5_0_7  (mixColumns_port_state_out_5_0_7 ), //o
    .port_state_out_5_1_0  (mixColumns_port_state_out_5_1_0 ), //o
    .port_state_out_5_1_1  (mixColumns_port_state_out_5_1_1 ), //o
    .port_state_out_5_1_2  (mixColumns_port_state_out_5_1_2 ), //o
    .port_state_out_5_1_3  (mixColumns_port_state_out_5_1_3 ), //o
    .port_state_out_5_1_4  (mixColumns_port_state_out_5_1_4 ), //o
    .port_state_out_5_1_5  (mixColumns_port_state_out_5_1_5 ), //o
    .port_state_out_5_1_6  (mixColumns_port_state_out_5_1_6 ), //o
    .port_state_out_5_1_7  (mixColumns_port_state_out_5_1_7 ), //o
    .port_state_out_6_0_0  (mixColumns_port_state_out_6_0_0 ), //o
    .port_state_out_6_0_1  (mixColumns_port_state_out_6_0_1 ), //o
    .port_state_out_6_0_2  (mixColumns_port_state_out_6_0_2 ), //o
    .port_state_out_6_0_3  (mixColumns_port_state_out_6_0_3 ), //o
    .port_state_out_6_0_4  (mixColumns_port_state_out_6_0_4 ), //o
    .port_state_out_6_0_5  (mixColumns_port_state_out_6_0_5 ), //o
    .port_state_out_6_0_6  (mixColumns_port_state_out_6_0_6 ), //o
    .port_state_out_6_0_7  (mixColumns_port_state_out_6_0_7 ), //o
    .port_state_out_6_1_0  (mixColumns_port_state_out_6_1_0 ), //o
    .port_state_out_6_1_1  (mixColumns_port_state_out_6_1_1 ), //o
    .port_state_out_6_1_2  (mixColumns_port_state_out_6_1_2 ), //o
    .port_state_out_6_1_3  (mixColumns_port_state_out_6_1_3 ), //o
    .port_state_out_6_1_4  (mixColumns_port_state_out_6_1_4 ), //o
    .port_state_out_6_1_5  (mixColumns_port_state_out_6_1_5 ), //o
    .port_state_out_6_1_6  (mixColumns_port_state_out_6_1_6 ), //o
    .port_state_out_6_1_7  (mixColumns_port_state_out_6_1_7 ), //o
    .port_state_out_7_0_0  (mixColumns_port_state_out_7_0_0 ), //o
    .port_state_out_7_0_1  (mixColumns_port_state_out_7_0_1 ), //o
    .port_state_out_7_0_2  (mixColumns_port_state_out_7_0_2 ), //o
    .port_state_out_7_0_3  (mixColumns_port_state_out_7_0_3 ), //o
    .port_state_out_7_0_4  (mixColumns_port_state_out_7_0_4 ), //o
    .port_state_out_7_0_5  (mixColumns_port_state_out_7_0_5 ), //o
    .port_state_out_7_0_6  (mixColumns_port_state_out_7_0_6 ), //o
    .port_state_out_7_0_7  (mixColumns_port_state_out_7_0_7 ), //o
    .port_state_out_7_1_0  (mixColumns_port_state_out_7_1_0 ), //o
    .port_state_out_7_1_1  (mixColumns_port_state_out_7_1_1 ), //o
    .port_state_out_7_1_2  (mixColumns_port_state_out_7_1_2 ), //o
    .port_state_out_7_1_3  (mixColumns_port_state_out_7_1_3 ), //o
    .port_state_out_7_1_4  (mixColumns_port_state_out_7_1_4 ), //o
    .port_state_out_7_1_5  (mixColumns_port_state_out_7_1_5 ), //o
    .port_state_out_7_1_6  (mixColumns_port_state_out_7_1_6 ), //o
    .port_state_out_7_1_7  (mixColumns_port_state_out_7_1_7 ), //o
    .port_state_out_8_0_0  (mixColumns_port_state_out_8_0_0 ), //o
    .port_state_out_8_0_1  (mixColumns_port_state_out_8_0_1 ), //o
    .port_state_out_8_0_2  (mixColumns_port_state_out_8_0_2 ), //o
    .port_state_out_8_0_3  (mixColumns_port_state_out_8_0_3 ), //o
    .port_state_out_8_0_4  (mixColumns_port_state_out_8_0_4 ), //o
    .port_state_out_8_0_5  (mixColumns_port_state_out_8_0_5 ), //o
    .port_state_out_8_0_6  (mixColumns_port_state_out_8_0_6 ), //o
    .port_state_out_8_0_7  (mixColumns_port_state_out_8_0_7 ), //o
    .port_state_out_8_1_0  (mixColumns_port_state_out_8_1_0 ), //o
    .port_state_out_8_1_1  (mixColumns_port_state_out_8_1_1 ), //o
    .port_state_out_8_1_2  (mixColumns_port_state_out_8_1_2 ), //o
    .port_state_out_8_1_3  (mixColumns_port_state_out_8_1_3 ), //o
    .port_state_out_8_1_4  (mixColumns_port_state_out_8_1_4 ), //o
    .port_state_out_8_1_5  (mixColumns_port_state_out_8_1_5 ), //o
    .port_state_out_8_1_6  (mixColumns_port_state_out_8_1_6 ), //o
    .port_state_out_8_1_7  (mixColumns_port_state_out_8_1_7 ), //o
    .port_state_out_9_0_0  (mixColumns_port_state_out_9_0_0 ), //o
    .port_state_out_9_0_1  (mixColumns_port_state_out_9_0_1 ), //o
    .port_state_out_9_0_2  (mixColumns_port_state_out_9_0_2 ), //o
    .port_state_out_9_0_3  (mixColumns_port_state_out_9_0_3 ), //o
    .port_state_out_9_0_4  (mixColumns_port_state_out_9_0_4 ), //o
    .port_state_out_9_0_5  (mixColumns_port_state_out_9_0_5 ), //o
    .port_state_out_9_0_6  (mixColumns_port_state_out_9_0_6 ), //o
    .port_state_out_9_0_7  (mixColumns_port_state_out_9_0_7 ), //o
    .port_state_out_9_1_0  (mixColumns_port_state_out_9_1_0 ), //o
    .port_state_out_9_1_1  (mixColumns_port_state_out_9_1_1 ), //o
    .port_state_out_9_1_2  (mixColumns_port_state_out_9_1_2 ), //o
    .port_state_out_9_1_3  (mixColumns_port_state_out_9_1_3 ), //o
    .port_state_out_9_1_4  (mixColumns_port_state_out_9_1_4 ), //o
    .port_state_out_9_1_5  (mixColumns_port_state_out_9_1_5 ), //o
    .port_state_out_9_1_6  (mixColumns_port_state_out_9_1_6 ), //o
    .port_state_out_9_1_7  (mixColumns_port_state_out_9_1_7 ), //o
    .port_state_out_10_0_0 (mixColumns_port_state_out_10_0_0), //o
    .port_state_out_10_0_1 (mixColumns_port_state_out_10_0_1), //o
    .port_state_out_10_0_2 (mixColumns_port_state_out_10_0_2), //o
    .port_state_out_10_0_3 (mixColumns_port_state_out_10_0_3), //o
    .port_state_out_10_0_4 (mixColumns_port_state_out_10_0_4), //o
    .port_state_out_10_0_5 (mixColumns_port_state_out_10_0_5), //o
    .port_state_out_10_0_6 (mixColumns_port_state_out_10_0_6), //o
    .port_state_out_10_0_7 (mixColumns_port_state_out_10_0_7), //o
    .port_state_out_10_1_0 (mixColumns_port_state_out_10_1_0), //o
    .port_state_out_10_1_1 (mixColumns_port_state_out_10_1_1), //o
    .port_state_out_10_1_2 (mixColumns_port_state_out_10_1_2), //o
    .port_state_out_10_1_3 (mixColumns_port_state_out_10_1_3), //o
    .port_state_out_10_1_4 (mixColumns_port_state_out_10_1_4), //o
    .port_state_out_10_1_5 (mixColumns_port_state_out_10_1_5), //o
    .port_state_out_10_1_6 (mixColumns_port_state_out_10_1_6), //o
    .port_state_out_10_1_7 (mixColumns_port_state_out_10_1_7), //o
    .port_state_out_11_0_0 (mixColumns_port_state_out_11_0_0), //o
    .port_state_out_11_0_1 (mixColumns_port_state_out_11_0_1), //o
    .port_state_out_11_0_2 (mixColumns_port_state_out_11_0_2), //o
    .port_state_out_11_0_3 (mixColumns_port_state_out_11_0_3), //o
    .port_state_out_11_0_4 (mixColumns_port_state_out_11_0_4), //o
    .port_state_out_11_0_5 (mixColumns_port_state_out_11_0_5), //o
    .port_state_out_11_0_6 (mixColumns_port_state_out_11_0_6), //o
    .port_state_out_11_0_7 (mixColumns_port_state_out_11_0_7), //o
    .port_state_out_11_1_0 (mixColumns_port_state_out_11_1_0), //o
    .port_state_out_11_1_1 (mixColumns_port_state_out_11_1_1), //o
    .port_state_out_11_1_2 (mixColumns_port_state_out_11_1_2), //o
    .port_state_out_11_1_3 (mixColumns_port_state_out_11_1_3), //o
    .port_state_out_11_1_4 (mixColumns_port_state_out_11_1_4), //o
    .port_state_out_11_1_5 (mixColumns_port_state_out_11_1_5), //o
    .port_state_out_11_1_6 (mixColumns_port_state_out_11_1_6), //o
    .port_state_out_11_1_7 (mixColumns_port_state_out_11_1_7), //o
    .port_state_out_12_0_0 (mixColumns_port_state_out_12_0_0), //o
    .port_state_out_12_0_1 (mixColumns_port_state_out_12_0_1), //o
    .port_state_out_12_0_2 (mixColumns_port_state_out_12_0_2), //o
    .port_state_out_12_0_3 (mixColumns_port_state_out_12_0_3), //o
    .port_state_out_12_0_4 (mixColumns_port_state_out_12_0_4), //o
    .port_state_out_12_0_5 (mixColumns_port_state_out_12_0_5), //o
    .port_state_out_12_0_6 (mixColumns_port_state_out_12_0_6), //o
    .port_state_out_12_0_7 (mixColumns_port_state_out_12_0_7), //o
    .port_state_out_12_1_0 (mixColumns_port_state_out_12_1_0), //o
    .port_state_out_12_1_1 (mixColumns_port_state_out_12_1_1), //o
    .port_state_out_12_1_2 (mixColumns_port_state_out_12_1_2), //o
    .port_state_out_12_1_3 (mixColumns_port_state_out_12_1_3), //o
    .port_state_out_12_1_4 (mixColumns_port_state_out_12_1_4), //o
    .port_state_out_12_1_5 (mixColumns_port_state_out_12_1_5), //o
    .port_state_out_12_1_6 (mixColumns_port_state_out_12_1_6), //o
    .port_state_out_12_1_7 (mixColumns_port_state_out_12_1_7), //o
    .port_state_out_13_0_0 (mixColumns_port_state_out_13_0_0), //o
    .port_state_out_13_0_1 (mixColumns_port_state_out_13_0_1), //o
    .port_state_out_13_0_2 (mixColumns_port_state_out_13_0_2), //o
    .port_state_out_13_0_3 (mixColumns_port_state_out_13_0_3), //o
    .port_state_out_13_0_4 (mixColumns_port_state_out_13_0_4), //o
    .port_state_out_13_0_5 (mixColumns_port_state_out_13_0_5), //o
    .port_state_out_13_0_6 (mixColumns_port_state_out_13_0_6), //o
    .port_state_out_13_0_7 (mixColumns_port_state_out_13_0_7), //o
    .port_state_out_13_1_0 (mixColumns_port_state_out_13_1_0), //o
    .port_state_out_13_1_1 (mixColumns_port_state_out_13_1_1), //o
    .port_state_out_13_1_2 (mixColumns_port_state_out_13_1_2), //o
    .port_state_out_13_1_3 (mixColumns_port_state_out_13_1_3), //o
    .port_state_out_13_1_4 (mixColumns_port_state_out_13_1_4), //o
    .port_state_out_13_1_5 (mixColumns_port_state_out_13_1_5), //o
    .port_state_out_13_1_6 (mixColumns_port_state_out_13_1_6), //o
    .port_state_out_13_1_7 (mixColumns_port_state_out_13_1_7), //o
    .port_state_out_14_0_0 (mixColumns_port_state_out_14_0_0), //o
    .port_state_out_14_0_1 (mixColumns_port_state_out_14_0_1), //o
    .port_state_out_14_0_2 (mixColumns_port_state_out_14_0_2), //o
    .port_state_out_14_0_3 (mixColumns_port_state_out_14_0_3), //o
    .port_state_out_14_0_4 (mixColumns_port_state_out_14_0_4), //o
    .port_state_out_14_0_5 (mixColumns_port_state_out_14_0_5), //o
    .port_state_out_14_0_6 (mixColumns_port_state_out_14_0_6), //o
    .port_state_out_14_0_7 (mixColumns_port_state_out_14_0_7), //o
    .port_state_out_14_1_0 (mixColumns_port_state_out_14_1_0), //o
    .port_state_out_14_1_1 (mixColumns_port_state_out_14_1_1), //o
    .port_state_out_14_1_2 (mixColumns_port_state_out_14_1_2), //o
    .port_state_out_14_1_3 (mixColumns_port_state_out_14_1_3), //o
    .port_state_out_14_1_4 (mixColumns_port_state_out_14_1_4), //o
    .port_state_out_14_1_5 (mixColumns_port_state_out_14_1_5), //o
    .port_state_out_14_1_6 (mixColumns_port_state_out_14_1_6), //o
    .port_state_out_14_1_7 (mixColumns_port_state_out_14_1_7), //o
    .port_state_out_15_0_0 (mixColumns_port_state_out_15_0_0), //o
    .port_state_out_15_0_1 (mixColumns_port_state_out_15_0_1), //o
    .port_state_out_15_0_2 (mixColumns_port_state_out_15_0_2), //o
    .port_state_out_15_0_3 (mixColumns_port_state_out_15_0_3), //o
    .port_state_out_15_0_4 (mixColumns_port_state_out_15_0_4), //o
    .port_state_out_15_0_5 (mixColumns_port_state_out_15_0_5), //o
    .port_state_out_15_0_6 (mixColumns_port_state_out_15_0_6), //o
    .port_state_out_15_0_7 (mixColumns_port_state_out_15_0_7), //o
    .port_state_out_15_1_0 (mixColumns_port_state_out_15_1_0), //o
    .port_state_out_15_1_1 (mixColumns_port_state_out_15_1_1), //o
    .port_state_out_15_1_2 (mixColumns_port_state_out_15_1_2), //o
    .port_state_out_15_1_3 (mixColumns_port_state_out_15_1_3), //o
    .port_state_out_15_1_4 (mixColumns_port_state_out_15_1_4), //o
    .port_state_out_15_1_5 (mixColumns_port_state_out_15_1_5), //o
    .port_state_out_15_1_6 (mixColumns_port_state_out_15_1_6), //o
    .port_state_out_15_1_7 (mixColumns_port_state_out_15_1_7)  //o
  );
  assign subBytes_out_0_0_0 = sbox_AES_Canright_CMS_2shares_16_port_o_0_0;
  assign subBytes_out_0_0_1 = sbox_AES_Canright_CMS_2shares_16_port_o_0_1;
  assign subBytes_out_0_0_2 = sbox_AES_Canright_CMS_2shares_16_port_o_0_2;
  assign subBytes_out_0_0_3 = sbox_AES_Canright_CMS_2shares_16_port_o_0_3;
  assign subBytes_out_0_0_4 = sbox_AES_Canright_CMS_2shares_16_port_o_0_4;
  assign subBytes_out_0_0_5 = sbox_AES_Canright_CMS_2shares_16_port_o_0_5;
  assign subBytes_out_0_0_6 = sbox_AES_Canright_CMS_2shares_16_port_o_0_6;
  assign subBytes_out_0_0_7 = sbox_AES_Canright_CMS_2shares_16_port_o_0_7;
  assign subBytes_out_0_1_0 = sbox_AES_Canright_CMS_2shares_16_port_o_1_0;
  assign subBytes_out_0_1_1 = sbox_AES_Canright_CMS_2shares_16_port_o_1_1;
  assign subBytes_out_0_1_2 = sbox_AES_Canright_CMS_2shares_16_port_o_1_2;
  assign subBytes_out_0_1_3 = sbox_AES_Canright_CMS_2shares_16_port_o_1_3;
  assign subBytes_out_0_1_4 = sbox_AES_Canright_CMS_2shares_16_port_o_1_4;
  assign subBytes_out_0_1_5 = sbox_AES_Canright_CMS_2shares_16_port_o_1_5;
  assign subBytes_out_0_1_6 = sbox_AES_Canright_CMS_2shares_16_port_o_1_6;
  assign subBytes_out_0_1_7 = sbox_AES_Canright_CMS_2shares_16_port_o_1_7;
  assign subBytes_out_1_0_0 = sbox_AES_Canright_CMS_2shares_17_port_o_0_0;
  assign subBytes_out_1_0_1 = sbox_AES_Canright_CMS_2shares_17_port_o_0_1;
  assign subBytes_out_1_0_2 = sbox_AES_Canright_CMS_2shares_17_port_o_0_2;
  assign subBytes_out_1_0_3 = sbox_AES_Canright_CMS_2shares_17_port_o_0_3;
  assign subBytes_out_1_0_4 = sbox_AES_Canright_CMS_2shares_17_port_o_0_4;
  assign subBytes_out_1_0_5 = sbox_AES_Canright_CMS_2shares_17_port_o_0_5;
  assign subBytes_out_1_0_6 = sbox_AES_Canright_CMS_2shares_17_port_o_0_6;
  assign subBytes_out_1_0_7 = sbox_AES_Canright_CMS_2shares_17_port_o_0_7;
  assign subBytes_out_1_1_0 = sbox_AES_Canright_CMS_2shares_17_port_o_1_0;
  assign subBytes_out_1_1_1 = sbox_AES_Canright_CMS_2shares_17_port_o_1_1;
  assign subBytes_out_1_1_2 = sbox_AES_Canright_CMS_2shares_17_port_o_1_2;
  assign subBytes_out_1_1_3 = sbox_AES_Canright_CMS_2shares_17_port_o_1_3;
  assign subBytes_out_1_1_4 = sbox_AES_Canright_CMS_2shares_17_port_o_1_4;
  assign subBytes_out_1_1_5 = sbox_AES_Canright_CMS_2shares_17_port_o_1_5;
  assign subBytes_out_1_1_6 = sbox_AES_Canright_CMS_2shares_17_port_o_1_6;
  assign subBytes_out_1_1_7 = sbox_AES_Canright_CMS_2shares_17_port_o_1_7;
  assign subBytes_out_2_0_0 = sbox_AES_Canright_CMS_2shares_18_port_o_0_0;
  assign subBytes_out_2_0_1 = sbox_AES_Canright_CMS_2shares_18_port_o_0_1;
  assign subBytes_out_2_0_2 = sbox_AES_Canright_CMS_2shares_18_port_o_0_2;
  assign subBytes_out_2_0_3 = sbox_AES_Canright_CMS_2shares_18_port_o_0_3;
  assign subBytes_out_2_0_4 = sbox_AES_Canright_CMS_2shares_18_port_o_0_4;
  assign subBytes_out_2_0_5 = sbox_AES_Canright_CMS_2shares_18_port_o_0_5;
  assign subBytes_out_2_0_6 = sbox_AES_Canright_CMS_2shares_18_port_o_0_6;
  assign subBytes_out_2_0_7 = sbox_AES_Canright_CMS_2shares_18_port_o_0_7;
  assign subBytes_out_2_1_0 = sbox_AES_Canright_CMS_2shares_18_port_o_1_0;
  assign subBytes_out_2_1_1 = sbox_AES_Canright_CMS_2shares_18_port_o_1_1;
  assign subBytes_out_2_1_2 = sbox_AES_Canright_CMS_2shares_18_port_o_1_2;
  assign subBytes_out_2_1_3 = sbox_AES_Canright_CMS_2shares_18_port_o_1_3;
  assign subBytes_out_2_1_4 = sbox_AES_Canright_CMS_2shares_18_port_o_1_4;
  assign subBytes_out_2_1_5 = sbox_AES_Canright_CMS_2shares_18_port_o_1_5;
  assign subBytes_out_2_1_6 = sbox_AES_Canright_CMS_2shares_18_port_o_1_6;
  assign subBytes_out_2_1_7 = sbox_AES_Canright_CMS_2shares_18_port_o_1_7;
  assign subBytes_out_3_0_0 = sbox_AES_Canright_CMS_2shares_19_port_o_0_0;
  assign subBytes_out_3_0_1 = sbox_AES_Canright_CMS_2shares_19_port_o_0_1;
  assign subBytes_out_3_0_2 = sbox_AES_Canright_CMS_2shares_19_port_o_0_2;
  assign subBytes_out_3_0_3 = sbox_AES_Canright_CMS_2shares_19_port_o_0_3;
  assign subBytes_out_3_0_4 = sbox_AES_Canright_CMS_2shares_19_port_o_0_4;
  assign subBytes_out_3_0_5 = sbox_AES_Canright_CMS_2shares_19_port_o_0_5;
  assign subBytes_out_3_0_6 = sbox_AES_Canright_CMS_2shares_19_port_o_0_6;
  assign subBytes_out_3_0_7 = sbox_AES_Canright_CMS_2shares_19_port_o_0_7;
  assign subBytes_out_3_1_0 = sbox_AES_Canright_CMS_2shares_19_port_o_1_0;
  assign subBytes_out_3_1_1 = sbox_AES_Canright_CMS_2shares_19_port_o_1_1;
  assign subBytes_out_3_1_2 = sbox_AES_Canright_CMS_2shares_19_port_o_1_2;
  assign subBytes_out_3_1_3 = sbox_AES_Canright_CMS_2shares_19_port_o_1_3;
  assign subBytes_out_3_1_4 = sbox_AES_Canright_CMS_2shares_19_port_o_1_4;
  assign subBytes_out_3_1_5 = sbox_AES_Canright_CMS_2shares_19_port_o_1_5;
  assign subBytes_out_3_1_6 = sbox_AES_Canright_CMS_2shares_19_port_o_1_6;
  assign subBytes_out_3_1_7 = sbox_AES_Canright_CMS_2shares_19_port_o_1_7;
  assign subBytes_out_4_0_0 = sbox_AES_Canright_CMS_2shares_20_port_o_0_0;
  assign subBytes_out_4_0_1 = sbox_AES_Canright_CMS_2shares_20_port_o_0_1;
  assign subBytes_out_4_0_2 = sbox_AES_Canright_CMS_2shares_20_port_o_0_2;
  assign subBytes_out_4_0_3 = sbox_AES_Canright_CMS_2shares_20_port_o_0_3;
  assign subBytes_out_4_0_4 = sbox_AES_Canright_CMS_2shares_20_port_o_0_4;
  assign subBytes_out_4_0_5 = sbox_AES_Canright_CMS_2shares_20_port_o_0_5;
  assign subBytes_out_4_0_6 = sbox_AES_Canright_CMS_2shares_20_port_o_0_6;
  assign subBytes_out_4_0_7 = sbox_AES_Canright_CMS_2shares_20_port_o_0_7;
  assign subBytes_out_4_1_0 = sbox_AES_Canright_CMS_2shares_20_port_o_1_0;
  assign subBytes_out_4_1_1 = sbox_AES_Canright_CMS_2shares_20_port_o_1_1;
  assign subBytes_out_4_1_2 = sbox_AES_Canright_CMS_2shares_20_port_o_1_2;
  assign subBytes_out_4_1_3 = sbox_AES_Canright_CMS_2shares_20_port_o_1_3;
  assign subBytes_out_4_1_4 = sbox_AES_Canright_CMS_2shares_20_port_o_1_4;
  assign subBytes_out_4_1_5 = sbox_AES_Canright_CMS_2shares_20_port_o_1_5;
  assign subBytes_out_4_1_6 = sbox_AES_Canright_CMS_2shares_20_port_o_1_6;
  assign subBytes_out_4_1_7 = sbox_AES_Canright_CMS_2shares_20_port_o_1_7;
  assign subBytes_out_5_0_0 = sbox_AES_Canright_CMS_2shares_21_port_o_0_0;
  assign subBytes_out_5_0_1 = sbox_AES_Canright_CMS_2shares_21_port_o_0_1;
  assign subBytes_out_5_0_2 = sbox_AES_Canright_CMS_2shares_21_port_o_0_2;
  assign subBytes_out_5_0_3 = sbox_AES_Canright_CMS_2shares_21_port_o_0_3;
  assign subBytes_out_5_0_4 = sbox_AES_Canright_CMS_2shares_21_port_o_0_4;
  assign subBytes_out_5_0_5 = sbox_AES_Canright_CMS_2shares_21_port_o_0_5;
  assign subBytes_out_5_0_6 = sbox_AES_Canright_CMS_2shares_21_port_o_0_6;
  assign subBytes_out_5_0_7 = sbox_AES_Canright_CMS_2shares_21_port_o_0_7;
  assign subBytes_out_5_1_0 = sbox_AES_Canright_CMS_2shares_21_port_o_1_0;
  assign subBytes_out_5_1_1 = sbox_AES_Canright_CMS_2shares_21_port_o_1_1;
  assign subBytes_out_5_1_2 = sbox_AES_Canright_CMS_2shares_21_port_o_1_2;
  assign subBytes_out_5_1_3 = sbox_AES_Canright_CMS_2shares_21_port_o_1_3;
  assign subBytes_out_5_1_4 = sbox_AES_Canright_CMS_2shares_21_port_o_1_4;
  assign subBytes_out_5_1_5 = sbox_AES_Canright_CMS_2shares_21_port_o_1_5;
  assign subBytes_out_5_1_6 = sbox_AES_Canright_CMS_2shares_21_port_o_1_6;
  assign subBytes_out_5_1_7 = sbox_AES_Canright_CMS_2shares_21_port_o_1_7;
  assign subBytes_out_6_0_0 = sbox_AES_Canright_CMS_2shares_22_port_o_0_0;
  assign subBytes_out_6_0_1 = sbox_AES_Canright_CMS_2shares_22_port_o_0_1;
  assign subBytes_out_6_0_2 = sbox_AES_Canright_CMS_2shares_22_port_o_0_2;
  assign subBytes_out_6_0_3 = sbox_AES_Canright_CMS_2shares_22_port_o_0_3;
  assign subBytes_out_6_0_4 = sbox_AES_Canright_CMS_2shares_22_port_o_0_4;
  assign subBytes_out_6_0_5 = sbox_AES_Canright_CMS_2shares_22_port_o_0_5;
  assign subBytes_out_6_0_6 = sbox_AES_Canright_CMS_2shares_22_port_o_0_6;
  assign subBytes_out_6_0_7 = sbox_AES_Canright_CMS_2shares_22_port_o_0_7;
  assign subBytes_out_6_1_0 = sbox_AES_Canright_CMS_2shares_22_port_o_1_0;
  assign subBytes_out_6_1_1 = sbox_AES_Canright_CMS_2shares_22_port_o_1_1;
  assign subBytes_out_6_1_2 = sbox_AES_Canright_CMS_2shares_22_port_o_1_2;
  assign subBytes_out_6_1_3 = sbox_AES_Canright_CMS_2shares_22_port_o_1_3;
  assign subBytes_out_6_1_4 = sbox_AES_Canright_CMS_2shares_22_port_o_1_4;
  assign subBytes_out_6_1_5 = sbox_AES_Canright_CMS_2shares_22_port_o_1_5;
  assign subBytes_out_6_1_6 = sbox_AES_Canright_CMS_2shares_22_port_o_1_6;
  assign subBytes_out_6_1_7 = sbox_AES_Canright_CMS_2shares_22_port_o_1_7;
  assign subBytes_out_7_0_0 = sbox_AES_Canright_CMS_2shares_23_port_o_0_0;
  assign subBytes_out_7_0_1 = sbox_AES_Canright_CMS_2shares_23_port_o_0_1;
  assign subBytes_out_7_0_2 = sbox_AES_Canright_CMS_2shares_23_port_o_0_2;
  assign subBytes_out_7_0_3 = sbox_AES_Canright_CMS_2shares_23_port_o_0_3;
  assign subBytes_out_7_0_4 = sbox_AES_Canright_CMS_2shares_23_port_o_0_4;
  assign subBytes_out_7_0_5 = sbox_AES_Canright_CMS_2shares_23_port_o_0_5;
  assign subBytes_out_7_0_6 = sbox_AES_Canright_CMS_2shares_23_port_o_0_6;
  assign subBytes_out_7_0_7 = sbox_AES_Canright_CMS_2shares_23_port_o_0_7;
  assign subBytes_out_7_1_0 = sbox_AES_Canright_CMS_2shares_23_port_o_1_0;
  assign subBytes_out_7_1_1 = sbox_AES_Canright_CMS_2shares_23_port_o_1_1;
  assign subBytes_out_7_1_2 = sbox_AES_Canright_CMS_2shares_23_port_o_1_2;
  assign subBytes_out_7_1_3 = sbox_AES_Canright_CMS_2shares_23_port_o_1_3;
  assign subBytes_out_7_1_4 = sbox_AES_Canright_CMS_2shares_23_port_o_1_4;
  assign subBytes_out_7_1_5 = sbox_AES_Canright_CMS_2shares_23_port_o_1_5;
  assign subBytes_out_7_1_6 = sbox_AES_Canright_CMS_2shares_23_port_o_1_6;
  assign subBytes_out_7_1_7 = sbox_AES_Canright_CMS_2shares_23_port_o_1_7;
  assign subBytes_out_8_0_0 = sbox_AES_Canright_CMS_2shares_24_port_o_0_0;
  assign subBytes_out_8_0_1 = sbox_AES_Canright_CMS_2shares_24_port_o_0_1;
  assign subBytes_out_8_0_2 = sbox_AES_Canright_CMS_2shares_24_port_o_0_2;
  assign subBytes_out_8_0_3 = sbox_AES_Canright_CMS_2shares_24_port_o_0_3;
  assign subBytes_out_8_0_4 = sbox_AES_Canright_CMS_2shares_24_port_o_0_4;
  assign subBytes_out_8_0_5 = sbox_AES_Canright_CMS_2shares_24_port_o_0_5;
  assign subBytes_out_8_0_6 = sbox_AES_Canright_CMS_2shares_24_port_o_0_6;
  assign subBytes_out_8_0_7 = sbox_AES_Canright_CMS_2shares_24_port_o_0_7;
  assign subBytes_out_8_1_0 = sbox_AES_Canright_CMS_2shares_24_port_o_1_0;
  assign subBytes_out_8_1_1 = sbox_AES_Canright_CMS_2shares_24_port_o_1_1;
  assign subBytes_out_8_1_2 = sbox_AES_Canright_CMS_2shares_24_port_o_1_2;
  assign subBytes_out_8_1_3 = sbox_AES_Canright_CMS_2shares_24_port_o_1_3;
  assign subBytes_out_8_1_4 = sbox_AES_Canright_CMS_2shares_24_port_o_1_4;
  assign subBytes_out_8_1_5 = sbox_AES_Canright_CMS_2shares_24_port_o_1_5;
  assign subBytes_out_8_1_6 = sbox_AES_Canright_CMS_2shares_24_port_o_1_6;
  assign subBytes_out_8_1_7 = sbox_AES_Canright_CMS_2shares_24_port_o_1_7;
  assign subBytes_out_9_0_0 = sbox_AES_Canright_CMS_2shares_25_port_o_0_0;
  assign subBytes_out_9_0_1 = sbox_AES_Canright_CMS_2shares_25_port_o_0_1;
  assign subBytes_out_9_0_2 = sbox_AES_Canright_CMS_2shares_25_port_o_0_2;
  assign subBytes_out_9_0_3 = sbox_AES_Canright_CMS_2shares_25_port_o_0_3;
  assign subBytes_out_9_0_4 = sbox_AES_Canright_CMS_2shares_25_port_o_0_4;
  assign subBytes_out_9_0_5 = sbox_AES_Canright_CMS_2shares_25_port_o_0_5;
  assign subBytes_out_9_0_6 = sbox_AES_Canright_CMS_2shares_25_port_o_0_6;
  assign subBytes_out_9_0_7 = sbox_AES_Canright_CMS_2shares_25_port_o_0_7;
  assign subBytes_out_9_1_0 = sbox_AES_Canright_CMS_2shares_25_port_o_1_0;
  assign subBytes_out_9_1_1 = sbox_AES_Canright_CMS_2shares_25_port_o_1_1;
  assign subBytes_out_9_1_2 = sbox_AES_Canright_CMS_2shares_25_port_o_1_2;
  assign subBytes_out_9_1_3 = sbox_AES_Canright_CMS_2shares_25_port_o_1_3;
  assign subBytes_out_9_1_4 = sbox_AES_Canright_CMS_2shares_25_port_o_1_4;
  assign subBytes_out_9_1_5 = sbox_AES_Canright_CMS_2shares_25_port_o_1_5;
  assign subBytes_out_9_1_6 = sbox_AES_Canright_CMS_2shares_25_port_o_1_6;
  assign subBytes_out_9_1_7 = sbox_AES_Canright_CMS_2shares_25_port_o_1_7;
  assign subBytes_out_10_0_0 = sbox_AES_Canright_CMS_2shares_26_port_o_0_0;
  assign subBytes_out_10_0_1 = sbox_AES_Canright_CMS_2shares_26_port_o_0_1;
  assign subBytes_out_10_0_2 = sbox_AES_Canright_CMS_2shares_26_port_o_0_2;
  assign subBytes_out_10_0_3 = sbox_AES_Canright_CMS_2shares_26_port_o_0_3;
  assign subBytes_out_10_0_4 = sbox_AES_Canright_CMS_2shares_26_port_o_0_4;
  assign subBytes_out_10_0_5 = sbox_AES_Canright_CMS_2shares_26_port_o_0_5;
  assign subBytes_out_10_0_6 = sbox_AES_Canright_CMS_2shares_26_port_o_0_6;
  assign subBytes_out_10_0_7 = sbox_AES_Canright_CMS_2shares_26_port_o_0_7;
  assign subBytes_out_10_1_0 = sbox_AES_Canright_CMS_2shares_26_port_o_1_0;
  assign subBytes_out_10_1_1 = sbox_AES_Canright_CMS_2shares_26_port_o_1_1;
  assign subBytes_out_10_1_2 = sbox_AES_Canright_CMS_2shares_26_port_o_1_2;
  assign subBytes_out_10_1_3 = sbox_AES_Canright_CMS_2shares_26_port_o_1_3;
  assign subBytes_out_10_1_4 = sbox_AES_Canright_CMS_2shares_26_port_o_1_4;
  assign subBytes_out_10_1_5 = sbox_AES_Canright_CMS_2shares_26_port_o_1_5;
  assign subBytes_out_10_1_6 = sbox_AES_Canright_CMS_2shares_26_port_o_1_6;
  assign subBytes_out_10_1_7 = sbox_AES_Canright_CMS_2shares_26_port_o_1_7;
  assign subBytes_out_11_0_0 = sbox_AES_Canright_CMS_2shares_27_port_o_0_0;
  assign subBytes_out_11_0_1 = sbox_AES_Canright_CMS_2shares_27_port_o_0_1;
  assign subBytes_out_11_0_2 = sbox_AES_Canright_CMS_2shares_27_port_o_0_2;
  assign subBytes_out_11_0_3 = sbox_AES_Canright_CMS_2shares_27_port_o_0_3;
  assign subBytes_out_11_0_4 = sbox_AES_Canright_CMS_2shares_27_port_o_0_4;
  assign subBytes_out_11_0_5 = sbox_AES_Canright_CMS_2shares_27_port_o_0_5;
  assign subBytes_out_11_0_6 = sbox_AES_Canright_CMS_2shares_27_port_o_0_6;
  assign subBytes_out_11_0_7 = sbox_AES_Canright_CMS_2shares_27_port_o_0_7;
  assign subBytes_out_11_1_0 = sbox_AES_Canright_CMS_2shares_27_port_o_1_0;
  assign subBytes_out_11_1_1 = sbox_AES_Canright_CMS_2shares_27_port_o_1_1;
  assign subBytes_out_11_1_2 = sbox_AES_Canright_CMS_2shares_27_port_o_1_2;
  assign subBytes_out_11_1_3 = sbox_AES_Canright_CMS_2shares_27_port_o_1_3;
  assign subBytes_out_11_1_4 = sbox_AES_Canright_CMS_2shares_27_port_o_1_4;
  assign subBytes_out_11_1_5 = sbox_AES_Canright_CMS_2shares_27_port_o_1_5;
  assign subBytes_out_11_1_6 = sbox_AES_Canright_CMS_2shares_27_port_o_1_6;
  assign subBytes_out_11_1_7 = sbox_AES_Canright_CMS_2shares_27_port_o_1_7;
  assign subBytes_out_12_0_0 = sbox_AES_Canright_CMS_2shares_28_port_o_0_0;
  assign subBytes_out_12_0_1 = sbox_AES_Canright_CMS_2shares_28_port_o_0_1;
  assign subBytes_out_12_0_2 = sbox_AES_Canright_CMS_2shares_28_port_o_0_2;
  assign subBytes_out_12_0_3 = sbox_AES_Canright_CMS_2shares_28_port_o_0_3;
  assign subBytes_out_12_0_4 = sbox_AES_Canright_CMS_2shares_28_port_o_0_4;
  assign subBytes_out_12_0_5 = sbox_AES_Canright_CMS_2shares_28_port_o_0_5;
  assign subBytes_out_12_0_6 = sbox_AES_Canright_CMS_2shares_28_port_o_0_6;
  assign subBytes_out_12_0_7 = sbox_AES_Canright_CMS_2shares_28_port_o_0_7;
  assign subBytes_out_12_1_0 = sbox_AES_Canright_CMS_2shares_28_port_o_1_0;
  assign subBytes_out_12_1_1 = sbox_AES_Canright_CMS_2shares_28_port_o_1_1;
  assign subBytes_out_12_1_2 = sbox_AES_Canright_CMS_2shares_28_port_o_1_2;
  assign subBytes_out_12_1_3 = sbox_AES_Canright_CMS_2shares_28_port_o_1_3;
  assign subBytes_out_12_1_4 = sbox_AES_Canright_CMS_2shares_28_port_o_1_4;
  assign subBytes_out_12_1_5 = sbox_AES_Canright_CMS_2shares_28_port_o_1_5;
  assign subBytes_out_12_1_6 = sbox_AES_Canright_CMS_2shares_28_port_o_1_6;
  assign subBytes_out_12_1_7 = sbox_AES_Canright_CMS_2shares_28_port_o_1_7;
  assign subBytes_out_13_0_0 = sbox_AES_Canright_CMS_2shares_29_port_o_0_0;
  assign subBytes_out_13_0_1 = sbox_AES_Canright_CMS_2shares_29_port_o_0_1;
  assign subBytes_out_13_0_2 = sbox_AES_Canright_CMS_2shares_29_port_o_0_2;
  assign subBytes_out_13_0_3 = sbox_AES_Canright_CMS_2shares_29_port_o_0_3;
  assign subBytes_out_13_0_4 = sbox_AES_Canright_CMS_2shares_29_port_o_0_4;
  assign subBytes_out_13_0_5 = sbox_AES_Canright_CMS_2shares_29_port_o_0_5;
  assign subBytes_out_13_0_6 = sbox_AES_Canright_CMS_2shares_29_port_o_0_6;
  assign subBytes_out_13_0_7 = sbox_AES_Canright_CMS_2shares_29_port_o_0_7;
  assign subBytes_out_13_1_0 = sbox_AES_Canright_CMS_2shares_29_port_o_1_0;
  assign subBytes_out_13_1_1 = sbox_AES_Canright_CMS_2shares_29_port_o_1_1;
  assign subBytes_out_13_1_2 = sbox_AES_Canright_CMS_2shares_29_port_o_1_2;
  assign subBytes_out_13_1_3 = sbox_AES_Canright_CMS_2shares_29_port_o_1_3;
  assign subBytes_out_13_1_4 = sbox_AES_Canright_CMS_2shares_29_port_o_1_4;
  assign subBytes_out_13_1_5 = sbox_AES_Canright_CMS_2shares_29_port_o_1_5;
  assign subBytes_out_13_1_6 = sbox_AES_Canright_CMS_2shares_29_port_o_1_6;
  assign subBytes_out_13_1_7 = sbox_AES_Canright_CMS_2shares_29_port_o_1_7;
  assign subBytes_out_14_0_0 = sbox_AES_Canright_CMS_2shares_30_port_o_0_0;
  assign subBytes_out_14_0_1 = sbox_AES_Canright_CMS_2shares_30_port_o_0_1;
  assign subBytes_out_14_0_2 = sbox_AES_Canright_CMS_2shares_30_port_o_0_2;
  assign subBytes_out_14_0_3 = sbox_AES_Canright_CMS_2shares_30_port_o_0_3;
  assign subBytes_out_14_0_4 = sbox_AES_Canright_CMS_2shares_30_port_o_0_4;
  assign subBytes_out_14_0_5 = sbox_AES_Canright_CMS_2shares_30_port_o_0_5;
  assign subBytes_out_14_0_6 = sbox_AES_Canright_CMS_2shares_30_port_o_0_6;
  assign subBytes_out_14_0_7 = sbox_AES_Canright_CMS_2shares_30_port_o_0_7;
  assign subBytes_out_14_1_0 = sbox_AES_Canright_CMS_2shares_30_port_o_1_0;
  assign subBytes_out_14_1_1 = sbox_AES_Canright_CMS_2shares_30_port_o_1_1;
  assign subBytes_out_14_1_2 = sbox_AES_Canright_CMS_2shares_30_port_o_1_2;
  assign subBytes_out_14_1_3 = sbox_AES_Canright_CMS_2shares_30_port_o_1_3;
  assign subBytes_out_14_1_4 = sbox_AES_Canright_CMS_2shares_30_port_o_1_4;
  assign subBytes_out_14_1_5 = sbox_AES_Canright_CMS_2shares_30_port_o_1_5;
  assign subBytes_out_14_1_6 = sbox_AES_Canright_CMS_2shares_30_port_o_1_6;
  assign subBytes_out_14_1_7 = sbox_AES_Canright_CMS_2shares_30_port_o_1_7;
  assign subBytes_out_15_0_0 = sbox_AES_Canright_CMS_2shares_31_port_o_0_0;
  assign subBytes_out_15_0_1 = sbox_AES_Canright_CMS_2shares_31_port_o_0_1;
  assign subBytes_out_15_0_2 = sbox_AES_Canright_CMS_2shares_31_port_o_0_2;
  assign subBytes_out_15_0_3 = sbox_AES_Canright_CMS_2shares_31_port_o_0_3;
  assign subBytes_out_15_0_4 = sbox_AES_Canright_CMS_2shares_31_port_o_0_4;
  assign subBytes_out_15_0_5 = sbox_AES_Canright_CMS_2shares_31_port_o_0_5;
  assign subBytes_out_15_0_6 = sbox_AES_Canright_CMS_2shares_31_port_o_0_6;
  assign subBytes_out_15_0_7 = sbox_AES_Canright_CMS_2shares_31_port_o_0_7;
  assign subBytes_out_15_1_0 = sbox_AES_Canright_CMS_2shares_31_port_o_1_0;
  assign subBytes_out_15_1_1 = sbox_AES_Canright_CMS_2shares_31_port_o_1_1;
  assign subBytes_out_15_1_2 = sbox_AES_Canright_CMS_2shares_31_port_o_1_2;
  assign subBytes_out_15_1_3 = sbox_AES_Canright_CMS_2shares_31_port_o_1_3;
  assign subBytes_out_15_1_4 = sbox_AES_Canright_CMS_2shares_31_port_o_1_4;
  assign subBytes_out_15_1_5 = sbox_AES_Canright_CMS_2shares_31_port_o_1_5;
  assign subBytes_out_15_1_6 = sbox_AES_Canright_CMS_2shares_31_port_o_1_6;
  assign subBytes_out_15_1_7 = sbox_AES_Canright_CMS_2shares_31_port_o_1_7;
  assign port_state_out_0_0_0 = roundReg_0_0_0;
  assign port_state_out_0_0_1 = roundReg_0_0_1;
  assign port_state_out_0_0_2 = roundReg_0_0_2;
  assign port_state_out_0_0_3 = roundReg_0_0_3;
  assign port_state_out_0_0_4 = roundReg_0_0_4;
  assign port_state_out_0_0_5 = roundReg_0_0_5;
  assign port_state_out_0_0_6 = roundReg_0_0_6;
  assign port_state_out_0_0_7 = roundReg_0_0_7;
  assign port_state_out_0_1_0 = roundReg_0_1_0;
  assign port_state_out_0_1_1 = roundReg_0_1_1;
  assign port_state_out_0_1_2 = roundReg_0_1_2;
  assign port_state_out_0_1_3 = roundReg_0_1_3;
  assign port_state_out_0_1_4 = roundReg_0_1_4;
  assign port_state_out_0_1_5 = roundReg_0_1_5;
  assign port_state_out_0_1_6 = roundReg_0_1_6;
  assign port_state_out_0_1_7 = roundReg_0_1_7;
  assign port_state_out_1_0_0 = roundReg_1_0_0;
  assign port_state_out_1_0_1 = roundReg_1_0_1;
  assign port_state_out_1_0_2 = roundReg_1_0_2;
  assign port_state_out_1_0_3 = roundReg_1_0_3;
  assign port_state_out_1_0_4 = roundReg_1_0_4;
  assign port_state_out_1_0_5 = roundReg_1_0_5;
  assign port_state_out_1_0_6 = roundReg_1_0_6;
  assign port_state_out_1_0_7 = roundReg_1_0_7;
  assign port_state_out_1_1_0 = roundReg_1_1_0;
  assign port_state_out_1_1_1 = roundReg_1_1_1;
  assign port_state_out_1_1_2 = roundReg_1_1_2;
  assign port_state_out_1_1_3 = roundReg_1_1_3;
  assign port_state_out_1_1_4 = roundReg_1_1_4;
  assign port_state_out_1_1_5 = roundReg_1_1_5;
  assign port_state_out_1_1_6 = roundReg_1_1_6;
  assign port_state_out_1_1_7 = roundReg_1_1_7;
  assign port_state_out_2_0_0 = roundReg_2_0_0;
  assign port_state_out_2_0_1 = roundReg_2_0_1;
  assign port_state_out_2_0_2 = roundReg_2_0_2;
  assign port_state_out_2_0_3 = roundReg_2_0_3;
  assign port_state_out_2_0_4 = roundReg_2_0_4;
  assign port_state_out_2_0_5 = roundReg_2_0_5;
  assign port_state_out_2_0_6 = roundReg_2_0_6;
  assign port_state_out_2_0_7 = roundReg_2_0_7;
  assign port_state_out_2_1_0 = roundReg_2_1_0;
  assign port_state_out_2_1_1 = roundReg_2_1_1;
  assign port_state_out_2_1_2 = roundReg_2_1_2;
  assign port_state_out_2_1_3 = roundReg_2_1_3;
  assign port_state_out_2_1_4 = roundReg_2_1_4;
  assign port_state_out_2_1_5 = roundReg_2_1_5;
  assign port_state_out_2_1_6 = roundReg_2_1_6;
  assign port_state_out_2_1_7 = roundReg_2_1_7;
  assign port_state_out_3_0_0 = roundReg_3_0_0;
  assign port_state_out_3_0_1 = roundReg_3_0_1;
  assign port_state_out_3_0_2 = roundReg_3_0_2;
  assign port_state_out_3_0_3 = roundReg_3_0_3;
  assign port_state_out_3_0_4 = roundReg_3_0_4;
  assign port_state_out_3_0_5 = roundReg_3_0_5;
  assign port_state_out_3_0_6 = roundReg_3_0_6;
  assign port_state_out_3_0_7 = roundReg_3_0_7;
  assign port_state_out_3_1_0 = roundReg_3_1_0;
  assign port_state_out_3_1_1 = roundReg_3_1_1;
  assign port_state_out_3_1_2 = roundReg_3_1_2;
  assign port_state_out_3_1_3 = roundReg_3_1_3;
  assign port_state_out_3_1_4 = roundReg_3_1_4;
  assign port_state_out_3_1_5 = roundReg_3_1_5;
  assign port_state_out_3_1_6 = roundReg_3_1_6;
  assign port_state_out_3_1_7 = roundReg_3_1_7;
  assign port_state_out_4_0_0 = roundReg_4_0_0;
  assign port_state_out_4_0_1 = roundReg_4_0_1;
  assign port_state_out_4_0_2 = roundReg_4_0_2;
  assign port_state_out_4_0_3 = roundReg_4_0_3;
  assign port_state_out_4_0_4 = roundReg_4_0_4;
  assign port_state_out_4_0_5 = roundReg_4_0_5;
  assign port_state_out_4_0_6 = roundReg_4_0_6;
  assign port_state_out_4_0_7 = roundReg_4_0_7;
  assign port_state_out_4_1_0 = roundReg_4_1_0;
  assign port_state_out_4_1_1 = roundReg_4_1_1;
  assign port_state_out_4_1_2 = roundReg_4_1_2;
  assign port_state_out_4_1_3 = roundReg_4_1_3;
  assign port_state_out_4_1_4 = roundReg_4_1_4;
  assign port_state_out_4_1_5 = roundReg_4_1_5;
  assign port_state_out_4_1_6 = roundReg_4_1_6;
  assign port_state_out_4_1_7 = roundReg_4_1_7;
  assign port_state_out_5_0_0 = roundReg_5_0_0;
  assign port_state_out_5_0_1 = roundReg_5_0_1;
  assign port_state_out_5_0_2 = roundReg_5_0_2;
  assign port_state_out_5_0_3 = roundReg_5_0_3;
  assign port_state_out_5_0_4 = roundReg_5_0_4;
  assign port_state_out_5_0_5 = roundReg_5_0_5;
  assign port_state_out_5_0_6 = roundReg_5_0_6;
  assign port_state_out_5_0_7 = roundReg_5_0_7;
  assign port_state_out_5_1_0 = roundReg_5_1_0;
  assign port_state_out_5_1_1 = roundReg_5_1_1;
  assign port_state_out_5_1_2 = roundReg_5_1_2;
  assign port_state_out_5_1_3 = roundReg_5_1_3;
  assign port_state_out_5_1_4 = roundReg_5_1_4;
  assign port_state_out_5_1_5 = roundReg_5_1_5;
  assign port_state_out_5_1_6 = roundReg_5_1_6;
  assign port_state_out_5_1_7 = roundReg_5_1_7;
  assign port_state_out_6_0_0 = roundReg_6_0_0;
  assign port_state_out_6_0_1 = roundReg_6_0_1;
  assign port_state_out_6_0_2 = roundReg_6_0_2;
  assign port_state_out_6_0_3 = roundReg_6_0_3;
  assign port_state_out_6_0_4 = roundReg_6_0_4;
  assign port_state_out_6_0_5 = roundReg_6_0_5;
  assign port_state_out_6_0_6 = roundReg_6_0_6;
  assign port_state_out_6_0_7 = roundReg_6_0_7;
  assign port_state_out_6_1_0 = roundReg_6_1_0;
  assign port_state_out_6_1_1 = roundReg_6_1_1;
  assign port_state_out_6_1_2 = roundReg_6_1_2;
  assign port_state_out_6_1_3 = roundReg_6_1_3;
  assign port_state_out_6_1_4 = roundReg_6_1_4;
  assign port_state_out_6_1_5 = roundReg_6_1_5;
  assign port_state_out_6_1_6 = roundReg_6_1_6;
  assign port_state_out_6_1_7 = roundReg_6_1_7;
  assign port_state_out_7_0_0 = roundReg_7_0_0;
  assign port_state_out_7_0_1 = roundReg_7_0_1;
  assign port_state_out_7_0_2 = roundReg_7_0_2;
  assign port_state_out_7_0_3 = roundReg_7_0_3;
  assign port_state_out_7_0_4 = roundReg_7_0_4;
  assign port_state_out_7_0_5 = roundReg_7_0_5;
  assign port_state_out_7_0_6 = roundReg_7_0_6;
  assign port_state_out_7_0_7 = roundReg_7_0_7;
  assign port_state_out_7_1_0 = roundReg_7_1_0;
  assign port_state_out_7_1_1 = roundReg_7_1_1;
  assign port_state_out_7_1_2 = roundReg_7_1_2;
  assign port_state_out_7_1_3 = roundReg_7_1_3;
  assign port_state_out_7_1_4 = roundReg_7_1_4;
  assign port_state_out_7_1_5 = roundReg_7_1_5;
  assign port_state_out_7_1_6 = roundReg_7_1_6;
  assign port_state_out_7_1_7 = roundReg_7_1_7;
  assign port_state_out_8_0_0 = roundReg_8_0_0;
  assign port_state_out_8_0_1 = roundReg_8_0_1;
  assign port_state_out_8_0_2 = roundReg_8_0_2;
  assign port_state_out_8_0_3 = roundReg_8_0_3;
  assign port_state_out_8_0_4 = roundReg_8_0_4;
  assign port_state_out_8_0_5 = roundReg_8_0_5;
  assign port_state_out_8_0_6 = roundReg_8_0_6;
  assign port_state_out_8_0_7 = roundReg_8_0_7;
  assign port_state_out_8_1_0 = roundReg_8_1_0;
  assign port_state_out_8_1_1 = roundReg_8_1_1;
  assign port_state_out_8_1_2 = roundReg_8_1_2;
  assign port_state_out_8_1_3 = roundReg_8_1_3;
  assign port_state_out_8_1_4 = roundReg_8_1_4;
  assign port_state_out_8_1_5 = roundReg_8_1_5;
  assign port_state_out_8_1_6 = roundReg_8_1_6;
  assign port_state_out_8_1_7 = roundReg_8_1_7;
  assign port_state_out_9_0_0 = roundReg_9_0_0;
  assign port_state_out_9_0_1 = roundReg_9_0_1;
  assign port_state_out_9_0_2 = roundReg_9_0_2;
  assign port_state_out_9_0_3 = roundReg_9_0_3;
  assign port_state_out_9_0_4 = roundReg_9_0_4;
  assign port_state_out_9_0_5 = roundReg_9_0_5;
  assign port_state_out_9_0_6 = roundReg_9_0_6;
  assign port_state_out_9_0_7 = roundReg_9_0_7;
  assign port_state_out_9_1_0 = roundReg_9_1_0;
  assign port_state_out_9_1_1 = roundReg_9_1_1;
  assign port_state_out_9_1_2 = roundReg_9_1_2;
  assign port_state_out_9_1_3 = roundReg_9_1_3;
  assign port_state_out_9_1_4 = roundReg_9_1_4;
  assign port_state_out_9_1_5 = roundReg_9_1_5;
  assign port_state_out_9_1_6 = roundReg_9_1_6;
  assign port_state_out_9_1_7 = roundReg_9_1_7;
  assign port_state_out_10_0_0 = roundReg_10_0_0;
  assign port_state_out_10_0_1 = roundReg_10_0_1;
  assign port_state_out_10_0_2 = roundReg_10_0_2;
  assign port_state_out_10_0_3 = roundReg_10_0_3;
  assign port_state_out_10_0_4 = roundReg_10_0_4;
  assign port_state_out_10_0_5 = roundReg_10_0_5;
  assign port_state_out_10_0_6 = roundReg_10_0_6;
  assign port_state_out_10_0_7 = roundReg_10_0_7;
  assign port_state_out_10_1_0 = roundReg_10_1_0;
  assign port_state_out_10_1_1 = roundReg_10_1_1;
  assign port_state_out_10_1_2 = roundReg_10_1_2;
  assign port_state_out_10_1_3 = roundReg_10_1_3;
  assign port_state_out_10_1_4 = roundReg_10_1_4;
  assign port_state_out_10_1_5 = roundReg_10_1_5;
  assign port_state_out_10_1_6 = roundReg_10_1_6;
  assign port_state_out_10_1_7 = roundReg_10_1_7;
  assign port_state_out_11_0_0 = roundReg_11_0_0;
  assign port_state_out_11_0_1 = roundReg_11_0_1;
  assign port_state_out_11_0_2 = roundReg_11_0_2;
  assign port_state_out_11_0_3 = roundReg_11_0_3;
  assign port_state_out_11_0_4 = roundReg_11_0_4;
  assign port_state_out_11_0_5 = roundReg_11_0_5;
  assign port_state_out_11_0_6 = roundReg_11_0_6;
  assign port_state_out_11_0_7 = roundReg_11_0_7;
  assign port_state_out_11_1_0 = roundReg_11_1_0;
  assign port_state_out_11_1_1 = roundReg_11_1_1;
  assign port_state_out_11_1_2 = roundReg_11_1_2;
  assign port_state_out_11_1_3 = roundReg_11_1_3;
  assign port_state_out_11_1_4 = roundReg_11_1_4;
  assign port_state_out_11_1_5 = roundReg_11_1_5;
  assign port_state_out_11_1_6 = roundReg_11_1_6;
  assign port_state_out_11_1_7 = roundReg_11_1_7;
  assign port_state_out_12_0_0 = roundReg_12_0_0;
  assign port_state_out_12_0_1 = roundReg_12_0_1;
  assign port_state_out_12_0_2 = roundReg_12_0_2;
  assign port_state_out_12_0_3 = roundReg_12_0_3;
  assign port_state_out_12_0_4 = roundReg_12_0_4;
  assign port_state_out_12_0_5 = roundReg_12_0_5;
  assign port_state_out_12_0_6 = roundReg_12_0_6;
  assign port_state_out_12_0_7 = roundReg_12_0_7;
  assign port_state_out_12_1_0 = roundReg_12_1_0;
  assign port_state_out_12_1_1 = roundReg_12_1_1;
  assign port_state_out_12_1_2 = roundReg_12_1_2;
  assign port_state_out_12_1_3 = roundReg_12_1_3;
  assign port_state_out_12_1_4 = roundReg_12_1_4;
  assign port_state_out_12_1_5 = roundReg_12_1_5;
  assign port_state_out_12_1_6 = roundReg_12_1_6;
  assign port_state_out_12_1_7 = roundReg_12_1_7;
  assign port_state_out_13_0_0 = roundReg_13_0_0;
  assign port_state_out_13_0_1 = roundReg_13_0_1;
  assign port_state_out_13_0_2 = roundReg_13_0_2;
  assign port_state_out_13_0_3 = roundReg_13_0_3;
  assign port_state_out_13_0_4 = roundReg_13_0_4;
  assign port_state_out_13_0_5 = roundReg_13_0_5;
  assign port_state_out_13_0_6 = roundReg_13_0_6;
  assign port_state_out_13_0_7 = roundReg_13_0_7;
  assign port_state_out_13_1_0 = roundReg_13_1_0;
  assign port_state_out_13_1_1 = roundReg_13_1_1;
  assign port_state_out_13_1_2 = roundReg_13_1_2;
  assign port_state_out_13_1_3 = roundReg_13_1_3;
  assign port_state_out_13_1_4 = roundReg_13_1_4;
  assign port_state_out_13_1_5 = roundReg_13_1_5;
  assign port_state_out_13_1_6 = roundReg_13_1_6;
  assign port_state_out_13_1_7 = roundReg_13_1_7;
  assign port_state_out_14_0_0 = roundReg_14_0_0;
  assign port_state_out_14_0_1 = roundReg_14_0_1;
  assign port_state_out_14_0_2 = roundReg_14_0_2;
  assign port_state_out_14_0_3 = roundReg_14_0_3;
  assign port_state_out_14_0_4 = roundReg_14_0_4;
  assign port_state_out_14_0_5 = roundReg_14_0_5;
  assign port_state_out_14_0_6 = roundReg_14_0_6;
  assign port_state_out_14_0_7 = roundReg_14_0_7;
  assign port_state_out_14_1_0 = roundReg_14_1_0;
  assign port_state_out_14_1_1 = roundReg_14_1_1;
  assign port_state_out_14_1_2 = roundReg_14_1_2;
  assign port_state_out_14_1_3 = roundReg_14_1_3;
  assign port_state_out_14_1_4 = roundReg_14_1_4;
  assign port_state_out_14_1_5 = roundReg_14_1_5;
  assign port_state_out_14_1_6 = roundReg_14_1_6;
  assign port_state_out_14_1_7 = roundReg_14_1_7;
  assign port_state_out_15_0_0 = roundReg_15_0_0;
  assign port_state_out_15_0_1 = roundReg_15_0_1;
  assign port_state_out_15_0_2 = roundReg_15_0_2;
  assign port_state_out_15_0_3 = roundReg_15_0_3;
  assign port_state_out_15_0_4 = roundReg_15_0_4;
  assign port_state_out_15_0_5 = roundReg_15_0_5;
  assign port_state_out_15_0_6 = roundReg_15_0_6;
  assign port_state_out_15_0_7 = roundReg_15_0_7;
  assign port_state_out_15_1_0 = roundReg_15_1_0;
  assign port_state_out_15_1_1 = roundReg_15_1_1;
  assign port_state_out_15_1_2 = roundReg_15_1_2;
  assign port_state_out_15_1_3 = roundReg_15_1_3;
  assign port_state_out_15_1_4 = roundReg_15_1_4;
  assign port_state_out_15_1_5 = roundReg_15_1_5;
  assign port_state_out_15_1_6 = roundReg_15_1_6;
  assign port_state_out_15_1_7 = roundReg_15_1_7;
  always @(posedge clk) begin
    roundReg_0_0_0 <= mixColumns_port_state_out_0_0_0;
    roundReg_0_0_1 <= mixColumns_port_state_out_0_0_1;
    roundReg_0_0_2 <= mixColumns_port_state_out_0_0_2;
    roundReg_0_0_3 <= mixColumns_port_state_out_0_0_3;
    roundReg_0_0_4 <= mixColumns_port_state_out_0_0_4;
    roundReg_0_0_5 <= mixColumns_port_state_out_0_0_5;
    roundReg_0_0_6 <= mixColumns_port_state_out_0_0_6;
    roundReg_0_0_7 <= mixColumns_port_state_out_0_0_7;
    roundReg_0_1_0 <= mixColumns_port_state_out_0_1_0;
    roundReg_0_1_1 <= mixColumns_port_state_out_0_1_1;
    roundReg_0_1_2 <= mixColumns_port_state_out_0_1_2;
    roundReg_0_1_3 <= mixColumns_port_state_out_0_1_3;
    roundReg_0_1_4 <= mixColumns_port_state_out_0_1_4;
    roundReg_0_1_5 <= mixColumns_port_state_out_0_1_5;
    roundReg_0_1_6 <= mixColumns_port_state_out_0_1_6;
    roundReg_0_1_7 <= mixColumns_port_state_out_0_1_7;
    roundReg_1_0_0 <= mixColumns_port_state_out_1_0_0;
    roundReg_1_0_1 <= mixColumns_port_state_out_1_0_1;
    roundReg_1_0_2 <= mixColumns_port_state_out_1_0_2;
    roundReg_1_0_3 <= mixColumns_port_state_out_1_0_3;
    roundReg_1_0_4 <= mixColumns_port_state_out_1_0_4;
    roundReg_1_0_5 <= mixColumns_port_state_out_1_0_5;
    roundReg_1_0_6 <= mixColumns_port_state_out_1_0_6;
    roundReg_1_0_7 <= mixColumns_port_state_out_1_0_7;
    roundReg_1_1_0 <= mixColumns_port_state_out_1_1_0;
    roundReg_1_1_1 <= mixColumns_port_state_out_1_1_1;
    roundReg_1_1_2 <= mixColumns_port_state_out_1_1_2;
    roundReg_1_1_3 <= mixColumns_port_state_out_1_1_3;
    roundReg_1_1_4 <= mixColumns_port_state_out_1_1_4;
    roundReg_1_1_5 <= mixColumns_port_state_out_1_1_5;
    roundReg_1_1_6 <= mixColumns_port_state_out_1_1_6;
    roundReg_1_1_7 <= mixColumns_port_state_out_1_1_7;
    roundReg_2_0_0 <= mixColumns_port_state_out_2_0_0;
    roundReg_2_0_1 <= mixColumns_port_state_out_2_0_1;
    roundReg_2_0_2 <= mixColumns_port_state_out_2_0_2;
    roundReg_2_0_3 <= mixColumns_port_state_out_2_0_3;
    roundReg_2_0_4 <= mixColumns_port_state_out_2_0_4;
    roundReg_2_0_5 <= mixColumns_port_state_out_2_0_5;
    roundReg_2_0_6 <= mixColumns_port_state_out_2_0_6;
    roundReg_2_0_7 <= mixColumns_port_state_out_2_0_7;
    roundReg_2_1_0 <= mixColumns_port_state_out_2_1_0;
    roundReg_2_1_1 <= mixColumns_port_state_out_2_1_1;
    roundReg_2_1_2 <= mixColumns_port_state_out_2_1_2;
    roundReg_2_1_3 <= mixColumns_port_state_out_2_1_3;
    roundReg_2_1_4 <= mixColumns_port_state_out_2_1_4;
    roundReg_2_1_5 <= mixColumns_port_state_out_2_1_5;
    roundReg_2_1_6 <= mixColumns_port_state_out_2_1_6;
    roundReg_2_1_7 <= mixColumns_port_state_out_2_1_7;
    roundReg_3_0_0 <= mixColumns_port_state_out_3_0_0;
    roundReg_3_0_1 <= mixColumns_port_state_out_3_0_1;
    roundReg_3_0_2 <= mixColumns_port_state_out_3_0_2;
    roundReg_3_0_3 <= mixColumns_port_state_out_3_0_3;
    roundReg_3_0_4 <= mixColumns_port_state_out_3_0_4;
    roundReg_3_0_5 <= mixColumns_port_state_out_3_0_5;
    roundReg_3_0_6 <= mixColumns_port_state_out_3_0_6;
    roundReg_3_0_7 <= mixColumns_port_state_out_3_0_7;
    roundReg_3_1_0 <= mixColumns_port_state_out_3_1_0;
    roundReg_3_1_1 <= mixColumns_port_state_out_3_1_1;
    roundReg_3_1_2 <= mixColumns_port_state_out_3_1_2;
    roundReg_3_1_3 <= mixColumns_port_state_out_3_1_3;
    roundReg_3_1_4 <= mixColumns_port_state_out_3_1_4;
    roundReg_3_1_5 <= mixColumns_port_state_out_3_1_5;
    roundReg_3_1_6 <= mixColumns_port_state_out_3_1_6;
    roundReg_3_1_7 <= mixColumns_port_state_out_3_1_7;
    roundReg_4_0_0 <= mixColumns_port_state_out_4_0_0;
    roundReg_4_0_1 <= mixColumns_port_state_out_4_0_1;
    roundReg_4_0_2 <= mixColumns_port_state_out_4_0_2;
    roundReg_4_0_3 <= mixColumns_port_state_out_4_0_3;
    roundReg_4_0_4 <= mixColumns_port_state_out_4_0_4;
    roundReg_4_0_5 <= mixColumns_port_state_out_4_0_5;
    roundReg_4_0_6 <= mixColumns_port_state_out_4_0_6;
    roundReg_4_0_7 <= mixColumns_port_state_out_4_0_7;
    roundReg_4_1_0 <= mixColumns_port_state_out_4_1_0;
    roundReg_4_1_1 <= mixColumns_port_state_out_4_1_1;
    roundReg_4_1_2 <= mixColumns_port_state_out_4_1_2;
    roundReg_4_1_3 <= mixColumns_port_state_out_4_1_3;
    roundReg_4_1_4 <= mixColumns_port_state_out_4_1_4;
    roundReg_4_1_5 <= mixColumns_port_state_out_4_1_5;
    roundReg_4_1_6 <= mixColumns_port_state_out_4_1_6;
    roundReg_4_1_7 <= mixColumns_port_state_out_4_1_7;
    roundReg_5_0_0 <= mixColumns_port_state_out_5_0_0;
    roundReg_5_0_1 <= mixColumns_port_state_out_5_0_1;
    roundReg_5_0_2 <= mixColumns_port_state_out_5_0_2;
    roundReg_5_0_3 <= mixColumns_port_state_out_5_0_3;
    roundReg_5_0_4 <= mixColumns_port_state_out_5_0_4;
    roundReg_5_0_5 <= mixColumns_port_state_out_5_0_5;
    roundReg_5_0_6 <= mixColumns_port_state_out_5_0_6;
    roundReg_5_0_7 <= mixColumns_port_state_out_5_0_7;
    roundReg_5_1_0 <= mixColumns_port_state_out_5_1_0;
    roundReg_5_1_1 <= mixColumns_port_state_out_5_1_1;
    roundReg_5_1_2 <= mixColumns_port_state_out_5_1_2;
    roundReg_5_1_3 <= mixColumns_port_state_out_5_1_3;
    roundReg_5_1_4 <= mixColumns_port_state_out_5_1_4;
    roundReg_5_1_5 <= mixColumns_port_state_out_5_1_5;
    roundReg_5_1_6 <= mixColumns_port_state_out_5_1_6;
    roundReg_5_1_7 <= mixColumns_port_state_out_5_1_7;
    roundReg_6_0_0 <= mixColumns_port_state_out_6_0_0;
    roundReg_6_0_1 <= mixColumns_port_state_out_6_0_1;
    roundReg_6_0_2 <= mixColumns_port_state_out_6_0_2;
    roundReg_6_0_3 <= mixColumns_port_state_out_6_0_3;
    roundReg_6_0_4 <= mixColumns_port_state_out_6_0_4;
    roundReg_6_0_5 <= mixColumns_port_state_out_6_0_5;
    roundReg_6_0_6 <= mixColumns_port_state_out_6_0_6;
    roundReg_6_0_7 <= mixColumns_port_state_out_6_0_7;
    roundReg_6_1_0 <= mixColumns_port_state_out_6_1_0;
    roundReg_6_1_1 <= mixColumns_port_state_out_6_1_1;
    roundReg_6_1_2 <= mixColumns_port_state_out_6_1_2;
    roundReg_6_1_3 <= mixColumns_port_state_out_6_1_3;
    roundReg_6_1_4 <= mixColumns_port_state_out_6_1_4;
    roundReg_6_1_5 <= mixColumns_port_state_out_6_1_5;
    roundReg_6_1_6 <= mixColumns_port_state_out_6_1_6;
    roundReg_6_1_7 <= mixColumns_port_state_out_6_1_7;
    roundReg_7_0_0 <= mixColumns_port_state_out_7_0_0;
    roundReg_7_0_1 <= mixColumns_port_state_out_7_0_1;
    roundReg_7_0_2 <= mixColumns_port_state_out_7_0_2;
    roundReg_7_0_3 <= mixColumns_port_state_out_7_0_3;
    roundReg_7_0_4 <= mixColumns_port_state_out_7_0_4;
    roundReg_7_0_5 <= mixColumns_port_state_out_7_0_5;
    roundReg_7_0_6 <= mixColumns_port_state_out_7_0_6;
    roundReg_7_0_7 <= mixColumns_port_state_out_7_0_7;
    roundReg_7_1_0 <= mixColumns_port_state_out_7_1_0;
    roundReg_7_1_1 <= mixColumns_port_state_out_7_1_1;
    roundReg_7_1_2 <= mixColumns_port_state_out_7_1_2;
    roundReg_7_1_3 <= mixColumns_port_state_out_7_1_3;
    roundReg_7_1_4 <= mixColumns_port_state_out_7_1_4;
    roundReg_7_1_5 <= mixColumns_port_state_out_7_1_5;
    roundReg_7_1_6 <= mixColumns_port_state_out_7_1_6;
    roundReg_7_1_7 <= mixColumns_port_state_out_7_1_7;
    roundReg_8_0_0 <= mixColumns_port_state_out_8_0_0;
    roundReg_8_0_1 <= mixColumns_port_state_out_8_0_1;
    roundReg_8_0_2 <= mixColumns_port_state_out_8_0_2;
    roundReg_8_0_3 <= mixColumns_port_state_out_8_0_3;
    roundReg_8_0_4 <= mixColumns_port_state_out_8_0_4;
    roundReg_8_0_5 <= mixColumns_port_state_out_8_0_5;
    roundReg_8_0_6 <= mixColumns_port_state_out_8_0_6;
    roundReg_8_0_7 <= mixColumns_port_state_out_8_0_7;
    roundReg_8_1_0 <= mixColumns_port_state_out_8_1_0;
    roundReg_8_1_1 <= mixColumns_port_state_out_8_1_1;
    roundReg_8_1_2 <= mixColumns_port_state_out_8_1_2;
    roundReg_8_1_3 <= mixColumns_port_state_out_8_1_3;
    roundReg_8_1_4 <= mixColumns_port_state_out_8_1_4;
    roundReg_8_1_5 <= mixColumns_port_state_out_8_1_5;
    roundReg_8_1_6 <= mixColumns_port_state_out_8_1_6;
    roundReg_8_1_7 <= mixColumns_port_state_out_8_1_7;
    roundReg_9_0_0 <= mixColumns_port_state_out_9_0_0;
    roundReg_9_0_1 <= mixColumns_port_state_out_9_0_1;
    roundReg_9_0_2 <= mixColumns_port_state_out_9_0_2;
    roundReg_9_0_3 <= mixColumns_port_state_out_9_0_3;
    roundReg_9_0_4 <= mixColumns_port_state_out_9_0_4;
    roundReg_9_0_5 <= mixColumns_port_state_out_9_0_5;
    roundReg_9_0_6 <= mixColumns_port_state_out_9_0_6;
    roundReg_9_0_7 <= mixColumns_port_state_out_9_0_7;
    roundReg_9_1_0 <= mixColumns_port_state_out_9_1_0;
    roundReg_9_1_1 <= mixColumns_port_state_out_9_1_1;
    roundReg_9_1_2 <= mixColumns_port_state_out_9_1_2;
    roundReg_9_1_3 <= mixColumns_port_state_out_9_1_3;
    roundReg_9_1_4 <= mixColumns_port_state_out_9_1_4;
    roundReg_9_1_5 <= mixColumns_port_state_out_9_1_5;
    roundReg_9_1_6 <= mixColumns_port_state_out_9_1_6;
    roundReg_9_1_7 <= mixColumns_port_state_out_9_1_7;
    roundReg_10_0_0 <= mixColumns_port_state_out_10_0_0;
    roundReg_10_0_1 <= mixColumns_port_state_out_10_0_1;
    roundReg_10_0_2 <= mixColumns_port_state_out_10_0_2;
    roundReg_10_0_3 <= mixColumns_port_state_out_10_0_3;
    roundReg_10_0_4 <= mixColumns_port_state_out_10_0_4;
    roundReg_10_0_5 <= mixColumns_port_state_out_10_0_5;
    roundReg_10_0_6 <= mixColumns_port_state_out_10_0_6;
    roundReg_10_0_7 <= mixColumns_port_state_out_10_0_7;
    roundReg_10_1_0 <= mixColumns_port_state_out_10_1_0;
    roundReg_10_1_1 <= mixColumns_port_state_out_10_1_1;
    roundReg_10_1_2 <= mixColumns_port_state_out_10_1_2;
    roundReg_10_1_3 <= mixColumns_port_state_out_10_1_3;
    roundReg_10_1_4 <= mixColumns_port_state_out_10_1_4;
    roundReg_10_1_5 <= mixColumns_port_state_out_10_1_5;
    roundReg_10_1_6 <= mixColumns_port_state_out_10_1_6;
    roundReg_10_1_7 <= mixColumns_port_state_out_10_1_7;
    roundReg_11_0_0 <= mixColumns_port_state_out_11_0_0;
    roundReg_11_0_1 <= mixColumns_port_state_out_11_0_1;
    roundReg_11_0_2 <= mixColumns_port_state_out_11_0_2;
    roundReg_11_0_3 <= mixColumns_port_state_out_11_0_3;
    roundReg_11_0_4 <= mixColumns_port_state_out_11_0_4;
    roundReg_11_0_5 <= mixColumns_port_state_out_11_0_5;
    roundReg_11_0_6 <= mixColumns_port_state_out_11_0_6;
    roundReg_11_0_7 <= mixColumns_port_state_out_11_0_7;
    roundReg_11_1_0 <= mixColumns_port_state_out_11_1_0;
    roundReg_11_1_1 <= mixColumns_port_state_out_11_1_1;
    roundReg_11_1_2 <= mixColumns_port_state_out_11_1_2;
    roundReg_11_1_3 <= mixColumns_port_state_out_11_1_3;
    roundReg_11_1_4 <= mixColumns_port_state_out_11_1_4;
    roundReg_11_1_5 <= mixColumns_port_state_out_11_1_5;
    roundReg_11_1_6 <= mixColumns_port_state_out_11_1_6;
    roundReg_11_1_7 <= mixColumns_port_state_out_11_1_7;
    roundReg_12_0_0 <= mixColumns_port_state_out_12_0_0;
    roundReg_12_0_1 <= mixColumns_port_state_out_12_0_1;
    roundReg_12_0_2 <= mixColumns_port_state_out_12_0_2;
    roundReg_12_0_3 <= mixColumns_port_state_out_12_0_3;
    roundReg_12_0_4 <= mixColumns_port_state_out_12_0_4;
    roundReg_12_0_5 <= mixColumns_port_state_out_12_0_5;
    roundReg_12_0_6 <= mixColumns_port_state_out_12_0_6;
    roundReg_12_0_7 <= mixColumns_port_state_out_12_0_7;
    roundReg_12_1_0 <= mixColumns_port_state_out_12_1_0;
    roundReg_12_1_1 <= mixColumns_port_state_out_12_1_1;
    roundReg_12_1_2 <= mixColumns_port_state_out_12_1_2;
    roundReg_12_1_3 <= mixColumns_port_state_out_12_1_3;
    roundReg_12_1_4 <= mixColumns_port_state_out_12_1_4;
    roundReg_12_1_5 <= mixColumns_port_state_out_12_1_5;
    roundReg_12_1_6 <= mixColumns_port_state_out_12_1_6;
    roundReg_12_1_7 <= mixColumns_port_state_out_12_1_7;
    roundReg_13_0_0 <= mixColumns_port_state_out_13_0_0;
    roundReg_13_0_1 <= mixColumns_port_state_out_13_0_1;
    roundReg_13_0_2 <= mixColumns_port_state_out_13_0_2;
    roundReg_13_0_3 <= mixColumns_port_state_out_13_0_3;
    roundReg_13_0_4 <= mixColumns_port_state_out_13_0_4;
    roundReg_13_0_5 <= mixColumns_port_state_out_13_0_5;
    roundReg_13_0_6 <= mixColumns_port_state_out_13_0_6;
    roundReg_13_0_7 <= mixColumns_port_state_out_13_0_7;
    roundReg_13_1_0 <= mixColumns_port_state_out_13_1_0;
    roundReg_13_1_1 <= mixColumns_port_state_out_13_1_1;
    roundReg_13_1_2 <= mixColumns_port_state_out_13_1_2;
    roundReg_13_1_3 <= mixColumns_port_state_out_13_1_3;
    roundReg_13_1_4 <= mixColumns_port_state_out_13_1_4;
    roundReg_13_1_5 <= mixColumns_port_state_out_13_1_5;
    roundReg_13_1_6 <= mixColumns_port_state_out_13_1_6;
    roundReg_13_1_7 <= mixColumns_port_state_out_13_1_7;
    roundReg_14_0_0 <= mixColumns_port_state_out_14_0_0;
    roundReg_14_0_1 <= mixColumns_port_state_out_14_0_1;
    roundReg_14_0_2 <= mixColumns_port_state_out_14_0_2;
    roundReg_14_0_3 <= mixColumns_port_state_out_14_0_3;
    roundReg_14_0_4 <= mixColumns_port_state_out_14_0_4;
    roundReg_14_0_5 <= mixColumns_port_state_out_14_0_5;
    roundReg_14_0_6 <= mixColumns_port_state_out_14_0_6;
    roundReg_14_0_7 <= mixColumns_port_state_out_14_0_7;
    roundReg_14_1_0 <= mixColumns_port_state_out_14_1_0;
    roundReg_14_1_1 <= mixColumns_port_state_out_14_1_1;
    roundReg_14_1_2 <= mixColumns_port_state_out_14_1_2;
    roundReg_14_1_3 <= mixColumns_port_state_out_14_1_3;
    roundReg_14_1_4 <= mixColumns_port_state_out_14_1_4;
    roundReg_14_1_5 <= mixColumns_port_state_out_14_1_5;
    roundReg_14_1_6 <= mixColumns_port_state_out_14_1_6;
    roundReg_14_1_7 <= mixColumns_port_state_out_14_1_7;
    roundReg_15_0_0 <= mixColumns_port_state_out_15_0_0;
    roundReg_15_0_1 <= mixColumns_port_state_out_15_0_1;
    roundReg_15_0_2 <= mixColumns_port_state_out_15_0_2;
    roundReg_15_0_3 <= mixColumns_port_state_out_15_0_3;
    roundReg_15_0_4 <= mixColumns_port_state_out_15_0_4;
    roundReg_15_0_5 <= mixColumns_port_state_out_15_0_5;
    roundReg_15_0_6 <= mixColumns_port_state_out_15_0_6;
    roundReg_15_0_7 <= mixColumns_port_state_out_15_0_7;
    roundReg_15_1_0 <= mixColumns_port_state_out_15_1_0;
    roundReg_15_1_1 <= mixColumns_port_state_out_15_1_1;
    roundReg_15_1_2 <= mixColumns_port_state_out_15_1_2;
    roundReg_15_1_3 <= mixColumns_port_state_out_15_1_3;
    roundReg_15_1_4 <= mixColumns_port_state_out_15_1_4;
    roundReg_15_1_5 <= mixColumns_port_state_out_15_1_5;
    roundReg_15_1_6 <= mixColumns_port_state_out_15_1_6;
    roundReg_15_1_7 <= mixColumns_port_state_out_15_1_7;
  end


endmodule

module Aes_MixColumn (
  input      [0:0]    port_state_in_0_0_0,
  input      [0:0]    port_state_in_0_0_1,
  input      [0:0]    port_state_in_0_0_2,
  input      [0:0]    port_state_in_0_0_3,
  input      [0:0]    port_state_in_0_0_4,
  input      [0:0]    port_state_in_0_0_5,
  input      [0:0]    port_state_in_0_0_6,
  input      [0:0]    port_state_in_0_0_7,
  input      [0:0]    port_state_in_0_1_0,
  input      [0:0]    port_state_in_0_1_1,
  input      [0:0]    port_state_in_0_1_2,
  input      [0:0]    port_state_in_0_1_3,
  input      [0:0]    port_state_in_0_1_4,
  input      [0:0]    port_state_in_0_1_5,
  input      [0:0]    port_state_in_0_1_6,
  input      [0:0]    port_state_in_0_1_7,
  input      [0:0]    port_state_in_1_0_0,
  input      [0:0]    port_state_in_1_0_1,
  input      [0:0]    port_state_in_1_0_2,
  input      [0:0]    port_state_in_1_0_3,
  input      [0:0]    port_state_in_1_0_4,
  input      [0:0]    port_state_in_1_0_5,
  input      [0:0]    port_state_in_1_0_6,
  input      [0:0]    port_state_in_1_0_7,
  input      [0:0]    port_state_in_1_1_0,
  input      [0:0]    port_state_in_1_1_1,
  input      [0:0]    port_state_in_1_1_2,
  input      [0:0]    port_state_in_1_1_3,
  input      [0:0]    port_state_in_1_1_4,
  input      [0:0]    port_state_in_1_1_5,
  input      [0:0]    port_state_in_1_1_6,
  input      [0:0]    port_state_in_1_1_7,
  input      [0:0]    port_state_in_2_0_0,
  input      [0:0]    port_state_in_2_0_1,
  input      [0:0]    port_state_in_2_0_2,
  input      [0:0]    port_state_in_2_0_3,
  input      [0:0]    port_state_in_2_0_4,
  input      [0:0]    port_state_in_2_0_5,
  input      [0:0]    port_state_in_2_0_6,
  input      [0:0]    port_state_in_2_0_7,
  input      [0:0]    port_state_in_2_1_0,
  input      [0:0]    port_state_in_2_1_1,
  input      [0:0]    port_state_in_2_1_2,
  input      [0:0]    port_state_in_2_1_3,
  input      [0:0]    port_state_in_2_1_4,
  input      [0:0]    port_state_in_2_1_5,
  input      [0:0]    port_state_in_2_1_6,
  input      [0:0]    port_state_in_2_1_7,
  input      [0:0]    port_state_in_3_0_0,
  input      [0:0]    port_state_in_3_0_1,
  input      [0:0]    port_state_in_3_0_2,
  input      [0:0]    port_state_in_3_0_3,
  input      [0:0]    port_state_in_3_0_4,
  input      [0:0]    port_state_in_3_0_5,
  input      [0:0]    port_state_in_3_0_6,
  input      [0:0]    port_state_in_3_0_7,
  input      [0:0]    port_state_in_3_1_0,
  input      [0:0]    port_state_in_3_1_1,
  input      [0:0]    port_state_in_3_1_2,
  input      [0:0]    port_state_in_3_1_3,
  input      [0:0]    port_state_in_3_1_4,
  input      [0:0]    port_state_in_3_1_5,
  input      [0:0]    port_state_in_3_1_6,
  input      [0:0]    port_state_in_3_1_7,
  input      [0:0]    port_state_in_4_0_0,
  input      [0:0]    port_state_in_4_0_1,
  input      [0:0]    port_state_in_4_0_2,
  input      [0:0]    port_state_in_4_0_3,
  input      [0:0]    port_state_in_4_0_4,
  input      [0:0]    port_state_in_4_0_5,
  input      [0:0]    port_state_in_4_0_6,
  input      [0:0]    port_state_in_4_0_7,
  input      [0:0]    port_state_in_4_1_0,
  input      [0:0]    port_state_in_4_1_1,
  input      [0:0]    port_state_in_4_1_2,
  input      [0:0]    port_state_in_4_1_3,
  input      [0:0]    port_state_in_4_1_4,
  input      [0:0]    port_state_in_4_1_5,
  input      [0:0]    port_state_in_4_1_6,
  input      [0:0]    port_state_in_4_1_7,
  input      [0:0]    port_state_in_5_0_0,
  input      [0:0]    port_state_in_5_0_1,
  input      [0:0]    port_state_in_5_0_2,
  input      [0:0]    port_state_in_5_0_3,
  input      [0:0]    port_state_in_5_0_4,
  input      [0:0]    port_state_in_5_0_5,
  input      [0:0]    port_state_in_5_0_6,
  input      [0:0]    port_state_in_5_0_7,
  input      [0:0]    port_state_in_5_1_0,
  input      [0:0]    port_state_in_5_1_1,
  input      [0:0]    port_state_in_5_1_2,
  input      [0:0]    port_state_in_5_1_3,
  input      [0:0]    port_state_in_5_1_4,
  input      [0:0]    port_state_in_5_1_5,
  input      [0:0]    port_state_in_5_1_6,
  input      [0:0]    port_state_in_5_1_7,
  input      [0:0]    port_state_in_6_0_0,
  input      [0:0]    port_state_in_6_0_1,
  input      [0:0]    port_state_in_6_0_2,
  input      [0:0]    port_state_in_6_0_3,
  input      [0:0]    port_state_in_6_0_4,
  input      [0:0]    port_state_in_6_0_5,
  input      [0:0]    port_state_in_6_0_6,
  input      [0:0]    port_state_in_6_0_7,
  input      [0:0]    port_state_in_6_1_0,
  input      [0:0]    port_state_in_6_1_1,
  input      [0:0]    port_state_in_6_1_2,
  input      [0:0]    port_state_in_6_1_3,
  input      [0:0]    port_state_in_6_1_4,
  input      [0:0]    port_state_in_6_1_5,
  input      [0:0]    port_state_in_6_1_6,
  input      [0:0]    port_state_in_6_1_7,
  input      [0:0]    port_state_in_7_0_0,
  input      [0:0]    port_state_in_7_0_1,
  input      [0:0]    port_state_in_7_0_2,
  input      [0:0]    port_state_in_7_0_3,
  input      [0:0]    port_state_in_7_0_4,
  input      [0:0]    port_state_in_7_0_5,
  input      [0:0]    port_state_in_7_0_6,
  input      [0:0]    port_state_in_7_0_7,
  input      [0:0]    port_state_in_7_1_0,
  input      [0:0]    port_state_in_7_1_1,
  input      [0:0]    port_state_in_7_1_2,
  input      [0:0]    port_state_in_7_1_3,
  input      [0:0]    port_state_in_7_1_4,
  input      [0:0]    port_state_in_7_1_5,
  input      [0:0]    port_state_in_7_1_6,
  input      [0:0]    port_state_in_7_1_7,
  input      [0:0]    port_state_in_8_0_0,
  input      [0:0]    port_state_in_8_0_1,
  input      [0:0]    port_state_in_8_0_2,
  input      [0:0]    port_state_in_8_0_3,
  input      [0:0]    port_state_in_8_0_4,
  input      [0:0]    port_state_in_8_0_5,
  input      [0:0]    port_state_in_8_0_6,
  input      [0:0]    port_state_in_8_0_7,
  input      [0:0]    port_state_in_8_1_0,
  input      [0:0]    port_state_in_8_1_1,
  input      [0:0]    port_state_in_8_1_2,
  input      [0:0]    port_state_in_8_1_3,
  input      [0:0]    port_state_in_8_1_4,
  input      [0:0]    port_state_in_8_1_5,
  input      [0:0]    port_state_in_8_1_6,
  input      [0:0]    port_state_in_8_1_7,
  input      [0:0]    port_state_in_9_0_0,
  input      [0:0]    port_state_in_9_0_1,
  input      [0:0]    port_state_in_9_0_2,
  input      [0:0]    port_state_in_9_0_3,
  input      [0:0]    port_state_in_9_0_4,
  input      [0:0]    port_state_in_9_0_5,
  input      [0:0]    port_state_in_9_0_6,
  input      [0:0]    port_state_in_9_0_7,
  input      [0:0]    port_state_in_9_1_0,
  input      [0:0]    port_state_in_9_1_1,
  input      [0:0]    port_state_in_9_1_2,
  input      [0:0]    port_state_in_9_1_3,
  input      [0:0]    port_state_in_9_1_4,
  input      [0:0]    port_state_in_9_1_5,
  input      [0:0]    port_state_in_9_1_6,
  input      [0:0]    port_state_in_9_1_7,
  input      [0:0]    port_state_in_10_0_0,
  input      [0:0]    port_state_in_10_0_1,
  input      [0:0]    port_state_in_10_0_2,
  input      [0:0]    port_state_in_10_0_3,
  input      [0:0]    port_state_in_10_0_4,
  input      [0:0]    port_state_in_10_0_5,
  input      [0:0]    port_state_in_10_0_6,
  input      [0:0]    port_state_in_10_0_7,
  input      [0:0]    port_state_in_10_1_0,
  input      [0:0]    port_state_in_10_1_1,
  input      [0:0]    port_state_in_10_1_2,
  input      [0:0]    port_state_in_10_1_3,
  input      [0:0]    port_state_in_10_1_4,
  input      [0:0]    port_state_in_10_1_5,
  input      [0:0]    port_state_in_10_1_6,
  input      [0:0]    port_state_in_10_1_7,
  input      [0:0]    port_state_in_11_0_0,
  input      [0:0]    port_state_in_11_0_1,
  input      [0:0]    port_state_in_11_0_2,
  input      [0:0]    port_state_in_11_0_3,
  input      [0:0]    port_state_in_11_0_4,
  input      [0:0]    port_state_in_11_0_5,
  input      [0:0]    port_state_in_11_0_6,
  input      [0:0]    port_state_in_11_0_7,
  input      [0:0]    port_state_in_11_1_0,
  input      [0:0]    port_state_in_11_1_1,
  input      [0:0]    port_state_in_11_1_2,
  input      [0:0]    port_state_in_11_1_3,
  input      [0:0]    port_state_in_11_1_4,
  input      [0:0]    port_state_in_11_1_5,
  input      [0:0]    port_state_in_11_1_6,
  input      [0:0]    port_state_in_11_1_7,
  input      [0:0]    port_state_in_12_0_0,
  input      [0:0]    port_state_in_12_0_1,
  input      [0:0]    port_state_in_12_0_2,
  input      [0:0]    port_state_in_12_0_3,
  input      [0:0]    port_state_in_12_0_4,
  input      [0:0]    port_state_in_12_0_5,
  input      [0:0]    port_state_in_12_0_6,
  input      [0:0]    port_state_in_12_0_7,
  input      [0:0]    port_state_in_12_1_0,
  input      [0:0]    port_state_in_12_1_1,
  input      [0:0]    port_state_in_12_1_2,
  input      [0:0]    port_state_in_12_1_3,
  input      [0:0]    port_state_in_12_1_4,
  input      [0:0]    port_state_in_12_1_5,
  input      [0:0]    port_state_in_12_1_6,
  input      [0:0]    port_state_in_12_1_7,
  input      [0:0]    port_state_in_13_0_0,
  input      [0:0]    port_state_in_13_0_1,
  input      [0:0]    port_state_in_13_0_2,
  input      [0:0]    port_state_in_13_0_3,
  input      [0:0]    port_state_in_13_0_4,
  input      [0:0]    port_state_in_13_0_5,
  input      [0:0]    port_state_in_13_0_6,
  input      [0:0]    port_state_in_13_0_7,
  input      [0:0]    port_state_in_13_1_0,
  input      [0:0]    port_state_in_13_1_1,
  input      [0:0]    port_state_in_13_1_2,
  input      [0:0]    port_state_in_13_1_3,
  input      [0:0]    port_state_in_13_1_4,
  input      [0:0]    port_state_in_13_1_5,
  input      [0:0]    port_state_in_13_1_6,
  input      [0:0]    port_state_in_13_1_7,
  input      [0:0]    port_state_in_14_0_0,
  input      [0:0]    port_state_in_14_0_1,
  input      [0:0]    port_state_in_14_0_2,
  input      [0:0]    port_state_in_14_0_3,
  input      [0:0]    port_state_in_14_0_4,
  input      [0:0]    port_state_in_14_0_5,
  input      [0:0]    port_state_in_14_0_6,
  input      [0:0]    port_state_in_14_0_7,
  input      [0:0]    port_state_in_14_1_0,
  input      [0:0]    port_state_in_14_1_1,
  input      [0:0]    port_state_in_14_1_2,
  input      [0:0]    port_state_in_14_1_3,
  input      [0:0]    port_state_in_14_1_4,
  input      [0:0]    port_state_in_14_1_5,
  input      [0:0]    port_state_in_14_1_6,
  input      [0:0]    port_state_in_14_1_7,
  input      [0:0]    port_state_in_15_0_0,
  input      [0:0]    port_state_in_15_0_1,
  input      [0:0]    port_state_in_15_0_2,
  input      [0:0]    port_state_in_15_0_3,
  input      [0:0]    port_state_in_15_0_4,
  input      [0:0]    port_state_in_15_0_5,
  input      [0:0]    port_state_in_15_0_6,
  input      [0:0]    port_state_in_15_0_7,
  input      [0:0]    port_state_in_15_1_0,
  input      [0:0]    port_state_in_15_1_1,
  input      [0:0]    port_state_in_15_1_2,
  input      [0:0]    port_state_in_15_1_3,
  input      [0:0]    port_state_in_15_1_4,
  input      [0:0]    port_state_in_15_1_5,
  input      [0:0]    port_state_in_15_1_6,
  input      [0:0]    port_state_in_15_1_7,
  output     [0:0]    port_state_out_0_0_0,
  output     [0:0]    port_state_out_0_0_1,
  output     [0:0]    port_state_out_0_0_2,
  output     [0:0]    port_state_out_0_0_3,
  output     [0:0]    port_state_out_0_0_4,
  output     [0:0]    port_state_out_0_0_5,
  output     [0:0]    port_state_out_0_0_6,
  output     [0:0]    port_state_out_0_0_7,
  output     [0:0]    port_state_out_0_1_0,
  output     [0:0]    port_state_out_0_1_1,
  output     [0:0]    port_state_out_0_1_2,
  output     [0:0]    port_state_out_0_1_3,
  output     [0:0]    port_state_out_0_1_4,
  output     [0:0]    port_state_out_0_1_5,
  output     [0:0]    port_state_out_0_1_6,
  output     [0:0]    port_state_out_0_1_7,
  output     [0:0]    port_state_out_1_0_0,
  output     [0:0]    port_state_out_1_0_1,
  output     [0:0]    port_state_out_1_0_2,
  output     [0:0]    port_state_out_1_0_3,
  output     [0:0]    port_state_out_1_0_4,
  output     [0:0]    port_state_out_1_0_5,
  output     [0:0]    port_state_out_1_0_6,
  output     [0:0]    port_state_out_1_0_7,
  output     [0:0]    port_state_out_1_1_0,
  output     [0:0]    port_state_out_1_1_1,
  output     [0:0]    port_state_out_1_1_2,
  output     [0:0]    port_state_out_1_1_3,
  output     [0:0]    port_state_out_1_1_4,
  output     [0:0]    port_state_out_1_1_5,
  output     [0:0]    port_state_out_1_1_6,
  output     [0:0]    port_state_out_1_1_7,
  output     [0:0]    port_state_out_2_0_0,
  output     [0:0]    port_state_out_2_0_1,
  output     [0:0]    port_state_out_2_0_2,
  output     [0:0]    port_state_out_2_0_3,
  output     [0:0]    port_state_out_2_0_4,
  output     [0:0]    port_state_out_2_0_5,
  output     [0:0]    port_state_out_2_0_6,
  output     [0:0]    port_state_out_2_0_7,
  output     [0:0]    port_state_out_2_1_0,
  output     [0:0]    port_state_out_2_1_1,
  output     [0:0]    port_state_out_2_1_2,
  output     [0:0]    port_state_out_2_1_3,
  output     [0:0]    port_state_out_2_1_4,
  output     [0:0]    port_state_out_2_1_5,
  output     [0:0]    port_state_out_2_1_6,
  output     [0:0]    port_state_out_2_1_7,
  output     [0:0]    port_state_out_3_0_0,
  output     [0:0]    port_state_out_3_0_1,
  output     [0:0]    port_state_out_3_0_2,
  output     [0:0]    port_state_out_3_0_3,
  output     [0:0]    port_state_out_3_0_4,
  output     [0:0]    port_state_out_3_0_5,
  output     [0:0]    port_state_out_3_0_6,
  output     [0:0]    port_state_out_3_0_7,
  output     [0:0]    port_state_out_3_1_0,
  output     [0:0]    port_state_out_3_1_1,
  output     [0:0]    port_state_out_3_1_2,
  output     [0:0]    port_state_out_3_1_3,
  output     [0:0]    port_state_out_3_1_4,
  output     [0:0]    port_state_out_3_1_5,
  output     [0:0]    port_state_out_3_1_6,
  output     [0:0]    port_state_out_3_1_7,
  output     [0:0]    port_state_out_4_0_0,
  output     [0:0]    port_state_out_4_0_1,
  output     [0:0]    port_state_out_4_0_2,
  output     [0:0]    port_state_out_4_0_3,
  output     [0:0]    port_state_out_4_0_4,
  output     [0:0]    port_state_out_4_0_5,
  output     [0:0]    port_state_out_4_0_6,
  output     [0:0]    port_state_out_4_0_7,
  output     [0:0]    port_state_out_4_1_0,
  output     [0:0]    port_state_out_4_1_1,
  output     [0:0]    port_state_out_4_1_2,
  output     [0:0]    port_state_out_4_1_3,
  output     [0:0]    port_state_out_4_1_4,
  output     [0:0]    port_state_out_4_1_5,
  output     [0:0]    port_state_out_4_1_6,
  output     [0:0]    port_state_out_4_1_7,
  output     [0:0]    port_state_out_5_0_0,
  output     [0:0]    port_state_out_5_0_1,
  output     [0:0]    port_state_out_5_0_2,
  output     [0:0]    port_state_out_5_0_3,
  output     [0:0]    port_state_out_5_0_4,
  output     [0:0]    port_state_out_5_0_5,
  output     [0:0]    port_state_out_5_0_6,
  output     [0:0]    port_state_out_5_0_7,
  output     [0:0]    port_state_out_5_1_0,
  output     [0:0]    port_state_out_5_1_1,
  output     [0:0]    port_state_out_5_1_2,
  output     [0:0]    port_state_out_5_1_3,
  output     [0:0]    port_state_out_5_1_4,
  output     [0:0]    port_state_out_5_1_5,
  output     [0:0]    port_state_out_5_1_6,
  output     [0:0]    port_state_out_5_1_7,
  output     [0:0]    port_state_out_6_0_0,
  output     [0:0]    port_state_out_6_0_1,
  output     [0:0]    port_state_out_6_0_2,
  output     [0:0]    port_state_out_6_0_3,
  output     [0:0]    port_state_out_6_0_4,
  output     [0:0]    port_state_out_6_0_5,
  output     [0:0]    port_state_out_6_0_6,
  output     [0:0]    port_state_out_6_0_7,
  output     [0:0]    port_state_out_6_1_0,
  output     [0:0]    port_state_out_6_1_1,
  output     [0:0]    port_state_out_6_1_2,
  output     [0:0]    port_state_out_6_1_3,
  output     [0:0]    port_state_out_6_1_4,
  output     [0:0]    port_state_out_6_1_5,
  output     [0:0]    port_state_out_6_1_6,
  output     [0:0]    port_state_out_6_1_7,
  output     [0:0]    port_state_out_7_0_0,
  output     [0:0]    port_state_out_7_0_1,
  output     [0:0]    port_state_out_7_0_2,
  output     [0:0]    port_state_out_7_0_3,
  output     [0:0]    port_state_out_7_0_4,
  output     [0:0]    port_state_out_7_0_5,
  output     [0:0]    port_state_out_7_0_6,
  output     [0:0]    port_state_out_7_0_7,
  output     [0:0]    port_state_out_7_1_0,
  output     [0:0]    port_state_out_7_1_1,
  output     [0:0]    port_state_out_7_1_2,
  output     [0:0]    port_state_out_7_1_3,
  output     [0:0]    port_state_out_7_1_4,
  output     [0:0]    port_state_out_7_1_5,
  output     [0:0]    port_state_out_7_1_6,
  output     [0:0]    port_state_out_7_1_7,
  output     [0:0]    port_state_out_8_0_0,
  output     [0:0]    port_state_out_8_0_1,
  output     [0:0]    port_state_out_8_0_2,
  output     [0:0]    port_state_out_8_0_3,
  output     [0:0]    port_state_out_8_0_4,
  output     [0:0]    port_state_out_8_0_5,
  output     [0:0]    port_state_out_8_0_6,
  output     [0:0]    port_state_out_8_0_7,
  output     [0:0]    port_state_out_8_1_0,
  output     [0:0]    port_state_out_8_1_1,
  output     [0:0]    port_state_out_8_1_2,
  output     [0:0]    port_state_out_8_1_3,
  output     [0:0]    port_state_out_8_1_4,
  output     [0:0]    port_state_out_8_1_5,
  output     [0:0]    port_state_out_8_1_6,
  output     [0:0]    port_state_out_8_1_7,
  output     [0:0]    port_state_out_9_0_0,
  output     [0:0]    port_state_out_9_0_1,
  output     [0:0]    port_state_out_9_0_2,
  output     [0:0]    port_state_out_9_0_3,
  output     [0:0]    port_state_out_9_0_4,
  output     [0:0]    port_state_out_9_0_5,
  output     [0:0]    port_state_out_9_0_6,
  output     [0:0]    port_state_out_9_0_7,
  output     [0:0]    port_state_out_9_1_0,
  output     [0:0]    port_state_out_9_1_1,
  output     [0:0]    port_state_out_9_1_2,
  output     [0:0]    port_state_out_9_1_3,
  output     [0:0]    port_state_out_9_1_4,
  output     [0:0]    port_state_out_9_1_5,
  output     [0:0]    port_state_out_9_1_6,
  output     [0:0]    port_state_out_9_1_7,
  output     [0:0]    port_state_out_10_0_0,
  output     [0:0]    port_state_out_10_0_1,
  output     [0:0]    port_state_out_10_0_2,
  output     [0:0]    port_state_out_10_0_3,
  output     [0:0]    port_state_out_10_0_4,
  output     [0:0]    port_state_out_10_0_5,
  output     [0:0]    port_state_out_10_0_6,
  output     [0:0]    port_state_out_10_0_7,
  output     [0:0]    port_state_out_10_1_0,
  output     [0:0]    port_state_out_10_1_1,
  output     [0:0]    port_state_out_10_1_2,
  output     [0:0]    port_state_out_10_1_3,
  output     [0:0]    port_state_out_10_1_4,
  output     [0:0]    port_state_out_10_1_5,
  output     [0:0]    port_state_out_10_1_6,
  output     [0:0]    port_state_out_10_1_7,
  output     [0:0]    port_state_out_11_0_0,
  output     [0:0]    port_state_out_11_0_1,
  output     [0:0]    port_state_out_11_0_2,
  output     [0:0]    port_state_out_11_0_3,
  output     [0:0]    port_state_out_11_0_4,
  output     [0:0]    port_state_out_11_0_5,
  output     [0:0]    port_state_out_11_0_6,
  output     [0:0]    port_state_out_11_0_7,
  output     [0:0]    port_state_out_11_1_0,
  output     [0:0]    port_state_out_11_1_1,
  output     [0:0]    port_state_out_11_1_2,
  output     [0:0]    port_state_out_11_1_3,
  output     [0:0]    port_state_out_11_1_4,
  output     [0:0]    port_state_out_11_1_5,
  output     [0:0]    port_state_out_11_1_6,
  output     [0:0]    port_state_out_11_1_7,
  output     [0:0]    port_state_out_12_0_0,
  output     [0:0]    port_state_out_12_0_1,
  output     [0:0]    port_state_out_12_0_2,
  output     [0:0]    port_state_out_12_0_3,
  output     [0:0]    port_state_out_12_0_4,
  output     [0:0]    port_state_out_12_0_5,
  output     [0:0]    port_state_out_12_0_6,
  output     [0:0]    port_state_out_12_0_7,
  output     [0:0]    port_state_out_12_1_0,
  output     [0:0]    port_state_out_12_1_1,
  output     [0:0]    port_state_out_12_1_2,
  output     [0:0]    port_state_out_12_1_3,
  output     [0:0]    port_state_out_12_1_4,
  output     [0:0]    port_state_out_12_1_5,
  output     [0:0]    port_state_out_12_1_6,
  output     [0:0]    port_state_out_12_1_7,
  output     [0:0]    port_state_out_13_0_0,
  output     [0:0]    port_state_out_13_0_1,
  output     [0:0]    port_state_out_13_0_2,
  output     [0:0]    port_state_out_13_0_3,
  output     [0:0]    port_state_out_13_0_4,
  output     [0:0]    port_state_out_13_0_5,
  output     [0:0]    port_state_out_13_0_6,
  output     [0:0]    port_state_out_13_0_7,
  output     [0:0]    port_state_out_13_1_0,
  output     [0:0]    port_state_out_13_1_1,
  output     [0:0]    port_state_out_13_1_2,
  output     [0:0]    port_state_out_13_1_3,
  output     [0:0]    port_state_out_13_1_4,
  output     [0:0]    port_state_out_13_1_5,
  output     [0:0]    port_state_out_13_1_6,
  output     [0:0]    port_state_out_13_1_7,
  output     [0:0]    port_state_out_14_0_0,
  output     [0:0]    port_state_out_14_0_1,
  output     [0:0]    port_state_out_14_0_2,
  output     [0:0]    port_state_out_14_0_3,
  output     [0:0]    port_state_out_14_0_4,
  output     [0:0]    port_state_out_14_0_5,
  output     [0:0]    port_state_out_14_0_6,
  output     [0:0]    port_state_out_14_0_7,
  output     [0:0]    port_state_out_14_1_0,
  output     [0:0]    port_state_out_14_1_1,
  output     [0:0]    port_state_out_14_1_2,
  output     [0:0]    port_state_out_14_1_3,
  output     [0:0]    port_state_out_14_1_4,
  output     [0:0]    port_state_out_14_1_5,
  output     [0:0]    port_state_out_14_1_6,
  output     [0:0]    port_state_out_14_1_7,
  output     [0:0]    port_state_out_15_0_0,
  output     [0:0]    port_state_out_15_0_1,
  output     [0:0]    port_state_out_15_0_2,
  output     [0:0]    port_state_out_15_0_3,
  output     [0:0]    port_state_out_15_0_4,
  output     [0:0]    port_state_out_15_0_5,
  output     [0:0]    port_state_out_15_0_6,
  output     [0:0]    port_state_out_15_0_7,
  output     [0:0]    port_state_out_15_1_0,
  output     [0:0]    port_state_out_15_1_1,
  output     [0:0]    port_state_out_15_1_2,
  output     [0:0]    port_state_out_15_1_3,
  output     [0:0]    port_state_out_15_1_4,
  output     [0:0]    port_state_out_15_1_5,
  output     [0:0]    port_state_out_15_1_6,
  output     [0:0]    port_state_out_15_1_7
);

  wire       [0:0]    mul2_32_port_byte_out_0;
  wire       [0:0]    mul2_32_port_byte_out_1;
  wire       [0:0]    mul2_32_port_byte_out_2;
  wire       [0:0]    mul2_32_port_byte_out_3;
  wire       [0:0]    mul2_32_port_byte_out_4;
  wire       [0:0]    mul2_32_port_byte_out_5;
  wire       [0:0]    mul2_32_port_byte_out_6;
  wire       [0:0]    mul2_32_port_byte_out_7;
  wire       [0:0]    mul3_32_port_byte_out_0;
  wire       [0:0]    mul3_32_port_byte_out_1;
  wire       [0:0]    mul3_32_port_byte_out_2;
  wire       [0:0]    mul3_32_port_byte_out_3;
  wire       [0:0]    mul3_32_port_byte_out_4;
  wire       [0:0]    mul3_32_port_byte_out_5;
  wire       [0:0]    mul3_32_port_byte_out_6;
  wire       [0:0]    mul3_32_port_byte_out_7;
  wire       [0:0]    mul2_33_port_byte_out_0;
  wire       [0:0]    mul2_33_port_byte_out_1;
  wire       [0:0]    mul2_33_port_byte_out_2;
  wire       [0:0]    mul2_33_port_byte_out_3;
  wire       [0:0]    mul2_33_port_byte_out_4;
  wire       [0:0]    mul2_33_port_byte_out_5;
  wire       [0:0]    mul2_33_port_byte_out_6;
  wire       [0:0]    mul2_33_port_byte_out_7;
  wire       [0:0]    mul3_33_port_byte_out_0;
  wire       [0:0]    mul3_33_port_byte_out_1;
  wire       [0:0]    mul3_33_port_byte_out_2;
  wire       [0:0]    mul3_33_port_byte_out_3;
  wire       [0:0]    mul3_33_port_byte_out_4;
  wire       [0:0]    mul3_33_port_byte_out_5;
  wire       [0:0]    mul3_33_port_byte_out_6;
  wire       [0:0]    mul3_33_port_byte_out_7;
  wire       [0:0]    mul2_34_port_byte_out_0;
  wire       [0:0]    mul2_34_port_byte_out_1;
  wire       [0:0]    mul2_34_port_byte_out_2;
  wire       [0:0]    mul2_34_port_byte_out_3;
  wire       [0:0]    mul2_34_port_byte_out_4;
  wire       [0:0]    mul2_34_port_byte_out_5;
  wire       [0:0]    mul2_34_port_byte_out_6;
  wire       [0:0]    mul2_34_port_byte_out_7;
  wire       [0:0]    mul3_34_port_byte_out_0;
  wire       [0:0]    mul3_34_port_byte_out_1;
  wire       [0:0]    mul3_34_port_byte_out_2;
  wire       [0:0]    mul3_34_port_byte_out_3;
  wire       [0:0]    mul3_34_port_byte_out_4;
  wire       [0:0]    mul3_34_port_byte_out_5;
  wire       [0:0]    mul3_34_port_byte_out_6;
  wire       [0:0]    mul3_34_port_byte_out_7;
  wire       [0:0]    mul2_35_port_byte_out_0;
  wire       [0:0]    mul2_35_port_byte_out_1;
  wire       [0:0]    mul2_35_port_byte_out_2;
  wire       [0:0]    mul2_35_port_byte_out_3;
  wire       [0:0]    mul2_35_port_byte_out_4;
  wire       [0:0]    mul2_35_port_byte_out_5;
  wire       [0:0]    mul2_35_port_byte_out_6;
  wire       [0:0]    mul2_35_port_byte_out_7;
  wire       [0:0]    mul3_35_port_byte_out_0;
  wire       [0:0]    mul3_35_port_byte_out_1;
  wire       [0:0]    mul3_35_port_byte_out_2;
  wire       [0:0]    mul3_35_port_byte_out_3;
  wire       [0:0]    mul3_35_port_byte_out_4;
  wire       [0:0]    mul3_35_port_byte_out_5;
  wire       [0:0]    mul3_35_port_byte_out_6;
  wire       [0:0]    mul3_35_port_byte_out_7;
  wire       [0:0]    mul2_36_port_byte_out_0;
  wire       [0:0]    mul2_36_port_byte_out_1;
  wire       [0:0]    mul2_36_port_byte_out_2;
  wire       [0:0]    mul2_36_port_byte_out_3;
  wire       [0:0]    mul2_36_port_byte_out_4;
  wire       [0:0]    mul2_36_port_byte_out_5;
  wire       [0:0]    mul2_36_port_byte_out_6;
  wire       [0:0]    mul2_36_port_byte_out_7;
  wire       [0:0]    mul3_36_port_byte_out_0;
  wire       [0:0]    mul3_36_port_byte_out_1;
  wire       [0:0]    mul3_36_port_byte_out_2;
  wire       [0:0]    mul3_36_port_byte_out_3;
  wire       [0:0]    mul3_36_port_byte_out_4;
  wire       [0:0]    mul3_36_port_byte_out_5;
  wire       [0:0]    mul3_36_port_byte_out_6;
  wire       [0:0]    mul3_36_port_byte_out_7;
  wire       [0:0]    mul2_37_port_byte_out_0;
  wire       [0:0]    mul2_37_port_byte_out_1;
  wire       [0:0]    mul2_37_port_byte_out_2;
  wire       [0:0]    mul2_37_port_byte_out_3;
  wire       [0:0]    mul2_37_port_byte_out_4;
  wire       [0:0]    mul2_37_port_byte_out_5;
  wire       [0:0]    mul2_37_port_byte_out_6;
  wire       [0:0]    mul2_37_port_byte_out_7;
  wire       [0:0]    mul3_37_port_byte_out_0;
  wire       [0:0]    mul3_37_port_byte_out_1;
  wire       [0:0]    mul3_37_port_byte_out_2;
  wire       [0:0]    mul3_37_port_byte_out_3;
  wire       [0:0]    mul3_37_port_byte_out_4;
  wire       [0:0]    mul3_37_port_byte_out_5;
  wire       [0:0]    mul3_37_port_byte_out_6;
  wire       [0:0]    mul3_37_port_byte_out_7;
  wire       [0:0]    mul2_38_port_byte_out_0;
  wire       [0:0]    mul2_38_port_byte_out_1;
  wire       [0:0]    mul2_38_port_byte_out_2;
  wire       [0:0]    mul2_38_port_byte_out_3;
  wire       [0:0]    mul2_38_port_byte_out_4;
  wire       [0:0]    mul2_38_port_byte_out_5;
  wire       [0:0]    mul2_38_port_byte_out_6;
  wire       [0:0]    mul2_38_port_byte_out_7;
  wire       [0:0]    mul3_38_port_byte_out_0;
  wire       [0:0]    mul3_38_port_byte_out_1;
  wire       [0:0]    mul3_38_port_byte_out_2;
  wire       [0:0]    mul3_38_port_byte_out_3;
  wire       [0:0]    mul3_38_port_byte_out_4;
  wire       [0:0]    mul3_38_port_byte_out_5;
  wire       [0:0]    mul3_38_port_byte_out_6;
  wire       [0:0]    mul3_38_port_byte_out_7;
  wire       [0:0]    mul2_39_port_byte_out_0;
  wire       [0:0]    mul2_39_port_byte_out_1;
  wire       [0:0]    mul2_39_port_byte_out_2;
  wire       [0:0]    mul2_39_port_byte_out_3;
  wire       [0:0]    mul2_39_port_byte_out_4;
  wire       [0:0]    mul2_39_port_byte_out_5;
  wire       [0:0]    mul2_39_port_byte_out_6;
  wire       [0:0]    mul2_39_port_byte_out_7;
  wire       [0:0]    mul3_39_port_byte_out_0;
  wire       [0:0]    mul3_39_port_byte_out_1;
  wire       [0:0]    mul3_39_port_byte_out_2;
  wire       [0:0]    mul3_39_port_byte_out_3;
  wire       [0:0]    mul3_39_port_byte_out_4;
  wire       [0:0]    mul3_39_port_byte_out_5;
  wire       [0:0]    mul3_39_port_byte_out_6;
  wire       [0:0]    mul3_39_port_byte_out_7;
  wire       [0:0]    mul2_40_port_byte_out_0;
  wire       [0:0]    mul2_40_port_byte_out_1;
  wire       [0:0]    mul2_40_port_byte_out_2;
  wire       [0:0]    mul2_40_port_byte_out_3;
  wire       [0:0]    mul2_40_port_byte_out_4;
  wire       [0:0]    mul2_40_port_byte_out_5;
  wire       [0:0]    mul2_40_port_byte_out_6;
  wire       [0:0]    mul2_40_port_byte_out_7;
  wire       [0:0]    mul3_40_port_byte_out_0;
  wire       [0:0]    mul3_40_port_byte_out_1;
  wire       [0:0]    mul3_40_port_byte_out_2;
  wire       [0:0]    mul3_40_port_byte_out_3;
  wire       [0:0]    mul3_40_port_byte_out_4;
  wire       [0:0]    mul3_40_port_byte_out_5;
  wire       [0:0]    mul3_40_port_byte_out_6;
  wire       [0:0]    mul3_40_port_byte_out_7;
  wire       [0:0]    mul2_41_port_byte_out_0;
  wire       [0:0]    mul2_41_port_byte_out_1;
  wire       [0:0]    mul2_41_port_byte_out_2;
  wire       [0:0]    mul2_41_port_byte_out_3;
  wire       [0:0]    mul2_41_port_byte_out_4;
  wire       [0:0]    mul2_41_port_byte_out_5;
  wire       [0:0]    mul2_41_port_byte_out_6;
  wire       [0:0]    mul2_41_port_byte_out_7;
  wire       [0:0]    mul3_41_port_byte_out_0;
  wire       [0:0]    mul3_41_port_byte_out_1;
  wire       [0:0]    mul3_41_port_byte_out_2;
  wire       [0:0]    mul3_41_port_byte_out_3;
  wire       [0:0]    mul3_41_port_byte_out_4;
  wire       [0:0]    mul3_41_port_byte_out_5;
  wire       [0:0]    mul3_41_port_byte_out_6;
  wire       [0:0]    mul3_41_port_byte_out_7;
  wire       [0:0]    mul2_42_port_byte_out_0;
  wire       [0:0]    mul2_42_port_byte_out_1;
  wire       [0:0]    mul2_42_port_byte_out_2;
  wire       [0:0]    mul2_42_port_byte_out_3;
  wire       [0:0]    mul2_42_port_byte_out_4;
  wire       [0:0]    mul2_42_port_byte_out_5;
  wire       [0:0]    mul2_42_port_byte_out_6;
  wire       [0:0]    mul2_42_port_byte_out_7;
  wire       [0:0]    mul3_42_port_byte_out_0;
  wire       [0:0]    mul3_42_port_byte_out_1;
  wire       [0:0]    mul3_42_port_byte_out_2;
  wire       [0:0]    mul3_42_port_byte_out_3;
  wire       [0:0]    mul3_42_port_byte_out_4;
  wire       [0:0]    mul3_42_port_byte_out_5;
  wire       [0:0]    mul3_42_port_byte_out_6;
  wire       [0:0]    mul3_42_port_byte_out_7;
  wire       [0:0]    mul2_43_port_byte_out_0;
  wire       [0:0]    mul2_43_port_byte_out_1;
  wire       [0:0]    mul2_43_port_byte_out_2;
  wire       [0:0]    mul2_43_port_byte_out_3;
  wire       [0:0]    mul2_43_port_byte_out_4;
  wire       [0:0]    mul2_43_port_byte_out_5;
  wire       [0:0]    mul2_43_port_byte_out_6;
  wire       [0:0]    mul2_43_port_byte_out_7;
  wire       [0:0]    mul3_43_port_byte_out_0;
  wire       [0:0]    mul3_43_port_byte_out_1;
  wire       [0:0]    mul3_43_port_byte_out_2;
  wire       [0:0]    mul3_43_port_byte_out_3;
  wire       [0:0]    mul3_43_port_byte_out_4;
  wire       [0:0]    mul3_43_port_byte_out_5;
  wire       [0:0]    mul3_43_port_byte_out_6;
  wire       [0:0]    mul3_43_port_byte_out_7;
  wire       [0:0]    mul2_44_port_byte_out_0;
  wire       [0:0]    mul2_44_port_byte_out_1;
  wire       [0:0]    mul2_44_port_byte_out_2;
  wire       [0:0]    mul2_44_port_byte_out_3;
  wire       [0:0]    mul2_44_port_byte_out_4;
  wire       [0:0]    mul2_44_port_byte_out_5;
  wire       [0:0]    mul2_44_port_byte_out_6;
  wire       [0:0]    mul2_44_port_byte_out_7;
  wire       [0:0]    mul3_44_port_byte_out_0;
  wire       [0:0]    mul3_44_port_byte_out_1;
  wire       [0:0]    mul3_44_port_byte_out_2;
  wire       [0:0]    mul3_44_port_byte_out_3;
  wire       [0:0]    mul3_44_port_byte_out_4;
  wire       [0:0]    mul3_44_port_byte_out_5;
  wire       [0:0]    mul3_44_port_byte_out_6;
  wire       [0:0]    mul3_44_port_byte_out_7;
  wire       [0:0]    mul2_45_port_byte_out_0;
  wire       [0:0]    mul2_45_port_byte_out_1;
  wire       [0:0]    mul2_45_port_byte_out_2;
  wire       [0:0]    mul2_45_port_byte_out_3;
  wire       [0:0]    mul2_45_port_byte_out_4;
  wire       [0:0]    mul2_45_port_byte_out_5;
  wire       [0:0]    mul2_45_port_byte_out_6;
  wire       [0:0]    mul2_45_port_byte_out_7;
  wire       [0:0]    mul3_45_port_byte_out_0;
  wire       [0:0]    mul3_45_port_byte_out_1;
  wire       [0:0]    mul3_45_port_byte_out_2;
  wire       [0:0]    mul3_45_port_byte_out_3;
  wire       [0:0]    mul3_45_port_byte_out_4;
  wire       [0:0]    mul3_45_port_byte_out_5;
  wire       [0:0]    mul3_45_port_byte_out_6;
  wire       [0:0]    mul3_45_port_byte_out_7;
  wire       [0:0]    mul2_46_port_byte_out_0;
  wire       [0:0]    mul2_46_port_byte_out_1;
  wire       [0:0]    mul2_46_port_byte_out_2;
  wire       [0:0]    mul2_46_port_byte_out_3;
  wire       [0:0]    mul2_46_port_byte_out_4;
  wire       [0:0]    mul2_46_port_byte_out_5;
  wire       [0:0]    mul2_46_port_byte_out_6;
  wire       [0:0]    mul2_46_port_byte_out_7;
  wire       [0:0]    mul3_46_port_byte_out_0;
  wire       [0:0]    mul3_46_port_byte_out_1;
  wire       [0:0]    mul3_46_port_byte_out_2;
  wire       [0:0]    mul3_46_port_byte_out_3;
  wire       [0:0]    mul3_46_port_byte_out_4;
  wire       [0:0]    mul3_46_port_byte_out_5;
  wire       [0:0]    mul3_46_port_byte_out_6;
  wire       [0:0]    mul3_46_port_byte_out_7;
  wire       [0:0]    mul2_47_port_byte_out_0;
  wire       [0:0]    mul2_47_port_byte_out_1;
  wire       [0:0]    mul2_47_port_byte_out_2;
  wire       [0:0]    mul2_47_port_byte_out_3;
  wire       [0:0]    mul2_47_port_byte_out_4;
  wire       [0:0]    mul2_47_port_byte_out_5;
  wire       [0:0]    mul2_47_port_byte_out_6;
  wire       [0:0]    mul2_47_port_byte_out_7;
  wire       [0:0]    mul3_47_port_byte_out_0;
  wire       [0:0]    mul3_47_port_byte_out_1;
  wire       [0:0]    mul3_47_port_byte_out_2;
  wire       [0:0]    mul3_47_port_byte_out_3;
  wire       [0:0]    mul3_47_port_byte_out_4;
  wire       [0:0]    mul3_47_port_byte_out_5;
  wire       [0:0]    mul3_47_port_byte_out_6;
  wire       [0:0]    mul3_47_port_byte_out_7;
  wire       [0:0]    mul2_48_port_byte_out_0;
  wire       [0:0]    mul2_48_port_byte_out_1;
  wire       [0:0]    mul2_48_port_byte_out_2;
  wire       [0:0]    mul2_48_port_byte_out_3;
  wire       [0:0]    mul2_48_port_byte_out_4;
  wire       [0:0]    mul2_48_port_byte_out_5;
  wire       [0:0]    mul2_48_port_byte_out_6;
  wire       [0:0]    mul2_48_port_byte_out_7;
  wire       [0:0]    mul3_48_port_byte_out_0;
  wire       [0:0]    mul3_48_port_byte_out_1;
  wire       [0:0]    mul3_48_port_byte_out_2;
  wire       [0:0]    mul3_48_port_byte_out_3;
  wire       [0:0]    mul3_48_port_byte_out_4;
  wire       [0:0]    mul3_48_port_byte_out_5;
  wire       [0:0]    mul3_48_port_byte_out_6;
  wire       [0:0]    mul3_48_port_byte_out_7;
  wire       [0:0]    mul2_49_port_byte_out_0;
  wire       [0:0]    mul2_49_port_byte_out_1;
  wire       [0:0]    mul2_49_port_byte_out_2;
  wire       [0:0]    mul2_49_port_byte_out_3;
  wire       [0:0]    mul2_49_port_byte_out_4;
  wire       [0:0]    mul2_49_port_byte_out_5;
  wire       [0:0]    mul2_49_port_byte_out_6;
  wire       [0:0]    mul2_49_port_byte_out_7;
  wire       [0:0]    mul3_49_port_byte_out_0;
  wire       [0:0]    mul3_49_port_byte_out_1;
  wire       [0:0]    mul3_49_port_byte_out_2;
  wire       [0:0]    mul3_49_port_byte_out_3;
  wire       [0:0]    mul3_49_port_byte_out_4;
  wire       [0:0]    mul3_49_port_byte_out_5;
  wire       [0:0]    mul3_49_port_byte_out_6;
  wire       [0:0]    mul3_49_port_byte_out_7;
  wire       [0:0]    mul2_50_port_byte_out_0;
  wire       [0:0]    mul2_50_port_byte_out_1;
  wire       [0:0]    mul2_50_port_byte_out_2;
  wire       [0:0]    mul2_50_port_byte_out_3;
  wire       [0:0]    mul2_50_port_byte_out_4;
  wire       [0:0]    mul2_50_port_byte_out_5;
  wire       [0:0]    mul2_50_port_byte_out_6;
  wire       [0:0]    mul2_50_port_byte_out_7;
  wire       [0:0]    mul3_50_port_byte_out_0;
  wire       [0:0]    mul3_50_port_byte_out_1;
  wire       [0:0]    mul3_50_port_byte_out_2;
  wire       [0:0]    mul3_50_port_byte_out_3;
  wire       [0:0]    mul3_50_port_byte_out_4;
  wire       [0:0]    mul3_50_port_byte_out_5;
  wire       [0:0]    mul3_50_port_byte_out_6;
  wire       [0:0]    mul3_50_port_byte_out_7;
  wire       [0:0]    mul2_51_port_byte_out_0;
  wire       [0:0]    mul2_51_port_byte_out_1;
  wire       [0:0]    mul2_51_port_byte_out_2;
  wire       [0:0]    mul2_51_port_byte_out_3;
  wire       [0:0]    mul2_51_port_byte_out_4;
  wire       [0:0]    mul2_51_port_byte_out_5;
  wire       [0:0]    mul2_51_port_byte_out_6;
  wire       [0:0]    mul2_51_port_byte_out_7;
  wire       [0:0]    mul3_51_port_byte_out_0;
  wire       [0:0]    mul3_51_port_byte_out_1;
  wire       [0:0]    mul3_51_port_byte_out_2;
  wire       [0:0]    mul3_51_port_byte_out_3;
  wire       [0:0]    mul3_51_port_byte_out_4;
  wire       [0:0]    mul3_51_port_byte_out_5;
  wire       [0:0]    mul3_51_port_byte_out_6;
  wire       [0:0]    mul3_51_port_byte_out_7;
  wire       [0:0]    mul2_52_port_byte_out_0;
  wire       [0:0]    mul2_52_port_byte_out_1;
  wire       [0:0]    mul2_52_port_byte_out_2;
  wire       [0:0]    mul2_52_port_byte_out_3;
  wire       [0:0]    mul2_52_port_byte_out_4;
  wire       [0:0]    mul2_52_port_byte_out_5;
  wire       [0:0]    mul2_52_port_byte_out_6;
  wire       [0:0]    mul2_52_port_byte_out_7;
  wire       [0:0]    mul3_52_port_byte_out_0;
  wire       [0:0]    mul3_52_port_byte_out_1;
  wire       [0:0]    mul3_52_port_byte_out_2;
  wire       [0:0]    mul3_52_port_byte_out_3;
  wire       [0:0]    mul3_52_port_byte_out_4;
  wire       [0:0]    mul3_52_port_byte_out_5;
  wire       [0:0]    mul3_52_port_byte_out_6;
  wire       [0:0]    mul3_52_port_byte_out_7;
  wire       [0:0]    mul2_53_port_byte_out_0;
  wire       [0:0]    mul2_53_port_byte_out_1;
  wire       [0:0]    mul2_53_port_byte_out_2;
  wire       [0:0]    mul2_53_port_byte_out_3;
  wire       [0:0]    mul2_53_port_byte_out_4;
  wire       [0:0]    mul2_53_port_byte_out_5;
  wire       [0:0]    mul2_53_port_byte_out_6;
  wire       [0:0]    mul2_53_port_byte_out_7;
  wire       [0:0]    mul3_53_port_byte_out_0;
  wire       [0:0]    mul3_53_port_byte_out_1;
  wire       [0:0]    mul3_53_port_byte_out_2;
  wire       [0:0]    mul3_53_port_byte_out_3;
  wire       [0:0]    mul3_53_port_byte_out_4;
  wire       [0:0]    mul3_53_port_byte_out_5;
  wire       [0:0]    mul3_53_port_byte_out_6;
  wire       [0:0]    mul3_53_port_byte_out_7;
  wire       [0:0]    mul2_54_port_byte_out_0;
  wire       [0:0]    mul2_54_port_byte_out_1;
  wire       [0:0]    mul2_54_port_byte_out_2;
  wire       [0:0]    mul2_54_port_byte_out_3;
  wire       [0:0]    mul2_54_port_byte_out_4;
  wire       [0:0]    mul2_54_port_byte_out_5;
  wire       [0:0]    mul2_54_port_byte_out_6;
  wire       [0:0]    mul2_54_port_byte_out_7;
  wire       [0:0]    mul3_54_port_byte_out_0;
  wire       [0:0]    mul3_54_port_byte_out_1;
  wire       [0:0]    mul3_54_port_byte_out_2;
  wire       [0:0]    mul3_54_port_byte_out_3;
  wire       [0:0]    mul3_54_port_byte_out_4;
  wire       [0:0]    mul3_54_port_byte_out_5;
  wire       [0:0]    mul3_54_port_byte_out_6;
  wire       [0:0]    mul3_54_port_byte_out_7;
  wire       [0:0]    mul2_55_port_byte_out_0;
  wire       [0:0]    mul2_55_port_byte_out_1;
  wire       [0:0]    mul2_55_port_byte_out_2;
  wire       [0:0]    mul2_55_port_byte_out_3;
  wire       [0:0]    mul2_55_port_byte_out_4;
  wire       [0:0]    mul2_55_port_byte_out_5;
  wire       [0:0]    mul2_55_port_byte_out_6;
  wire       [0:0]    mul2_55_port_byte_out_7;
  wire       [0:0]    mul3_55_port_byte_out_0;
  wire       [0:0]    mul3_55_port_byte_out_1;
  wire       [0:0]    mul3_55_port_byte_out_2;
  wire       [0:0]    mul3_55_port_byte_out_3;
  wire       [0:0]    mul3_55_port_byte_out_4;
  wire       [0:0]    mul3_55_port_byte_out_5;
  wire       [0:0]    mul3_55_port_byte_out_6;
  wire       [0:0]    mul3_55_port_byte_out_7;
  wire       [0:0]    mul2_56_port_byte_out_0;
  wire       [0:0]    mul2_56_port_byte_out_1;
  wire       [0:0]    mul2_56_port_byte_out_2;
  wire       [0:0]    mul2_56_port_byte_out_3;
  wire       [0:0]    mul2_56_port_byte_out_4;
  wire       [0:0]    mul2_56_port_byte_out_5;
  wire       [0:0]    mul2_56_port_byte_out_6;
  wire       [0:0]    mul2_56_port_byte_out_7;
  wire       [0:0]    mul3_56_port_byte_out_0;
  wire       [0:0]    mul3_56_port_byte_out_1;
  wire       [0:0]    mul3_56_port_byte_out_2;
  wire       [0:0]    mul3_56_port_byte_out_3;
  wire       [0:0]    mul3_56_port_byte_out_4;
  wire       [0:0]    mul3_56_port_byte_out_5;
  wire       [0:0]    mul3_56_port_byte_out_6;
  wire       [0:0]    mul3_56_port_byte_out_7;
  wire       [0:0]    mul2_57_port_byte_out_0;
  wire       [0:0]    mul2_57_port_byte_out_1;
  wire       [0:0]    mul2_57_port_byte_out_2;
  wire       [0:0]    mul2_57_port_byte_out_3;
  wire       [0:0]    mul2_57_port_byte_out_4;
  wire       [0:0]    mul2_57_port_byte_out_5;
  wire       [0:0]    mul2_57_port_byte_out_6;
  wire       [0:0]    mul2_57_port_byte_out_7;
  wire       [0:0]    mul3_57_port_byte_out_0;
  wire       [0:0]    mul3_57_port_byte_out_1;
  wire       [0:0]    mul3_57_port_byte_out_2;
  wire       [0:0]    mul3_57_port_byte_out_3;
  wire       [0:0]    mul3_57_port_byte_out_4;
  wire       [0:0]    mul3_57_port_byte_out_5;
  wire       [0:0]    mul3_57_port_byte_out_6;
  wire       [0:0]    mul3_57_port_byte_out_7;
  wire       [0:0]    mul2_58_port_byte_out_0;
  wire       [0:0]    mul2_58_port_byte_out_1;
  wire       [0:0]    mul2_58_port_byte_out_2;
  wire       [0:0]    mul2_58_port_byte_out_3;
  wire       [0:0]    mul2_58_port_byte_out_4;
  wire       [0:0]    mul2_58_port_byte_out_5;
  wire       [0:0]    mul2_58_port_byte_out_6;
  wire       [0:0]    mul2_58_port_byte_out_7;
  wire       [0:0]    mul3_58_port_byte_out_0;
  wire       [0:0]    mul3_58_port_byte_out_1;
  wire       [0:0]    mul3_58_port_byte_out_2;
  wire       [0:0]    mul3_58_port_byte_out_3;
  wire       [0:0]    mul3_58_port_byte_out_4;
  wire       [0:0]    mul3_58_port_byte_out_5;
  wire       [0:0]    mul3_58_port_byte_out_6;
  wire       [0:0]    mul3_58_port_byte_out_7;
  wire       [0:0]    mul2_59_port_byte_out_0;
  wire       [0:0]    mul2_59_port_byte_out_1;
  wire       [0:0]    mul2_59_port_byte_out_2;
  wire       [0:0]    mul2_59_port_byte_out_3;
  wire       [0:0]    mul2_59_port_byte_out_4;
  wire       [0:0]    mul2_59_port_byte_out_5;
  wire       [0:0]    mul2_59_port_byte_out_6;
  wire       [0:0]    mul2_59_port_byte_out_7;
  wire       [0:0]    mul3_59_port_byte_out_0;
  wire       [0:0]    mul3_59_port_byte_out_1;
  wire       [0:0]    mul3_59_port_byte_out_2;
  wire       [0:0]    mul3_59_port_byte_out_3;
  wire       [0:0]    mul3_59_port_byte_out_4;
  wire       [0:0]    mul3_59_port_byte_out_5;
  wire       [0:0]    mul3_59_port_byte_out_6;
  wire       [0:0]    mul3_59_port_byte_out_7;
  wire       [0:0]    mul2_60_port_byte_out_0;
  wire       [0:0]    mul2_60_port_byte_out_1;
  wire       [0:0]    mul2_60_port_byte_out_2;
  wire       [0:0]    mul2_60_port_byte_out_3;
  wire       [0:0]    mul2_60_port_byte_out_4;
  wire       [0:0]    mul2_60_port_byte_out_5;
  wire       [0:0]    mul2_60_port_byte_out_6;
  wire       [0:0]    mul2_60_port_byte_out_7;
  wire       [0:0]    mul3_60_port_byte_out_0;
  wire       [0:0]    mul3_60_port_byte_out_1;
  wire       [0:0]    mul3_60_port_byte_out_2;
  wire       [0:0]    mul3_60_port_byte_out_3;
  wire       [0:0]    mul3_60_port_byte_out_4;
  wire       [0:0]    mul3_60_port_byte_out_5;
  wire       [0:0]    mul3_60_port_byte_out_6;
  wire       [0:0]    mul3_60_port_byte_out_7;
  wire       [0:0]    mul2_61_port_byte_out_0;
  wire       [0:0]    mul2_61_port_byte_out_1;
  wire       [0:0]    mul2_61_port_byte_out_2;
  wire       [0:0]    mul2_61_port_byte_out_3;
  wire       [0:0]    mul2_61_port_byte_out_4;
  wire       [0:0]    mul2_61_port_byte_out_5;
  wire       [0:0]    mul2_61_port_byte_out_6;
  wire       [0:0]    mul2_61_port_byte_out_7;
  wire       [0:0]    mul3_61_port_byte_out_0;
  wire       [0:0]    mul3_61_port_byte_out_1;
  wire       [0:0]    mul3_61_port_byte_out_2;
  wire       [0:0]    mul3_61_port_byte_out_3;
  wire       [0:0]    mul3_61_port_byte_out_4;
  wire       [0:0]    mul3_61_port_byte_out_5;
  wire       [0:0]    mul3_61_port_byte_out_6;
  wire       [0:0]    mul3_61_port_byte_out_7;
  wire       [0:0]    mul2_62_port_byte_out_0;
  wire       [0:0]    mul2_62_port_byte_out_1;
  wire       [0:0]    mul2_62_port_byte_out_2;
  wire       [0:0]    mul2_62_port_byte_out_3;
  wire       [0:0]    mul2_62_port_byte_out_4;
  wire       [0:0]    mul2_62_port_byte_out_5;
  wire       [0:0]    mul2_62_port_byte_out_6;
  wire       [0:0]    mul2_62_port_byte_out_7;
  wire       [0:0]    mul3_62_port_byte_out_0;
  wire       [0:0]    mul3_62_port_byte_out_1;
  wire       [0:0]    mul3_62_port_byte_out_2;
  wire       [0:0]    mul3_62_port_byte_out_3;
  wire       [0:0]    mul3_62_port_byte_out_4;
  wire       [0:0]    mul3_62_port_byte_out_5;
  wire       [0:0]    mul3_62_port_byte_out_6;
  wire       [0:0]    mul3_62_port_byte_out_7;
  wire       [0:0]    mul2_63_port_byte_out_0;
  wire       [0:0]    mul2_63_port_byte_out_1;
  wire       [0:0]    mul2_63_port_byte_out_2;
  wire       [0:0]    mul2_63_port_byte_out_3;
  wire       [0:0]    mul2_63_port_byte_out_4;
  wire       [0:0]    mul2_63_port_byte_out_5;
  wire       [0:0]    mul2_63_port_byte_out_6;
  wire       [0:0]    mul2_63_port_byte_out_7;
  wire       [0:0]    mul3_63_port_byte_out_0;
  wire       [0:0]    mul3_63_port_byte_out_1;
  wire       [0:0]    mul3_63_port_byte_out_2;
  wire       [0:0]    mul3_63_port_byte_out_3;
  wire       [0:0]    mul3_63_port_byte_out_4;
  wire       [0:0]    mul3_63_port_byte_out_5;
  wire       [0:0]    mul3_63_port_byte_out_6;
  wire       [0:0]    mul3_63_port_byte_out_7;
  wire       [0:0]    state_out_0_0_0;
  wire       [0:0]    state_out_0_0_1;
  wire       [0:0]    state_out_0_0_2;
  wire       [0:0]    state_out_0_0_3;
  wire       [0:0]    state_out_0_0_4;
  wire       [0:0]    state_out_0_0_5;
  wire       [0:0]    state_out_0_0_6;
  wire       [0:0]    state_out_0_0_7;
  wire       [0:0]    state_out_0_1_0;
  wire       [0:0]    state_out_0_1_1;
  wire       [0:0]    state_out_0_1_2;
  wire       [0:0]    state_out_0_1_3;
  wire       [0:0]    state_out_0_1_4;
  wire       [0:0]    state_out_0_1_5;
  wire       [0:0]    state_out_0_1_6;
  wire       [0:0]    state_out_0_1_7;
  wire       [0:0]    state_out_1_0_0;
  wire       [0:0]    state_out_1_0_1;
  wire       [0:0]    state_out_1_0_2;
  wire       [0:0]    state_out_1_0_3;
  wire       [0:0]    state_out_1_0_4;
  wire       [0:0]    state_out_1_0_5;
  wire       [0:0]    state_out_1_0_6;
  wire       [0:0]    state_out_1_0_7;
  wire       [0:0]    state_out_1_1_0;
  wire       [0:0]    state_out_1_1_1;
  wire       [0:0]    state_out_1_1_2;
  wire       [0:0]    state_out_1_1_3;
  wire       [0:0]    state_out_1_1_4;
  wire       [0:0]    state_out_1_1_5;
  wire       [0:0]    state_out_1_1_6;
  wire       [0:0]    state_out_1_1_7;
  wire       [0:0]    state_out_2_0_0;
  wire       [0:0]    state_out_2_0_1;
  wire       [0:0]    state_out_2_0_2;
  wire       [0:0]    state_out_2_0_3;
  wire       [0:0]    state_out_2_0_4;
  wire       [0:0]    state_out_2_0_5;
  wire       [0:0]    state_out_2_0_6;
  wire       [0:0]    state_out_2_0_7;
  wire       [0:0]    state_out_2_1_0;
  wire       [0:0]    state_out_2_1_1;
  wire       [0:0]    state_out_2_1_2;
  wire       [0:0]    state_out_2_1_3;
  wire       [0:0]    state_out_2_1_4;
  wire       [0:0]    state_out_2_1_5;
  wire       [0:0]    state_out_2_1_6;
  wire       [0:0]    state_out_2_1_7;
  wire       [0:0]    state_out_3_0_0;
  wire       [0:0]    state_out_3_0_1;
  wire       [0:0]    state_out_3_0_2;
  wire       [0:0]    state_out_3_0_3;
  wire       [0:0]    state_out_3_0_4;
  wire       [0:0]    state_out_3_0_5;
  wire       [0:0]    state_out_3_0_6;
  wire       [0:0]    state_out_3_0_7;
  wire       [0:0]    state_out_3_1_0;
  wire       [0:0]    state_out_3_1_1;
  wire       [0:0]    state_out_3_1_2;
  wire       [0:0]    state_out_3_1_3;
  wire       [0:0]    state_out_3_1_4;
  wire       [0:0]    state_out_3_1_5;
  wire       [0:0]    state_out_3_1_6;
  wire       [0:0]    state_out_3_1_7;
  wire       [0:0]    state_out_4_0_0;
  wire       [0:0]    state_out_4_0_1;
  wire       [0:0]    state_out_4_0_2;
  wire       [0:0]    state_out_4_0_3;
  wire       [0:0]    state_out_4_0_4;
  wire       [0:0]    state_out_4_0_5;
  wire       [0:0]    state_out_4_0_6;
  wire       [0:0]    state_out_4_0_7;
  wire       [0:0]    state_out_4_1_0;
  wire       [0:0]    state_out_4_1_1;
  wire       [0:0]    state_out_4_1_2;
  wire       [0:0]    state_out_4_1_3;
  wire       [0:0]    state_out_4_1_4;
  wire       [0:0]    state_out_4_1_5;
  wire       [0:0]    state_out_4_1_6;
  wire       [0:0]    state_out_4_1_7;
  wire       [0:0]    state_out_5_0_0;
  wire       [0:0]    state_out_5_0_1;
  wire       [0:0]    state_out_5_0_2;
  wire       [0:0]    state_out_5_0_3;
  wire       [0:0]    state_out_5_0_4;
  wire       [0:0]    state_out_5_0_5;
  wire       [0:0]    state_out_5_0_6;
  wire       [0:0]    state_out_5_0_7;
  wire       [0:0]    state_out_5_1_0;
  wire       [0:0]    state_out_5_1_1;
  wire       [0:0]    state_out_5_1_2;
  wire       [0:0]    state_out_5_1_3;
  wire       [0:0]    state_out_5_1_4;
  wire       [0:0]    state_out_5_1_5;
  wire       [0:0]    state_out_5_1_6;
  wire       [0:0]    state_out_5_1_7;
  wire       [0:0]    state_out_6_0_0;
  wire       [0:0]    state_out_6_0_1;
  wire       [0:0]    state_out_6_0_2;
  wire       [0:0]    state_out_6_0_3;
  wire       [0:0]    state_out_6_0_4;
  wire       [0:0]    state_out_6_0_5;
  wire       [0:0]    state_out_6_0_6;
  wire       [0:0]    state_out_6_0_7;
  wire       [0:0]    state_out_6_1_0;
  wire       [0:0]    state_out_6_1_1;
  wire       [0:0]    state_out_6_1_2;
  wire       [0:0]    state_out_6_1_3;
  wire       [0:0]    state_out_6_1_4;
  wire       [0:0]    state_out_6_1_5;
  wire       [0:0]    state_out_6_1_6;
  wire       [0:0]    state_out_6_1_7;
  wire       [0:0]    state_out_7_0_0;
  wire       [0:0]    state_out_7_0_1;
  wire       [0:0]    state_out_7_0_2;
  wire       [0:0]    state_out_7_0_3;
  wire       [0:0]    state_out_7_0_4;
  wire       [0:0]    state_out_7_0_5;
  wire       [0:0]    state_out_7_0_6;
  wire       [0:0]    state_out_7_0_7;
  wire       [0:0]    state_out_7_1_0;
  wire       [0:0]    state_out_7_1_1;
  wire       [0:0]    state_out_7_1_2;
  wire       [0:0]    state_out_7_1_3;
  wire       [0:0]    state_out_7_1_4;
  wire       [0:0]    state_out_7_1_5;
  wire       [0:0]    state_out_7_1_6;
  wire       [0:0]    state_out_7_1_7;
  wire       [0:0]    state_out_8_0_0;
  wire       [0:0]    state_out_8_0_1;
  wire       [0:0]    state_out_8_0_2;
  wire       [0:0]    state_out_8_0_3;
  wire       [0:0]    state_out_8_0_4;
  wire       [0:0]    state_out_8_0_5;
  wire       [0:0]    state_out_8_0_6;
  wire       [0:0]    state_out_8_0_7;
  wire       [0:0]    state_out_8_1_0;
  wire       [0:0]    state_out_8_1_1;
  wire       [0:0]    state_out_8_1_2;
  wire       [0:0]    state_out_8_1_3;
  wire       [0:0]    state_out_8_1_4;
  wire       [0:0]    state_out_8_1_5;
  wire       [0:0]    state_out_8_1_6;
  wire       [0:0]    state_out_8_1_7;
  wire       [0:0]    state_out_9_0_0;
  wire       [0:0]    state_out_9_0_1;
  wire       [0:0]    state_out_9_0_2;
  wire       [0:0]    state_out_9_0_3;
  wire       [0:0]    state_out_9_0_4;
  wire       [0:0]    state_out_9_0_5;
  wire       [0:0]    state_out_9_0_6;
  wire       [0:0]    state_out_9_0_7;
  wire       [0:0]    state_out_9_1_0;
  wire       [0:0]    state_out_9_1_1;
  wire       [0:0]    state_out_9_1_2;
  wire       [0:0]    state_out_9_1_3;
  wire       [0:0]    state_out_9_1_4;
  wire       [0:0]    state_out_9_1_5;
  wire       [0:0]    state_out_9_1_6;
  wire       [0:0]    state_out_9_1_7;
  wire       [0:0]    state_out_10_0_0;
  wire       [0:0]    state_out_10_0_1;
  wire       [0:0]    state_out_10_0_2;
  wire       [0:0]    state_out_10_0_3;
  wire       [0:0]    state_out_10_0_4;
  wire       [0:0]    state_out_10_0_5;
  wire       [0:0]    state_out_10_0_6;
  wire       [0:0]    state_out_10_0_7;
  wire       [0:0]    state_out_10_1_0;
  wire       [0:0]    state_out_10_1_1;
  wire       [0:0]    state_out_10_1_2;
  wire       [0:0]    state_out_10_1_3;
  wire       [0:0]    state_out_10_1_4;
  wire       [0:0]    state_out_10_1_5;
  wire       [0:0]    state_out_10_1_6;
  wire       [0:0]    state_out_10_1_7;
  wire       [0:0]    state_out_11_0_0;
  wire       [0:0]    state_out_11_0_1;
  wire       [0:0]    state_out_11_0_2;
  wire       [0:0]    state_out_11_0_3;
  wire       [0:0]    state_out_11_0_4;
  wire       [0:0]    state_out_11_0_5;
  wire       [0:0]    state_out_11_0_6;
  wire       [0:0]    state_out_11_0_7;
  wire       [0:0]    state_out_11_1_0;
  wire       [0:0]    state_out_11_1_1;
  wire       [0:0]    state_out_11_1_2;
  wire       [0:0]    state_out_11_1_3;
  wire       [0:0]    state_out_11_1_4;
  wire       [0:0]    state_out_11_1_5;
  wire       [0:0]    state_out_11_1_6;
  wire       [0:0]    state_out_11_1_7;
  wire       [0:0]    state_out_12_0_0;
  wire       [0:0]    state_out_12_0_1;
  wire       [0:0]    state_out_12_0_2;
  wire       [0:0]    state_out_12_0_3;
  wire       [0:0]    state_out_12_0_4;
  wire       [0:0]    state_out_12_0_5;
  wire       [0:0]    state_out_12_0_6;
  wire       [0:0]    state_out_12_0_7;
  wire       [0:0]    state_out_12_1_0;
  wire       [0:0]    state_out_12_1_1;
  wire       [0:0]    state_out_12_1_2;
  wire       [0:0]    state_out_12_1_3;
  wire       [0:0]    state_out_12_1_4;
  wire       [0:0]    state_out_12_1_5;
  wire       [0:0]    state_out_12_1_6;
  wire       [0:0]    state_out_12_1_7;
  wire       [0:0]    state_out_13_0_0;
  wire       [0:0]    state_out_13_0_1;
  wire       [0:0]    state_out_13_0_2;
  wire       [0:0]    state_out_13_0_3;
  wire       [0:0]    state_out_13_0_4;
  wire       [0:0]    state_out_13_0_5;
  wire       [0:0]    state_out_13_0_6;
  wire       [0:0]    state_out_13_0_7;
  wire       [0:0]    state_out_13_1_0;
  wire       [0:0]    state_out_13_1_1;
  wire       [0:0]    state_out_13_1_2;
  wire       [0:0]    state_out_13_1_3;
  wire       [0:0]    state_out_13_1_4;
  wire       [0:0]    state_out_13_1_5;
  wire       [0:0]    state_out_13_1_6;
  wire       [0:0]    state_out_13_1_7;
  wire       [0:0]    state_out_14_0_0;
  wire       [0:0]    state_out_14_0_1;
  wire       [0:0]    state_out_14_0_2;
  wire       [0:0]    state_out_14_0_3;
  wire       [0:0]    state_out_14_0_4;
  wire       [0:0]    state_out_14_0_5;
  wire       [0:0]    state_out_14_0_6;
  wire       [0:0]    state_out_14_0_7;
  wire       [0:0]    state_out_14_1_0;
  wire       [0:0]    state_out_14_1_1;
  wire       [0:0]    state_out_14_1_2;
  wire       [0:0]    state_out_14_1_3;
  wire       [0:0]    state_out_14_1_4;
  wire       [0:0]    state_out_14_1_5;
  wire       [0:0]    state_out_14_1_6;
  wire       [0:0]    state_out_14_1_7;
  wire       [0:0]    state_out_15_0_0;
  wire       [0:0]    state_out_15_0_1;
  wire       [0:0]    state_out_15_0_2;
  wire       [0:0]    state_out_15_0_3;
  wire       [0:0]    state_out_15_0_4;
  wire       [0:0]    state_out_15_0_5;
  wire       [0:0]    state_out_15_0_6;
  wire       [0:0]    state_out_15_0_7;
  wire       [0:0]    state_out_15_1_0;
  wire       [0:0]    state_out_15_1_1;
  wire       [0:0]    state_out_15_1_2;
  wire       [0:0]    state_out_15_1_3;
  wire       [0:0]    state_out_15_1_4;
  wire       [0:0]    state_out_15_1_5;
  wire       [0:0]    state_out_15_1_6;
  wire       [0:0]    state_out_15_1_7;

  Mul2 mul2_32 (
    .port_byte_in_0  (port_state_in_0_0_0    ), //i
    .port_byte_in_1  (port_state_in_0_0_1    ), //i
    .port_byte_in_2  (port_state_in_0_0_2    ), //i
    .port_byte_in_3  (port_state_in_0_0_3    ), //i
    .port_byte_in_4  (port_state_in_0_0_4    ), //i
    .port_byte_in_5  (port_state_in_0_0_5    ), //i
    .port_byte_in_6  (port_state_in_0_0_6    ), //i
    .port_byte_in_7  (port_state_in_0_0_7    ), //i
    .port_byte_out_0 (mul2_32_port_byte_out_0), //o
    .port_byte_out_1 (mul2_32_port_byte_out_1), //o
    .port_byte_out_2 (mul2_32_port_byte_out_2), //o
    .port_byte_out_3 (mul2_32_port_byte_out_3), //o
    .port_byte_out_4 (mul2_32_port_byte_out_4), //o
    .port_byte_out_5 (mul2_32_port_byte_out_5), //o
    .port_byte_out_6 (mul2_32_port_byte_out_6), //o
    .port_byte_out_7 (mul2_32_port_byte_out_7)  //o
  );
  Mul3 mul3_32 (
    .port_byte_in_0  (port_state_in_1_0_0    ), //i
    .port_byte_in_1  (port_state_in_1_0_1    ), //i
    .port_byte_in_2  (port_state_in_1_0_2    ), //i
    .port_byte_in_3  (port_state_in_1_0_3    ), //i
    .port_byte_in_4  (port_state_in_1_0_4    ), //i
    .port_byte_in_5  (port_state_in_1_0_5    ), //i
    .port_byte_in_6  (port_state_in_1_0_6    ), //i
    .port_byte_in_7  (port_state_in_1_0_7    ), //i
    .port_byte_out_0 (mul3_32_port_byte_out_0), //o
    .port_byte_out_1 (mul3_32_port_byte_out_1), //o
    .port_byte_out_2 (mul3_32_port_byte_out_2), //o
    .port_byte_out_3 (mul3_32_port_byte_out_3), //o
    .port_byte_out_4 (mul3_32_port_byte_out_4), //o
    .port_byte_out_5 (mul3_32_port_byte_out_5), //o
    .port_byte_out_6 (mul3_32_port_byte_out_6), //o
    .port_byte_out_7 (mul3_32_port_byte_out_7)  //o
  );
  Mul2 mul2_33 (
    .port_byte_in_0  (port_state_in_1_0_0    ), //i
    .port_byte_in_1  (port_state_in_1_0_1    ), //i
    .port_byte_in_2  (port_state_in_1_0_2    ), //i
    .port_byte_in_3  (port_state_in_1_0_3    ), //i
    .port_byte_in_4  (port_state_in_1_0_4    ), //i
    .port_byte_in_5  (port_state_in_1_0_5    ), //i
    .port_byte_in_6  (port_state_in_1_0_6    ), //i
    .port_byte_in_7  (port_state_in_1_0_7    ), //i
    .port_byte_out_0 (mul2_33_port_byte_out_0), //o
    .port_byte_out_1 (mul2_33_port_byte_out_1), //o
    .port_byte_out_2 (mul2_33_port_byte_out_2), //o
    .port_byte_out_3 (mul2_33_port_byte_out_3), //o
    .port_byte_out_4 (mul2_33_port_byte_out_4), //o
    .port_byte_out_5 (mul2_33_port_byte_out_5), //o
    .port_byte_out_6 (mul2_33_port_byte_out_6), //o
    .port_byte_out_7 (mul2_33_port_byte_out_7)  //o
  );
  Mul3 mul3_33 (
    .port_byte_in_0  (port_state_in_2_0_0    ), //i
    .port_byte_in_1  (port_state_in_2_0_1    ), //i
    .port_byte_in_2  (port_state_in_2_0_2    ), //i
    .port_byte_in_3  (port_state_in_2_0_3    ), //i
    .port_byte_in_4  (port_state_in_2_0_4    ), //i
    .port_byte_in_5  (port_state_in_2_0_5    ), //i
    .port_byte_in_6  (port_state_in_2_0_6    ), //i
    .port_byte_in_7  (port_state_in_2_0_7    ), //i
    .port_byte_out_0 (mul3_33_port_byte_out_0), //o
    .port_byte_out_1 (mul3_33_port_byte_out_1), //o
    .port_byte_out_2 (mul3_33_port_byte_out_2), //o
    .port_byte_out_3 (mul3_33_port_byte_out_3), //o
    .port_byte_out_4 (mul3_33_port_byte_out_4), //o
    .port_byte_out_5 (mul3_33_port_byte_out_5), //o
    .port_byte_out_6 (mul3_33_port_byte_out_6), //o
    .port_byte_out_7 (mul3_33_port_byte_out_7)  //o
  );
  Mul2 mul2_34 (
    .port_byte_in_0  (port_state_in_2_0_0    ), //i
    .port_byte_in_1  (port_state_in_2_0_1    ), //i
    .port_byte_in_2  (port_state_in_2_0_2    ), //i
    .port_byte_in_3  (port_state_in_2_0_3    ), //i
    .port_byte_in_4  (port_state_in_2_0_4    ), //i
    .port_byte_in_5  (port_state_in_2_0_5    ), //i
    .port_byte_in_6  (port_state_in_2_0_6    ), //i
    .port_byte_in_7  (port_state_in_2_0_7    ), //i
    .port_byte_out_0 (mul2_34_port_byte_out_0), //o
    .port_byte_out_1 (mul2_34_port_byte_out_1), //o
    .port_byte_out_2 (mul2_34_port_byte_out_2), //o
    .port_byte_out_3 (mul2_34_port_byte_out_3), //o
    .port_byte_out_4 (mul2_34_port_byte_out_4), //o
    .port_byte_out_5 (mul2_34_port_byte_out_5), //o
    .port_byte_out_6 (mul2_34_port_byte_out_6), //o
    .port_byte_out_7 (mul2_34_port_byte_out_7)  //o
  );
  Mul3 mul3_34 (
    .port_byte_in_0  (port_state_in_3_0_0    ), //i
    .port_byte_in_1  (port_state_in_3_0_1    ), //i
    .port_byte_in_2  (port_state_in_3_0_2    ), //i
    .port_byte_in_3  (port_state_in_3_0_3    ), //i
    .port_byte_in_4  (port_state_in_3_0_4    ), //i
    .port_byte_in_5  (port_state_in_3_0_5    ), //i
    .port_byte_in_6  (port_state_in_3_0_6    ), //i
    .port_byte_in_7  (port_state_in_3_0_7    ), //i
    .port_byte_out_0 (mul3_34_port_byte_out_0), //o
    .port_byte_out_1 (mul3_34_port_byte_out_1), //o
    .port_byte_out_2 (mul3_34_port_byte_out_2), //o
    .port_byte_out_3 (mul3_34_port_byte_out_3), //o
    .port_byte_out_4 (mul3_34_port_byte_out_4), //o
    .port_byte_out_5 (mul3_34_port_byte_out_5), //o
    .port_byte_out_6 (mul3_34_port_byte_out_6), //o
    .port_byte_out_7 (mul3_34_port_byte_out_7)  //o
  );
  Mul2 mul2_35 (
    .port_byte_in_0  (port_state_in_3_0_0    ), //i
    .port_byte_in_1  (port_state_in_3_0_1    ), //i
    .port_byte_in_2  (port_state_in_3_0_2    ), //i
    .port_byte_in_3  (port_state_in_3_0_3    ), //i
    .port_byte_in_4  (port_state_in_3_0_4    ), //i
    .port_byte_in_5  (port_state_in_3_0_5    ), //i
    .port_byte_in_6  (port_state_in_3_0_6    ), //i
    .port_byte_in_7  (port_state_in_3_0_7    ), //i
    .port_byte_out_0 (mul2_35_port_byte_out_0), //o
    .port_byte_out_1 (mul2_35_port_byte_out_1), //o
    .port_byte_out_2 (mul2_35_port_byte_out_2), //o
    .port_byte_out_3 (mul2_35_port_byte_out_3), //o
    .port_byte_out_4 (mul2_35_port_byte_out_4), //o
    .port_byte_out_5 (mul2_35_port_byte_out_5), //o
    .port_byte_out_6 (mul2_35_port_byte_out_6), //o
    .port_byte_out_7 (mul2_35_port_byte_out_7)  //o
  );
  Mul3 mul3_35 (
    .port_byte_in_0  (port_state_in_0_0_0    ), //i
    .port_byte_in_1  (port_state_in_0_0_1    ), //i
    .port_byte_in_2  (port_state_in_0_0_2    ), //i
    .port_byte_in_3  (port_state_in_0_0_3    ), //i
    .port_byte_in_4  (port_state_in_0_0_4    ), //i
    .port_byte_in_5  (port_state_in_0_0_5    ), //i
    .port_byte_in_6  (port_state_in_0_0_6    ), //i
    .port_byte_in_7  (port_state_in_0_0_7    ), //i
    .port_byte_out_0 (mul3_35_port_byte_out_0), //o
    .port_byte_out_1 (mul3_35_port_byte_out_1), //o
    .port_byte_out_2 (mul3_35_port_byte_out_2), //o
    .port_byte_out_3 (mul3_35_port_byte_out_3), //o
    .port_byte_out_4 (mul3_35_port_byte_out_4), //o
    .port_byte_out_5 (mul3_35_port_byte_out_5), //o
    .port_byte_out_6 (mul3_35_port_byte_out_6), //o
    .port_byte_out_7 (mul3_35_port_byte_out_7)  //o
  );
  Mul2 mul2_36 (
    .port_byte_in_0  (port_state_in_0_1_0    ), //i
    .port_byte_in_1  (port_state_in_0_1_1    ), //i
    .port_byte_in_2  (port_state_in_0_1_2    ), //i
    .port_byte_in_3  (port_state_in_0_1_3    ), //i
    .port_byte_in_4  (port_state_in_0_1_4    ), //i
    .port_byte_in_5  (port_state_in_0_1_5    ), //i
    .port_byte_in_6  (port_state_in_0_1_6    ), //i
    .port_byte_in_7  (port_state_in_0_1_7    ), //i
    .port_byte_out_0 (mul2_36_port_byte_out_0), //o
    .port_byte_out_1 (mul2_36_port_byte_out_1), //o
    .port_byte_out_2 (mul2_36_port_byte_out_2), //o
    .port_byte_out_3 (mul2_36_port_byte_out_3), //o
    .port_byte_out_4 (mul2_36_port_byte_out_4), //o
    .port_byte_out_5 (mul2_36_port_byte_out_5), //o
    .port_byte_out_6 (mul2_36_port_byte_out_6), //o
    .port_byte_out_7 (mul2_36_port_byte_out_7)  //o
  );
  Mul3 mul3_36 (
    .port_byte_in_0  (port_state_in_1_1_0    ), //i
    .port_byte_in_1  (port_state_in_1_1_1    ), //i
    .port_byte_in_2  (port_state_in_1_1_2    ), //i
    .port_byte_in_3  (port_state_in_1_1_3    ), //i
    .port_byte_in_4  (port_state_in_1_1_4    ), //i
    .port_byte_in_5  (port_state_in_1_1_5    ), //i
    .port_byte_in_6  (port_state_in_1_1_6    ), //i
    .port_byte_in_7  (port_state_in_1_1_7    ), //i
    .port_byte_out_0 (mul3_36_port_byte_out_0), //o
    .port_byte_out_1 (mul3_36_port_byte_out_1), //o
    .port_byte_out_2 (mul3_36_port_byte_out_2), //o
    .port_byte_out_3 (mul3_36_port_byte_out_3), //o
    .port_byte_out_4 (mul3_36_port_byte_out_4), //o
    .port_byte_out_5 (mul3_36_port_byte_out_5), //o
    .port_byte_out_6 (mul3_36_port_byte_out_6), //o
    .port_byte_out_7 (mul3_36_port_byte_out_7)  //o
  );
  Mul2 mul2_37 (
    .port_byte_in_0  (port_state_in_1_1_0    ), //i
    .port_byte_in_1  (port_state_in_1_1_1    ), //i
    .port_byte_in_2  (port_state_in_1_1_2    ), //i
    .port_byte_in_3  (port_state_in_1_1_3    ), //i
    .port_byte_in_4  (port_state_in_1_1_4    ), //i
    .port_byte_in_5  (port_state_in_1_1_5    ), //i
    .port_byte_in_6  (port_state_in_1_1_6    ), //i
    .port_byte_in_7  (port_state_in_1_1_7    ), //i
    .port_byte_out_0 (mul2_37_port_byte_out_0), //o
    .port_byte_out_1 (mul2_37_port_byte_out_1), //o
    .port_byte_out_2 (mul2_37_port_byte_out_2), //o
    .port_byte_out_3 (mul2_37_port_byte_out_3), //o
    .port_byte_out_4 (mul2_37_port_byte_out_4), //o
    .port_byte_out_5 (mul2_37_port_byte_out_5), //o
    .port_byte_out_6 (mul2_37_port_byte_out_6), //o
    .port_byte_out_7 (mul2_37_port_byte_out_7)  //o
  );
  Mul3 mul3_37 (
    .port_byte_in_0  (port_state_in_2_1_0    ), //i
    .port_byte_in_1  (port_state_in_2_1_1    ), //i
    .port_byte_in_2  (port_state_in_2_1_2    ), //i
    .port_byte_in_3  (port_state_in_2_1_3    ), //i
    .port_byte_in_4  (port_state_in_2_1_4    ), //i
    .port_byte_in_5  (port_state_in_2_1_5    ), //i
    .port_byte_in_6  (port_state_in_2_1_6    ), //i
    .port_byte_in_7  (port_state_in_2_1_7    ), //i
    .port_byte_out_0 (mul3_37_port_byte_out_0), //o
    .port_byte_out_1 (mul3_37_port_byte_out_1), //o
    .port_byte_out_2 (mul3_37_port_byte_out_2), //o
    .port_byte_out_3 (mul3_37_port_byte_out_3), //o
    .port_byte_out_4 (mul3_37_port_byte_out_4), //o
    .port_byte_out_5 (mul3_37_port_byte_out_5), //o
    .port_byte_out_6 (mul3_37_port_byte_out_6), //o
    .port_byte_out_7 (mul3_37_port_byte_out_7)  //o
  );
  Mul2 mul2_38 (
    .port_byte_in_0  (port_state_in_2_1_0    ), //i
    .port_byte_in_1  (port_state_in_2_1_1    ), //i
    .port_byte_in_2  (port_state_in_2_1_2    ), //i
    .port_byte_in_3  (port_state_in_2_1_3    ), //i
    .port_byte_in_4  (port_state_in_2_1_4    ), //i
    .port_byte_in_5  (port_state_in_2_1_5    ), //i
    .port_byte_in_6  (port_state_in_2_1_6    ), //i
    .port_byte_in_7  (port_state_in_2_1_7    ), //i
    .port_byte_out_0 (mul2_38_port_byte_out_0), //o
    .port_byte_out_1 (mul2_38_port_byte_out_1), //o
    .port_byte_out_2 (mul2_38_port_byte_out_2), //o
    .port_byte_out_3 (mul2_38_port_byte_out_3), //o
    .port_byte_out_4 (mul2_38_port_byte_out_4), //o
    .port_byte_out_5 (mul2_38_port_byte_out_5), //o
    .port_byte_out_6 (mul2_38_port_byte_out_6), //o
    .port_byte_out_7 (mul2_38_port_byte_out_7)  //o
  );
  Mul3 mul3_38 (
    .port_byte_in_0  (port_state_in_3_1_0    ), //i
    .port_byte_in_1  (port_state_in_3_1_1    ), //i
    .port_byte_in_2  (port_state_in_3_1_2    ), //i
    .port_byte_in_3  (port_state_in_3_1_3    ), //i
    .port_byte_in_4  (port_state_in_3_1_4    ), //i
    .port_byte_in_5  (port_state_in_3_1_5    ), //i
    .port_byte_in_6  (port_state_in_3_1_6    ), //i
    .port_byte_in_7  (port_state_in_3_1_7    ), //i
    .port_byte_out_0 (mul3_38_port_byte_out_0), //o
    .port_byte_out_1 (mul3_38_port_byte_out_1), //o
    .port_byte_out_2 (mul3_38_port_byte_out_2), //o
    .port_byte_out_3 (mul3_38_port_byte_out_3), //o
    .port_byte_out_4 (mul3_38_port_byte_out_4), //o
    .port_byte_out_5 (mul3_38_port_byte_out_5), //o
    .port_byte_out_6 (mul3_38_port_byte_out_6), //o
    .port_byte_out_7 (mul3_38_port_byte_out_7)  //o
  );
  Mul2 mul2_39 (
    .port_byte_in_0  (port_state_in_3_1_0    ), //i
    .port_byte_in_1  (port_state_in_3_1_1    ), //i
    .port_byte_in_2  (port_state_in_3_1_2    ), //i
    .port_byte_in_3  (port_state_in_3_1_3    ), //i
    .port_byte_in_4  (port_state_in_3_1_4    ), //i
    .port_byte_in_5  (port_state_in_3_1_5    ), //i
    .port_byte_in_6  (port_state_in_3_1_6    ), //i
    .port_byte_in_7  (port_state_in_3_1_7    ), //i
    .port_byte_out_0 (mul2_39_port_byte_out_0), //o
    .port_byte_out_1 (mul2_39_port_byte_out_1), //o
    .port_byte_out_2 (mul2_39_port_byte_out_2), //o
    .port_byte_out_3 (mul2_39_port_byte_out_3), //o
    .port_byte_out_4 (mul2_39_port_byte_out_4), //o
    .port_byte_out_5 (mul2_39_port_byte_out_5), //o
    .port_byte_out_6 (mul2_39_port_byte_out_6), //o
    .port_byte_out_7 (mul2_39_port_byte_out_7)  //o
  );
  Mul3 mul3_39 (
    .port_byte_in_0  (port_state_in_0_1_0    ), //i
    .port_byte_in_1  (port_state_in_0_1_1    ), //i
    .port_byte_in_2  (port_state_in_0_1_2    ), //i
    .port_byte_in_3  (port_state_in_0_1_3    ), //i
    .port_byte_in_4  (port_state_in_0_1_4    ), //i
    .port_byte_in_5  (port_state_in_0_1_5    ), //i
    .port_byte_in_6  (port_state_in_0_1_6    ), //i
    .port_byte_in_7  (port_state_in_0_1_7    ), //i
    .port_byte_out_0 (mul3_39_port_byte_out_0), //o
    .port_byte_out_1 (mul3_39_port_byte_out_1), //o
    .port_byte_out_2 (mul3_39_port_byte_out_2), //o
    .port_byte_out_3 (mul3_39_port_byte_out_3), //o
    .port_byte_out_4 (mul3_39_port_byte_out_4), //o
    .port_byte_out_5 (mul3_39_port_byte_out_5), //o
    .port_byte_out_6 (mul3_39_port_byte_out_6), //o
    .port_byte_out_7 (mul3_39_port_byte_out_7)  //o
  );
  Mul2 mul2_40 (
    .port_byte_in_0  (port_state_in_4_0_0    ), //i
    .port_byte_in_1  (port_state_in_4_0_1    ), //i
    .port_byte_in_2  (port_state_in_4_0_2    ), //i
    .port_byte_in_3  (port_state_in_4_0_3    ), //i
    .port_byte_in_4  (port_state_in_4_0_4    ), //i
    .port_byte_in_5  (port_state_in_4_0_5    ), //i
    .port_byte_in_6  (port_state_in_4_0_6    ), //i
    .port_byte_in_7  (port_state_in_4_0_7    ), //i
    .port_byte_out_0 (mul2_40_port_byte_out_0), //o
    .port_byte_out_1 (mul2_40_port_byte_out_1), //o
    .port_byte_out_2 (mul2_40_port_byte_out_2), //o
    .port_byte_out_3 (mul2_40_port_byte_out_3), //o
    .port_byte_out_4 (mul2_40_port_byte_out_4), //o
    .port_byte_out_5 (mul2_40_port_byte_out_5), //o
    .port_byte_out_6 (mul2_40_port_byte_out_6), //o
    .port_byte_out_7 (mul2_40_port_byte_out_7)  //o
  );
  Mul3 mul3_40 (
    .port_byte_in_0  (port_state_in_5_0_0    ), //i
    .port_byte_in_1  (port_state_in_5_0_1    ), //i
    .port_byte_in_2  (port_state_in_5_0_2    ), //i
    .port_byte_in_3  (port_state_in_5_0_3    ), //i
    .port_byte_in_4  (port_state_in_5_0_4    ), //i
    .port_byte_in_5  (port_state_in_5_0_5    ), //i
    .port_byte_in_6  (port_state_in_5_0_6    ), //i
    .port_byte_in_7  (port_state_in_5_0_7    ), //i
    .port_byte_out_0 (mul3_40_port_byte_out_0), //o
    .port_byte_out_1 (mul3_40_port_byte_out_1), //o
    .port_byte_out_2 (mul3_40_port_byte_out_2), //o
    .port_byte_out_3 (mul3_40_port_byte_out_3), //o
    .port_byte_out_4 (mul3_40_port_byte_out_4), //o
    .port_byte_out_5 (mul3_40_port_byte_out_5), //o
    .port_byte_out_6 (mul3_40_port_byte_out_6), //o
    .port_byte_out_7 (mul3_40_port_byte_out_7)  //o
  );
  Mul2 mul2_41 (
    .port_byte_in_0  (port_state_in_5_0_0    ), //i
    .port_byte_in_1  (port_state_in_5_0_1    ), //i
    .port_byte_in_2  (port_state_in_5_0_2    ), //i
    .port_byte_in_3  (port_state_in_5_0_3    ), //i
    .port_byte_in_4  (port_state_in_5_0_4    ), //i
    .port_byte_in_5  (port_state_in_5_0_5    ), //i
    .port_byte_in_6  (port_state_in_5_0_6    ), //i
    .port_byte_in_7  (port_state_in_5_0_7    ), //i
    .port_byte_out_0 (mul2_41_port_byte_out_0), //o
    .port_byte_out_1 (mul2_41_port_byte_out_1), //o
    .port_byte_out_2 (mul2_41_port_byte_out_2), //o
    .port_byte_out_3 (mul2_41_port_byte_out_3), //o
    .port_byte_out_4 (mul2_41_port_byte_out_4), //o
    .port_byte_out_5 (mul2_41_port_byte_out_5), //o
    .port_byte_out_6 (mul2_41_port_byte_out_6), //o
    .port_byte_out_7 (mul2_41_port_byte_out_7)  //o
  );
  Mul3 mul3_41 (
    .port_byte_in_0  (port_state_in_6_0_0    ), //i
    .port_byte_in_1  (port_state_in_6_0_1    ), //i
    .port_byte_in_2  (port_state_in_6_0_2    ), //i
    .port_byte_in_3  (port_state_in_6_0_3    ), //i
    .port_byte_in_4  (port_state_in_6_0_4    ), //i
    .port_byte_in_5  (port_state_in_6_0_5    ), //i
    .port_byte_in_6  (port_state_in_6_0_6    ), //i
    .port_byte_in_7  (port_state_in_6_0_7    ), //i
    .port_byte_out_0 (mul3_41_port_byte_out_0), //o
    .port_byte_out_1 (mul3_41_port_byte_out_1), //o
    .port_byte_out_2 (mul3_41_port_byte_out_2), //o
    .port_byte_out_3 (mul3_41_port_byte_out_3), //o
    .port_byte_out_4 (mul3_41_port_byte_out_4), //o
    .port_byte_out_5 (mul3_41_port_byte_out_5), //o
    .port_byte_out_6 (mul3_41_port_byte_out_6), //o
    .port_byte_out_7 (mul3_41_port_byte_out_7)  //o
  );
  Mul2 mul2_42 (
    .port_byte_in_0  (port_state_in_6_0_0    ), //i
    .port_byte_in_1  (port_state_in_6_0_1    ), //i
    .port_byte_in_2  (port_state_in_6_0_2    ), //i
    .port_byte_in_3  (port_state_in_6_0_3    ), //i
    .port_byte_in_4  (port_state_in_6_0_4    ), //i
    .port_byte_in_5  (port_state_in_6_0_5    ), //i
    .port_byte_in_6  (port_state_in_6_0_6    ), //i
    .port_byte_in_7  (port_state_in_6_0_7    ), //i
    .port_byte_out_0 (mul2_42_port_byte_out_0), //o
    .port_byte_out_1 (mul2_42_port_byte_out_1), //o
    .port_byte_out_2 (mul2_42_port_byte_out_2), //o
    .port_byte_out_3 (mul2_42_port_byte_out_3), //o
    .port_byte_out_4 (mul2_42_port_byte_out_4), //o
    .port_byte_out_5 (mul2_42_port_byte_out_5), //o
    .port_byte_out_6 (mul2_42_port_byte_out_6), //o
    .port_byte_out_7 (mul2_42_port_byte_out_7)  //o
  );
  Mul3 mul3_42 (
    .port_byte_in_0  (port_state_in_7_0_0    ), //i
    .port_byte_in_1  (port_state_in_7_0_1    ), //i
    .port_byte_in_2  (port_state_in_7_0_2    ), //i
    .port_byte_in_3  (port_state_in_7_0_3    ), //i
    .port_byte_in_4  (port_state_in_7_0_4    ), //i
    .port_byte_in_5  (port_state_in_7_0_5    ), //i
    .port_byte_in_6  (port_state_in_7_0_6    ), //i
    .port_byte_in_7  (port_state_in_7_0_7    ), //i
    .port_byte_out_0 (mul3_42_port_byte_out_0), //o
    .port_byte_out_1 (mul3_42_port_byte_out_1), //o
    .port_byte_out_2 (mul3_42_port_byte_out_2), //o
    .port_byte_out_3 (mul3_42_port_byte_out_3), //o
    .port_byte_out_4 (mul3_42_port_byte_out_4), //o
    .port_byte_out_5 (mul3_42_port_byte_out_5), //o
    .port_byte_out_6 (mul3_42_port_byte_out_6), //o
    .port_byte_out_7 (mul3_42_port_byte_out_7)  //o
  );
  Mul2 mul2_43 (
    .port_byte_in_0  (port_state_in_7_0_0    ), //i
    .port_byte_in_1  (port_state_in_7_0_1    ), //i
    .port_byte_in_2  (port_state_in_7_0_2    ), //i
    .port_byte_in_3  (port_state_in_7_0_3    ), //i
    .port_byte_in_4  (port_state_in_7_0_4    ), //i
    .port_byte_in_5  (port_state_in_7_0_5    ), //i
    .port_byte_in_6  (port_state_in_7_0_6    ), //i
    .port_byte_in_7  (port_state_in_7_0_7    ), //i
    .port_byte_out_0 (mul2_43_port_byte_out_0), //o
    .port_byte_out_1 (mul2_43_port_byte_out_1), //o
    .port_byte_out_2 (mul2_43_port_byte_out_2), //o
    .port_byte_out_3 (mul2_43_port_byte_out_3), //o
    .port_byte_out_4 (mul2_43_port_byte_out_4), //o
    .port_byte_out_5 (mul2_43_port_byte_out_5), //o
    .port_byte_out_6 (mul2_43_port_byte_out_6), //o
    .port_byte_out_7 (mul2_43_port_byte_out_7)  //o
  );
  Mul3 mul3_43 (
    .port_byte_in_0  (port_state_in_4_0_0    ), //i
    .port_byte_in_1  (port_state_in_4_0_1    ), //i
    .port_byte_in_2  (port_state_in_4_0_2    ), //i
    .port_byte_in_3  (port_state_in_4_0_3    ), //i
    .port_byte_in_4  (port_state_in_4_0_4    ), //i
    .port_byte_in_5  (port_state_in_4_0_5    ), //i
    .port_byte_in_6  (port_state_in_4_0_6    ), //i
    .port_byte_in_7  (port_state_in_4_0_7    ), //i
    .port_byte_out_0 (mul3_43_port_byte_out_0), //o
    .port_byte_out_1 (mul3_43_port_byte_out_1), //o
    .port_byte_out_2 (mul3_43_port_byte_out_2), //o
    .port_byte_out_3 (mul3_43_port_byte_out_3), //o
    .port_byte_out_4 (mul3_43_port_byte_out_4), //o
    .port_byte_out_5 (mul3_43_port_byte_out_5), //o
    .port_byte_out_6 (mul3_43_port_byte_out_6), //o
    .port_byte_out_7 (mul3_43_port_byte_out_7)  //o
  );
  Mul2 mul2_44 (
    .port_byte_in_0  (port_state_in_4_1_0    ), //i
    .port_byte_in_1  (port_state_in_4_1_1    ), //i
    .port_byte_in_2  (port_state_in_4_1_2    ), //i
    .port_byte_in_3  (port_state_in_4_1_3    ), //i
    .port_byte_in_4  (port_state_in_4_1_4    ), //i
    .port_byte_in_5  (port_state_in_4_1_5    ), //i
    .port_byte_in_6  (port_state_in_4_1_6    ), //i
    .port_byte_in_7  (port_state_in_4_1_7    ), //i
    .port_byte_out_0 (mul2_44_port_byte_out_0), //o
    .port_byte_out_1 (mul2_44_port_byte_out_1), //o
    .port_byte_out_2 (mul2_44_port_byte_out_2), //o
    .port_byte_out_3 (mul2_44_port_byte_out_3), //o
    .port_byte_out_4 (mul2_44_port_byte_out_4), //o
    .port_byte_out_5 (mul2_44_port_byte_out_5), //o
    .port_byte_out_6 (mul2_44_port_byte_out_6), //o
    .port_byte_out_7 (mul2_44_port_byte_out_7)  //o
  );
  Mul3 mul3_44 (
    .port_byte_in_0  (port_state_in_5_1_0    ), //i
    .port_byte_in_1  (port_state_in_5_1_1    ), //i
    .port_byte_in_2  (port_state_in_5_1_2    ), //i
    .port_byte_in_3  (port_state_in_5_1_3    ), //i
    .port_byte_in_4  (port_state_in_5_1_4    ), //i
    .port_byte_in_5  (port_state_in_5_1_5    ), //i
    .port_byte_in_6  (port_state_in_5_1_6    ), //i
    .port_byte_in_7  (port_state_in_5_1_7    ), //i
    .port_byte_out_0 (mul3_44_port_byte_out_0), //o
    .port_byte_out_1 (mul3_44_port_byte_out_1), //o
    .port_byte_out_2 (mul3_44_port_byte_out_2), //o
    .port_byte_out_3 (mul3_44_port_byte_out_3), //o
    .port_byte_out_4 (mul3_44_port_byte_out_4), //o
    .port_byte_out_5 (mul3_44_port_byte_out_5), //o
    .port_byte_out_6 (mul3_44_port_byte_out_6), //o
    .port_byte_out_7 (mul3_44_port_byte_out_7)  //o
  );
  Mul2 mul2_45 (
    .port_byte_in_0  (port_state_in_5_1_0    ), //i
    .port_byte_in_1  (port_state_in_5_1_1    ), //i
    .port_byte_in_2  (port_state_in_5_1_2    ), //i
    .port_byte_in_3  (port_state_in_5_1_3    ), //i
    .port_byte_in_4  (port_state_in_5_1_4    ), //i
    .port_byte_in_5  (port_state_in_5_1_5    ), //i
    .port_byte_in_6  (port_state_in_5_1_6    ), //i
    .port_byte_in_7  (port_state_in_5_1_7    ), //i
    .port_byte_out_0 (mul2_45_port_byte_out_0), //o
    .port_byte_out_1 (mul2_45_port_byte_out_1), //o
    .port_byte_out_2 (mul2_45_port_byte_out_2), //o
    .port_byte_out_3 (mul2_45_port_byte_out_3), //o
    .port_byte_out_4 (mul2_45_port_byte_out_4), //o
    .port_byte_out_5 (mul2_45_port_byte_out_5), //o
    .port_byte_out_6 (mul2_45_port_byte_out_6), //o
    .port_byte_out_7 (mul2_45_port_byte_out_7)  //o
  );
  Mul3 mul3_45 (
    .port_byte_in_0  (port_state_in_6_1_0    ), //i
    .port_byte_in_1  (port_state_in_6_1_1    ), //i
    .port_byte_in_2  (port_state_in_6_1_2    ), //i
    .port_byte_in_3  (port_state_in_6_1_3    ), //i
    .port_byte_in_4  (port_state_in_6_1_4    ), //i
    .port_byte_in_5  (port_state_in_6_1_5    ), //i
    .port_byte_in_6  (port_state_in_6_1_6    ), //i
    .port_byte_in_7  (port_state_in_6_1_7    ), //i
    .port_byte_out_0 (mul3_45_port_byte_out_0), //o
    .port_byte_out_1 (mul3_45_port_byte_out_1), //o
    .port_byte_out_2 (mul3_45_port_byte_out_2), //o
    .port_byte_out_3 (mul3_45_port_byte_out_3), //o
    .port_byte_out_4 (mul3_45_port_byte_out_4), //o
    .port_byte_out_5 (mul3_45_port_byte_out_5), //o
    .port_byte_out_6 (mul3_45_port_byte_out_6), //o
    .port_byte_out_7 (mul3_45_port_byte_out_7)  //o
  );
  Mul2 mul2_46 (
    .port_byte_in_0  (port_state_in_6_1_0    ), //i
    .port_byte_in_1  (port_state_in_6_1_1    ), //i
    .port_byte_in_2  (port_state_in_6_1_2    ), //i
    .port_byte_in_3  (port_state_in_6_1_3    ), //i
    .port_byte_in_4  (port_state_in_6_1_4    ), //i
    .port_byte_in_5  (port_state_in_6_1_5    ), //i
    .port_byte_in_6  (port_state_in_6_1_6    ), //i
    .port_byte_in_7  (port_state_in_6_1_7    ), //i
    .port_byte_out_0 (mul2_46_port_byte_out_0), //o
    .port_byte_out_1 (mul2_46_port_byte_out_1), //o
    .port_byte_out_2 (mul2_46_port_byte_out_2), //o
    .port_byte_out_3 (mul2_46_port_byte_out_3), //o
    .port_byte_out_4 (mul2_46_port_byte_out_4), //o
    .port_byte_out_5 (mul2_46_port_byte_out_5), //o
    .port_byte_out_6 (mul2_46_port_byte_out_6), //o
    .port_byte_out_7 (mul2_46_port_byte_out_7)  //o
  );
  Mul3 mul3_46 (
    .port_byte_in_0  (port_state_in_7_1_0    ), //i
    .port_byte_in_1  (port_state_in_7_1_1    ), //i
    .port_byte_in_2  (port_state_in_7_1_2    ), //i
    .port_byte_in_3  (port_state_in_7_1_3    ), //i
    .port_byte_in_4  (port_state_in_7_1_4    ), //i
    .port_byte_in_5  (port_state_in_7_1_5    ), //i
    .port_byte_in_6  (port_state_in_7_1_6    ), //i
    .port_byte_in_7  (port_state_in_7_1_7    ), //i
    .port_byte_out_0 (mul3_46_port_byte_out_0), //o
    .port_byte_out_1 (mul3_46_port_byte_out_1), //o
    .port_byte_out_2 (mul3_46_port_byte_out_2), //o
    .port_byte_out_3 (mul3_46_port_byte_out_3), //o
    .port_byte_out_4 (mul3_46_port_byte_out_4), //o
    .port_byte_out_5 (mul3_46_port_byte_out_5), //o
    .port_byte_out_6 (mul3_46_port_byte_out_6), //o
    .port_byte_out_7 (mul3_46_port_byte_out_7)  //o
  );
  Mul2 mul2_47 (
    .port_byte_in_0  (port_state_in_7_1_0    ), //i
    .port_byte_in_1  (port_state_in_7_1_1    ), //i
    .port_byte_in_2  (port_state_in_7_1_2    ), //i
    .port_byte_in_3  (port_state_in_7_1_3    ), //i
    .port_byte_in_4  (port_state_in_7_1_4    ), //i
    .port_byte_in_5  (port_state_in_7_1_5    ), //i
    .port_byte_in_6  (port_state_in_7_1_6    ), //i
    .port_byte_in_7  (port_state_in_7_1_7    ), //i
    .port_byte_out_0 (mul2_47_port_byte_out_0), //o
    .port_byte_out_1 (mul2_47_port_byte_out_1), //o
    .port_byte_out_2 (mul2_47_port_byte_out_2), //o
    .port_byte_out_3 (mul2_47_port_byte_out_3), //o
    .port_byte_out_4 (mul2_47_port_byte_out_4), //o
    .port_byte_out_5 (mul2_47_port_byte_out_5), //o
    .port_byte_out_6 (mul2_47_port_byte_out_6), //o
    .port_byte_out_7 (mul2_47_port_byte_out_7)  //o
  );
  Mul3 mul3_47 (
    .port_byte_in_0  (port_state_in_4_1_0    ), //i
    .port_byte_in_1  (port_state_in_4_1_1    ), //i
    .port_byte_in_2  (port_state_in_4_1_2    ), //i
    .port_byte_in_3  (port_state_in_4_1_3    ), //i
    .port_byte_in_4  (port_state_in_4_1_4    ), //i
    .port_byte_in_5  (port_state_in_4_1_5    ), //i
    .port_byte_in_6  (port_state_in_4_1_6    ), //i
    .port_byte_in_7  (port_state_in_4_1_7    ), //i
    .port_byte_out_0 (mul3_47_port_byte_out_0), //o
    .port_byte_out_1 (mul3_47_port_byte_out_1), //o
    .port_byte_out_2 (mul3_47_port_byte_out_2), //o
    .port_byte_out_3 (mul3_47_port_byte_out_3), //o
    .port_byte_out_4 (mul3_47_port_byte_out_4), //o
    .port_byte_out_5 (mul3_47_port_byte_out_5), //o
    .port_byte_out_6 (mul3_47_port_byte_out_6), //o
    .port_byte_out_7 (mul3_47_port_byte_out_7)  //o
  );
  Mul2 mul2_48 (
    .port_byte_in_0  (port_state_in_8_0_0    ), //i
    .port_byte_in_1  (port_state_in_8_0_1    ), //i
    .port_byte_in_2  (port_state_in_8_0_2    ), //i
    .port_byte_in_3  (port_state_in_8_0_3    ), //i
    .port_byte_in_4  (port_state_in_8_0_4    ), //i
    .port_byte_in_5  (port_state_in_8_0_5    ), //i
    .port_byte_in_6  (port_state_in_8_0_6    ), //i
    .port_byte_in_7  (port_state_in_8_0_7    ), //i
    .port_byte_out_0 (mul2_48_port_byte_out_0), //o
    .port_byte_out_1 (mul2_48_port_byte_out_1), //o
    .port_byte_out_2 (mul2_48_port_byte_out_2), //o
    .port_byte_out_3 (mul2_48_port_byte_out_3), //o
    .port_byte_out_4 (mul2_48_port_byte_out_4), //o
    .port_byte_out_5 (mul2_48_port_byte_out_5), //o
    .port_byte_out_6 (mul2_48_port_byte_out_6), //o
    .port_byte_out_7 (mul2_48_port_byte_out_7)  //o
  );
  Mul3 mul3_48 (
    .port_byte_in_0  (port_state_in_9_0_0    ), //i
    .port_byte_in_1  (port_state_in_9_0_1    ), //i
    .port_byte_in_2  (port_state_in_9_0_2    ), //i
    .port_byte_in_3  (port_state_in_9_0_3    ), //i
    .port_byte_in_4  (port_state_in_9_0_4    ), //i
    .port_byte_in_5  (port_state_in_9_0_5    ), //i
    .port_byte_in_6  (port_state_in_9_0_6    ), //i
    .port_byte_in_7  (port_state_in_9_0_7    ), //i
    .port_byte_out_0 (mul3_48_port_byte_out_0), //o
    .port_byte_out_1 (mul3_48_port_byte_out_1), //o
    .port_byte_out_2 (mul3_48_port_byte_out_2), //o
    .port_byte_out_3 (mul3_48_port_byte_out_3), //o
    .port_byte_out_4 (mul3_48_port_byte_out_4), //o
    .port_byte_out_5 (mul3_48_port_byte_out_5), //o
    .port_byte_out_6 (mul3_48_port_byte_out_6), //o
    .port_byte_out_7 (mul3_48_port_byte_out_7)  //o
  );
  Mul2 mul2_49 (
    .port_byte_in_0  (port_state_in_9_0_0    ), //i
    .port_byte_in_1  (port_state_in_9_0_1    ), //i
    .port_byte_in_2  (port_state_in_9_0_2    ), //i
    .port_byte_in_3  (port_state_in_9_0_3    ), //i
    .port_byte_in_4  (port_state_in_9_0_4    ), //i
    .port_byte_in_5  (port_state_in_9_0_5    ), //i
    .port_byte_in_6  (port_state_in_9_0_6    ), //i
    .port_byte_in_7  (port_state_in_9_0_7    ), //i
    .port_byte_out_0 (mul2_49_port_byte_out_0), //o
    .port_byte_out_1 (mul2_49_port_byte_out_1), //o
    .port_byte_out_2 (mul2_49_port_byte_out_2), //o
    .port_byte_out_3 (mul2_49_port_byte_out_3), //o
    .port_byte_out_4 (mul2_49_port_byte_out_4), //o
    .port_byte_out_5 (mul2_49_port_byte_out_5), //o
    .port_byte_out_6 (mul2_49_port_byte_out_6), //o
    .port_byte_out_7 (mul2_49_port_byte_out_7)  //o
  );
  Mul3 mul3_49 (
    .port_byte_in_0  (port_state_in_10_0_0   ), //i
    .port_byte_in_1  (port_state_in_10_0_1   ), //i
    .port_byte_in_2  (port_state_in_10_0_2   ), //i
    .port_byte_in_3  (port_state_in_10_0_3   ), //i
    .port_byte_in_4  (port_state_in_10_0_4   ), //i
    .port_byte_in_5  (port_state_in_10_0_5   ), //i
    .port_byte_in_6  (port_state_in_10_0_6   ), //i
    .port_byte_in_7  (port_state_in_10_0_7   ), //i
    .port_byte_out_0 (mul3_49_port_byte_out_0), //o
    .port_byte_out_1 (mul3_49_port_byte_out_1), //o
    .port_byte_out_2 (mul3_49_port_byte_out_2), //o
    .port_byte_out_3 (mul3_49_port_byte_out_3), //o
    .port_byte_out_4 (mul3_49_port_byte_out_4), //o
    .port_byte_out_5 (mul3_49_port_byte_out_5), //o
    .port_byte_out_6 (mul3_49_port_byte_out_6), //o
    .port_byte_out_7 (mul3_49_port_byte_out_7)  //o
  );
  Mul2 mul2_50 (
    .port_byte_in_0  (port_state_in_10_0_0   ), //i
    .port_byte_in_1  (port_state_in_10_0_1   ), //i
    .port_byte_in_2  (port_state_in_10_0_2   ), //i
    .port_byte_in_3  (port_state_in_10_0_3   ), //i
    .port_byte_in_4  (port_state_in_10_0_4   ), //i
    .port_byte_in_5  (port_state_in_10_0_5   ), //i
    .port_byte_in_6  (port_state_in_10_0_6   ), //i
    .port_byte_in_7  (port_state_in_10_0_7   ), //i
    .port_byte_out_0 (mul2_50_port_byte_out_0), //o
    .port_byte_out_1 (mul2_50_port_byte_out_1), //o
    .port_byte_out_2 (mul2_50_port_byte_out_2), //o
    .port_byte_out_3 (mul2_50_port_byte_out_3), //o
    .port_byte_out_4 (mul2_50_port_byte_out_4), //o
    .port_byte_out_5 (mul2_50_port_byte_out_5), //o
    .port_byte_out_6 (mul2_50_port_byte_out_6), //o
    .port_byte_out_7 (mul2_50_port_byte_out_7)  //o
  );
  Mul3 mul3_50 (
    .port_byte_in_0  (port_state_in_11_0_0   ), //i
    .port_byte_in_1  (port_state_in_11_0_1   ), //i
    .port_byte_in_2  (port_state_in_11_0_2   ), //i
    .port_byte_in_3  (port_state_in_11_0_3   ), //i
    .port_byte_in_4  (port_state_in_11_0_4   ), //i
    .port_byte_in_5  (port_state_in_11_0_5   ), //i
    .port_byte_in_6  (port_state_in_11_0_6   ), //i
    .port_byte_in_7  (port_state_in_11_0_7   ), //i
    .port_byte_out_0 (mul3_50_port_byte_out_0), //o
    .port_byte_out_1 (mul3_50_port_byte_out_1), //o
    .port_byte_out_2 (mul3_50_port_byte_out_2), //o
    .port_byte_out_3 (mul3_50_port_byte_out_3), //o
    .port_byte_out_4 (mul3_50_port_byte_out_4), //o
    .port_byte_out_5 (mul3_50_port_byte_out_5), //o
    .port_byte_out_6 (mul3_50_port_byte_out_6), //o
    .port_byte_out_7 (mul3_50_port_byte_out_7)  //o
  );
  Mul2 mul2_51 (
    .port_byte_in_0  (port_state_in_11_0_0   ), //i
    .port_byte_in_1  (port_state_in_11_0_1   ), //i
    .port_byte_in_2  (port_state_in_11_0_2   ), //i
    .port_byte_in_3  (port_state_in_11_0_3   ), //i
    .port_byte_in_4  (port_state_in_11_0_4   ), //i
    .port_byte_in_5  (port_state_in_11_0_5   ), //i
    .port_byte_in_6  (port_state_in_11_0_6   ), //i
    .port_byte_in_7  (port_state_in_11_0_7   ), //i
    .port_byte_out_0 (mul2_51_port_byte_out_0), //o
    .port_byte_out_1 (mul2_51_port_byte_out_1), //o
    .port_byte_out_2 (mul2_51_port_byte_out_2), //o
    .port_byte_out_3 (mul2_51_port_byte_out_3), //o
    .port_byte_out_4 (mul2_51_port_byte_out_4), //o
    .port_byte_out_5 (mul2_51_port_byte_out_5), //o
    .port_byte_out_6 (mul2_51_port_byte_out_6), //o
    .port_byte_out_7 (mul2_51_port_byte_out_7)  //o
  );
  Mul3 mul3_51 (
    .port_byte_in_0  (port_state_in_8_0_0    ), //i
    .port_byte_in_1  (port_state_in_8_0_1    ), //i
    .port_byte_in_2  (port_state_in_8_0_2    ), //i
    .port_byte_in_3  (port_state_in_8_0_3    ), //i
    .port_byte_in_4  (port_state_in_8_0_4    ), //i
    .port_byte_in_5  (port_state_in_8_0_5    ), //i
    .port_byte_in_6  (port_state_in_8_0_6    ), //i
    .port_byte_in_7  (port_state_in_8_0_7    ), //i
    .port_byte_out_0 (mul3_51_port_byte_out_0), //o
    .port_byte_out_1 (mul3_51_port_byte_out_1), //o
    .port_byte_out_2 (mul3_51_port_byte_out_2), //o
    .port_byte_out_3 (mul3_51_port_byte_out_3), //o
    .port_byte_out_4 (mul3_51_port_byte_out_4), //o
    .port_byte_out_5 (mul3_51_port_byte_out_5), //o
    .port_byte_out_6 (mul3_51_port_byte_out_6), //o
    .port_byte_out_7 (mul3_51_port_byte_out_7)  //o
  );
  Mul2 mul2_52 (
    .port_byte_in_0  (port_state_in_8_1_0    ), //i
    .port_byte_in_1  (port_state_in_8_1_1    ), //i
    .port_byte_in_2  (port_state_in_8_1_2    ), //i
    .port_byte_in_3  (port_state_in_8_1_3    ), //i
    .port_byte_in_4  (port_state_in_8_1_4    ), //i
    .port_byte_in_5  (port_state_in_8_1_5    ), //i
    .port_byte_in_6  (port_state_in_8_1_6    ), //i
    .port_byte_in_7  (port_state_in_8_1_7    ), //i
    .port_byte_out_0 (mul2_52_port_byte_out_0), //o
    .port_byte_out_1 (mul2_52_port_byte_out_1), //o
    .port_byte_out_2 (mul2_52_port_byte_out_2), //o
    .port_byte_out_3 (mul2_52_port_byte_out_3), //o
    .port_byte_out_4 (mul2_52_port_byte_out_4), //o
    .port_byte_out_5 (mul2_52_port_byte_out_5), //o
    .port_byte_out_6 (mul2_52_port_byte_out_6), //o
    .port_byte_out_7 (mul2_52_port_byte_out_7)  //o
  );
  Mul3 mul3_52 (
    .port_byte_in_0  (port_state_in_9_1_0    ), //i
    .port_byte_in_1  (port_state_in_9_1_1    ), //i
    .port_byte_in_2  (port_state_in_9_1_2    ), //i
    .port_byte_in_3  (port_state_in_9_1_3    ), //i
    .port_byte_in_4  (port_state_in_9_1_4    ), //i
    .port_byte_in_5  (port_state_in_9_1_5    ), //i
    .port_byte_in_6  (port_state_in_9_1_6    ), //i
    .port_byte_in_7  (port_state_in_9_1_7    ), //i
    .port_byte_out_0 (mul3_52_port_byte_out_0), //o
    .port_byte_out_1 (mul3_52_port_byte_out_1), //o
    .port_byte_out_2 (mul3_52_port_byte_out_2), //o
    .port_byte_out_3 (mul3_52_port_byte_out_3), //o
    .port_byte_out_4 (mul3_52_port_byte_out_4), //o
    .port_byte_out_5 (mul3_52_port_byte_out_5), //o
    .port_byte_out_6 (mul3_52_port_byte_out_6), //o
    .port_byte_out_7 (mul3_52_port_byte_out_7)  //o
  );
  Mul2 mul2_53 (
    .port_byte_in_0  (port_state_in_9_1_0    ), //i
    .port_byte_in_1  (port_state_in_9_1_1    ), //i
    .port_byte_in_2  (port_state_in_9_1_2    ), //i
    .port_byte_in_3  (port_state_in_9_1_3    ), //i
    .port_byte_in_4  (port_state_in_9_1_4    ), //i
    .port_byte_in_5  (port_state_in_9_1_5    ), //i
    .port_byte_in_6  (port_state_in_9_1_6    ), //i
    .port_byte_in_7  (port_state_in_9_1_7    ), //i
    .port_byte_out_0 (mul2_53_port_byte_out_0), //o
    .port_byte_out_1 (mul2_53_port_byte_out_1), //o
    .port_byte_out_2 (mul2_53_port_byte_out_2), //o
    .port_byte_out_3 (mul2_53_port_byte_out_3), //o
    .port_byte_out_4 (mul2_53_port_byte_out_4), //o
    .port_byte_out_5 (mul2_53_port_byte_out_5), //o
    .port_byte_out_6 (mul2_53_port_byte_out_6), //o
    .port_byte_out_7 (mul2_53_port_byte_out_7)  //o
  );
  Mul3 mul3_53 (
    .port_byte_in_0  (port_state_in_10_1_0   ), //i
    .port_byte_in_1  (port_state_in_10_1_1   ), //i
    .port_byte_in_2  (port_state_in_10_1_2   ), //i
    .port_byte_in_3  (port_state_in_10_1_3   ), //i
    .port_byte_in_4  (port_state_in_10_1_4   ), //i
    .port_byte_in_5  (port_state_in_10_1_5   ), //i
    .port_byte_in_6  (port_state_in_10_1_6   ), //i
    .port_byte_in_7  (port_state_in_10_1_7   ), //i
    .port_byte_out_0 (mul3_53_port_byte_out_0), //o
    .port_byte_out_1 (mul3_53_port_byte_out_1), //o
    .port_byte_out_2 (mul3_53_port_byte_out_2), //o
    .port_byte_out_3 (mul3_53_port_byte_out_3), //o
    .port_byte_out_4 (mul3_53_port_byte_out_4), //o
    .port_byte_out_5 (mul3_53_port_byte_out_5), //o
    .port_byte_out_6 (mul3_53_port_byte_out_6), //o
    .port_byte_out_7 (mul3_53_port_byte_out_7)  //o
  );
  Mul2 mul2_54 (
    .port_byte_in_0  (port_state_in_10_1_0   ), //i
    .port_byte_in_1  (port_state_in_10_1_1   ), //i
    .port_byte_in_2  (port_state_in_10_1_2   ), //i
    .port_byte_in_3  (port_state_in_10_1_3   ), //i
    .port_byte_in_4  (port_state_in_10_1_4   ), //i
    .port_byte_in_5  (port_state_in_10_1_5   ), //i
    .port_byte_in_6  (port_state_in_10_1_6   ), //i
    .port_byte_in_7  (port_state_in_10_1_7   ), //i
    .port_byte_out_0 (mul2_54_port_byte_out_0), //o
    .port_byte_out_1 (mul2_54_port_byte_out_1), //o
    .port_byte_out_2 (mul2_54_port_byte_out_2), //o
    .port_byte_out_3 (mul2_54_port_byte_out_3), //o
    .port_byte_out_4 (mul2_54_port_byte_out_4), //o
    .port_byte_out_5 (mul2_54_port_byte_out_5), //o
    .port_byte_out_6 (mul2_54_port_byte_out_6), //o
    .port_byte_out_7 (mul2_54_port_byte_out_7)  //o
  );
  Mul3 mul3_54 (
    .port_byte_in_0  (port_state_in_11_1_0   ), //i
    .port_byte_in_1  (port_state_in_11_1_1   ), //i
    .port_byte_in_2  (port_state_in_11_1_2   ), //i
    .port_byte_in_3  (port_state_in_11_1_3   ), //i
    .port_byte_in_4  (port_state_in_11_1_4   ), //i
    .port_byte_in_5  (port_state_in_11_1_5   ), //i
    .port_byte_in_6  (port_state_in_11_1_6   ), //i
    .port_byte_in_7  (port_state_in_11_1_7   ), //i
    .port_byte_out_0 (mul3_54_port_byte_out_0), //o
    .port_byte_out_1 (mul3_54_port_byte_out_1), //o
    .port_byte_out_2 (mul3_54_port_byte_out_2), //o
    .port_byte_out_3 (mul3_54_port_byte_out_3), //o
    .port_byte_out_4 (mul3_54_port_byte_out_4), //o
    .port_byte_out_5 (mul3_54_port_byte_out_5), //o
    .port_byte_out_6 (mul3_54_port_byte_out_6), //o
    .port_byte_out_7 (mul3_54_port_byte_out_7)  //o
  );
  Mul2 mul2_55 (
    .port_byte_in_0  (port_state_in_11_1_0   ), //i
    .port_byte_in_1  (port_state_in_11_1_1   ), //i
    .port_byte_in_2  (port_state_in_11_1_2   ), //i
    .port_byte_in_3  (port_state_in_11_1_3   ), //i
    .port_byte_in_4  (port_state_in_11_1_4   ), //i
    .port_byte_in_5  (port_state_in_11_1_5   ), //i
    .port_byte_in_6  (port_state_in_11_1_6   ), //i
    .port_byte_in_7  (port_state_in_11_1_7   ), //i
    .port_byte_out_0 (mul2_55_port_byte_out_0), //o
    .port_byte_out_1 (mul2_55_port_byte_out_1), //o
    .port_byte_out_2 (mul2_55_port_byte_out_2), //o
    .port_byte_out_3 (mul2_55_port_byte_out_3), //o
    .port_byte_out_4 (mul2_55_port_byte_out_4), //o
    .port_byte_out_5 (mul2_55_port_byte_out_5), //o
    .port_byte_out_6 (mul2_55_port_byte_out_6), //o
    .port_byte_out_7 (mul2_55_port_byte_out_7)  //o
  );
  Mul3 mul3_55 (
    .port_byte_in_0  (port_state_in_8_1_0    ), //i
    .port_byte_in_1  (port_state_in_8_1_1    ), //i
    .port_byte_in_2  (port_state_in_8_1_2    ), //i
    .port_byte_in_3  (port_state_in_8_1_3    ), //i
    .port_byte_in_4  (port_state_in_8_1_4    ), //i
    .port_byte_in_5  (port_state_in_8_1_5    ), //i
    .port_byte_in_6  (port_state_in_8_1_6    ), //i
    .port_byte_in_7  (port_state_in_8_1_7    ), //i
    .port_byte_out_0 (mul3_55_port_byte_out_0), //o
    .port_byte_out_1 (mul3_55_port_byte_out_1), //o
    .port_byte_out_2 (mul3_55_port_byte_out_2), //o
    .port_byte_out_3 (mul3_55_port_byte_out_3), //o
    .port_byte_out_4 (mul3_55_port_byte_out_4), //o
    .port_byte_out_5 (mul3_55_port_byte_out_5), //o
    .port_byte_out_6 (mul3_55_port_byte_out_6), //o
    .port_byte_out_7 (mul3_55_port_byte_out_7)  //o
  );
  Mul2 mul2_56 (
    .port_byte_in_0  (port_state_in_12_0_0   ), //i
    .port_byte_in_1  (port_state_in_12_0_1   ), //i
    .port_byte_in_2  (port_state_in_12_0_2   ), //i
    .port_byte_in_3  (port_state_in_12_0_3   ), //i
    .port_byte_in_4  (port_state_in_12_0_4   ), //i
    .port_byte_in_5  (port_state_in_12_0_5   ), //i
    .port_byte_in_6  (port_state_in_12_0_6   ), //i
    .port_byte_in_7  (port_state_in_12_0_7   ), //i
    .port_byte_out_0 (mul2_56_port_byte_out_0), //o
    .port_byte_out_1 (mul2_56_port_byte_out_1), //o
    .port_byte_out_2 (mul2_56_port_byte_out_2), //o
    .port_byte_out_3 (mul2_56_port_byte_out_3), //o
    .port_byte_out_4 (mul2_56_port_byte_out_4), //o
    .port_byte_out_5 (mul2_56_port_byte_out_5), //o
    .port_byte_out_6 (mul2_56_port_byte_out_6), //o
    .port_byte_out_7 (mul2_56_port_byte_out_7)  //o
  );
  Mul3 mul3_56 (
    .port_byte_in_0  (port_state_in_13_0_0   ), //i
    .port_byte_in_1  (port_state_in_13_0_1   ), //i
    .port_byte_in_2  (port_state_in_13_0_2   ), //i
    .port_byte_in_3  (port_state_in_13_0_3   ), //i
    .port_byte_in_4  (port_state_in_13_0_4   ), //i
    .port_byte_in_5  (port_state_in_13_0_5   ), //i
    .port_byte_in_6  (port_state_in_13_0_6   ), //i
    .port_byte_in_7  (port_state_in_13_0_7   ), //i
    .port_byte_out_0 (mul3_56_port_byte_out_0), //o
    .port_byte_out_1 (mul3_56_port_byte_out_1), //o
    .port_byte_out_2 (mul3_56_port_byte_out_2), //o
    .port_byte_out_3 (mul3_56_port_byte_out_3), //o
    .port_byte_out_4 (mul3_56_port_byte_out_4), //o
    .port_byte_out_5 (mul3_56_port_byte_out_5), //o
    .port_byte_out_6 (mul3_56_port_byte_out_6), //o
    .port_byte_out_7 (mul3_56_port_byte_out_7)  //o
  );
  Mul2 mul2_57 (
    .port_byte_in_0  (port_state_in_13_0_0   ), //i
    .port_byte_in_1  (port_state_in_13_0_1   ), //i
    .port_byte_in_2  (port_state_in_13_0_2   ), //i
    .port_byte_in_3  (port_state_in_13_0_3   ), //i
    .port_byte_in_4  (port_state_in_13_0_4   ), //i
    .port_byte_in_5  (port_state_in_13_0_5   ), //i
    .port_byte_in_6  (port_state_in_13_0_6   ), //i
    .port_byte_in_7  (port_state_in_13_0_7   ), //i
    .port_byte_out_0 (mul2_57_port_byte_out_0), //o
    .port_byte_out_1 (mul2_57_port_byte_out_1), //o
    .port_byte_out_2 (mul2_57_port_byte_out_2), //o
    .port_byte_out_3 (mul2_57_port_byte_out_3), //o
    .port_byte_out_4 (mul2_57_port_byte_out_4), //o
    .port_byte_out_5 (mul2_57_port_byte_out_5), //o
    .port_byte_out_6 (mul2_57_port_byte_out_6), //o
    .port_byte_out_7 (mul2_57_port_byte_out_7)  //o
  );
  Mul3 mul3_57 (
    .port_byte_in_0  (port_state_in_14_0_0   ), //i
    .port_byte_in_1  (port_state_in_14_0_1   ), //i
    .port_byte_in_2  (port_state_in_14_0_2   ), //i
    .port_byte_in_3  (port_state_in_14_0_3   ), //i
    .port_byte_in_4  (port_state_in_14_0_4   ), //i
    .port_byte_in_5  (port_state_in_14_0_5   ), //i
    .port_byte_in_6  (port_state_in_14_0_6   ), //i
    .port_byte_in_7  (port_state_in_14_0_7   ), //i
    .port_byte_out_0 (mul3_57_port_byte_out_0), //o
    .port_byte_out_1 (mul3_57_port_byte_out_1), //o
    .port_byte_out_2 (mul3_57_port_byte_out_2), //o
    .port_byte_out_3 (mul3_57_port_byte_out_3), //o
    .port_byte_out_4 (mul3_57_port_byte_out_4), //o
    .port_byte_out_5 (mul3_57_port_byte_out_5), //o
    .port_byte_out_6 (mul3_57_port_byte_out_6), //o
    .port_byte_out_7 (mul3_57_port_byte_out_7)  //o
  );
  Mul2 mul2_58 (
    .port_byte_in_0  (port_state_in_14_0_0   ), //i
    .port_byte_in_1  (port_state_in_14_0_1   ), //i
    .port_byte_in_2  (port_state_in_14_0_2   ), //i
    .port_byte_in_3  (port_state_in_14_0_3   ), //i
    .port_byte_in_4  (port_state_in_14_0_4   ), //i
    .port_byte_in_5  (port_state_in_14_0_5   ), //i
    .port_byte_in_6  (port_state_in_14_0_6   ), //i
    .port_byte_in_7  (port_state_in_14_0_7   ), //i
    .port_byte_out_0 (mul2_58_port_byte_out_0), //o
    .port_byte_out_1 (mul2_58_port_byte_out_1), //o
    .port_byte_out_2 (mul2_58_port_byte_out_2), //o
    .port_byte_out_3 (mul2_58_port_byte_out_3), //o
    .port_byte_out_4 (mul2_58_port_byte_out_4), //o
    .port_byte_out_5 (mul2_58_port_byte_out_5), //o
    .port_byte_out_6 (mul2_58_port_byte_out_6), //o
    .port_byte_out_7 (mul2_58_port_byte_out_7)  //o
  );
  Mul3 mul3_58 (
    .port_byte_in_0  (port_state_in_15_0_0   ), //i
    .port_byte_in_1  (port_state_in_15_0_1   ), //i
    .port_byte_in_2  (port_state_in_15_0_2   ), //i
    .port_byte_in_3  (port_state_in_15_0_3   ), //i
    .port_byte_in_4  (port_state_in_15_0_4   ), //i
    .port_byte_in_5  (port_state_in_15_0_5   ), //i
    .port_byte_in_6  (port_state_in_15_0_6   ), //i
    .port_byte_in_7  (port_state_in_15_0_7   ), //i
    .port_byte_out_0 (mul3_58_port_byte_out_0), //o
    .port_byte_out_1 (mul3_58_port_byte_out_1), //o
    .port_byte_out_2 (mul3_58_port_byte_out_2), //o
    .port_byte_out_3 (mul3_58_port_byte_out_3), //o
    .port_byte_out_4 (mul3_58_port_byte_out_4), //o
    .port_byte_out_5 (mul3_58_port_byte_out_5), //o
    .port_byte_out_6 (mul3_58_port_byte_out_6), //o
    .port_byte_out_7 (mul3_58_port_byte_out_7)  //o
  );
  Mul2 mul2_59 (
    .port_byte_in_0  (port_state_in_15_0_0   ), //i
    .port_byte_in_1  (port_state_in_15_0_1   ), //i
    .port_byte_in_2  (port_state_in_15_0_2   ), //i
    .port_byte_in_3  (port_state_in_15_0_3   ), //i
    .port_byte_in_4  (port_state_in_15_0_4   ), //i
    .port_byte_in_5  (port_state_in_15_0_5   ), //i
    .port_byte_in_6  (port_state_in_15_0_6   ), //i
    .port_byte_in_7  (port_state_in_15_0_7   ), //i
    .port_byte_out_0 (mul2_59_port_byte_out_0), //o
    .port_byte_out_1 (mul2_59_port_byte_out_1), //o
    .port_byte_out_2 (mul2_59_port_byte_out_2), //o
    .port_byte_out_3 (mul2_59_port_byte_out_3), //o
    .port_byte_out_4 (mul2_59_port_byte_out_4), //o
    .port_byte_out_5 (mul2_59_port_byte_out_5), //o
    .port_byte_out_6 (mul2_59_port_byte_out_6), //o
    .port_byte_out_7 (mul2_59_port_byte_out_7)  //o
  );
  Mul3 mul3_59 (
    .port_byte_in_0  (port_state_in_12_0_0   ), //i
    .port_byte_in_1  (port_state_in_12_0_1   ), //i
    .port_byte_in_2  (port_state_in_12_0_2   ), //i
    .port_byte_in_3  (port_state_in_12_0_3   ), //i
    .port_byte_in_4  (port_state_in_12_0_4   ), //i
    .port_byte_in_5  (port_state_in_12_0_5   ), //i
    .port_byte_in_6  (port_state_in_12_0_6   ), //i
    .port_byte_in_7  (port_state_in_12_0_7   ), //i
    .port_byte_out_0 (mul3_59_port_byte_out_0), //o
    .port_byte_out_1 (mul3_59_port_byte_out_1), //o
    .port_byte_out_2 (mul3_59_port_byte_out_2), //o
    .port_byte_out_3 (mul3_59_port_byte_out_3), //o
    .port_byte_out_4 (mul3_59_port_byte_out_4), //o
    .port_byte_out_5 (mul3_59_port_byte_out_5), //o
    .port_byte_out_6 (mul3_59_port_byte_out_6), //o
    .port_byte_out_7 (mul3_59_port_byte_out_7)  //o
  );
  Mul2 mul2_60 (
    .port_byte_in_0  (port_state_in_12_1_0   ), //i
    .port_byte_in_1  (port_state_in_12_1_1   ), //i
    .port_byte_in_2  (port_state_in_12_1_2   ), //i
    .port_byte_in_3  (port_state_in_12_1_3   ), //i
    .port_byte_in_4  (port_state_in_12_1_4   ), //i
    .port_byte_in_5  (port_state_in_12_1_5   ), //i
    .port_byte_in_6  (port_state_in_12_1_6   ), //i
    .port_byte_in_7  (port_state_in_12_1_7   ), //i
    .port_byte_out_0 (mul2_60_port_byte_out_0), //o
    .port_byte_out_1 (mul2_60_port_byte_out_1), //o
    .port_byte_out_2 (mul2_60_port_byte_out_2), //o
    .port_byte_out_3 (mul2_60_port_byte_out_3), //o
    .port_byte_out_4 (mul2_60_port_byte_out_4), //o
    .port_byte_out_5 (mul2_60_port_byte_out_5), //o
    .port_byte_out_6 (mul2_60_port_byte_out_6), //o
    .port_byte_out_7 (mul2_60_port_byte_out_7)  //o
  );
  Mul3 mul3_60 (
    .port_byte_in_0  (port_state_in_13_1_0   ), //i
    .port_byte_in_1  (port_state_in_13_1_1   ), //i
    .port_byte_in_2  (port_state_in_13_1_2   ), //i
    .port_byte_in_3  (port_state_in_13_1_3   ), //i
    .port_byte_in_4  (port_state_in_13_1_4   ), //i
    .port_byte_in_5  (port_state_in_13_1_5   ), //i
    .port_byte_in_6  (port_state_in_13_1_6   ), //i
    .port_byte_in_7  (port_state_in_13_1_7   ), //i
    .port_byte_out_0 (mul3_60_port_byte_out_0), //o
    .port_byte_out_1 (mul3_60_port_byte_out_1), //o
    .port_byte_out_2 (mul3_60_port_byte_out_2), //o
    .port_byte_out_3 (mul3_60_port_byte_out_3), //o
    .port_byte_out_4 (mul3_60_port_byte_out_4), //o
    .port_byte_out_5 (mul3_60_port_byte_out_5), //o
    .port_byte_out_6 (mul3_60_port_byte_out_6), //o
    .port_byte_out_7 (mul3_60_port_byte_out_7)  //o
  );
  Mul2 mul2_61 (
    .port_byte_in_0  (port_state_in_13_1_0   ), //i
    .port_byte_in_1  (port_state_in_13_1_1   ), //i
    .port_byte_in_2  (port_state_in_13_1_2   ), //i
    .port_byte_in_3  (port_state_in_13_1_3   ), //i
    .port_byte_in_4  (port_state_in_13_1_4   ), //i
    .port_byte_in_5  (port_state_in_13_1_5   ), //i
    .port_byte_in_6  (port_state_in_13_1_6   ), //i
    .port_byte_in_7  (port_state_in_13_1_7   ), //i
    .port_byte_out_0 (mul2_61_port_byte_out_0), //o
    .port_byte_out_1 (mul2_61_port_byte_out_1), //o
    .port_byte_out_2 (mul2_61_port_byte_out_2), //o
    .port_byte_out_3 (mul2_61_port_byte_out_3), //o
    .port_byte_out_4 (mul2_61_port_byte_out_4), //o
    .port_byte_out_5 (mul2_61_port_byte_out_5), //o
    .port_byte_out_6 (mul2_61_port_byte_out_6), //o
    .port_byte_out_7 (mul2_61_port_byte_out_7)  //o
  );
  Mul3 mul3_61 (
    .port_byte_in_0  (port_state_in_14_1_0   ), //i
    .port_byte_in_1  (port_state_in_14_1_1   ), //i
    .port_byte_in_2  (port_state_in_14_1_2   ), //i
    .port_byte_in_3  (port_state_in_14_1_3   ), //i
    .port_byte_in_4  (port_state_in_14_1_4   ), //i
    .port_byte_in_5  (port_state_in_14_1_5   ), //i
    .port_byte_in_6  (port_state_in_14_1_6   ), //i
    .port_byte_in_7  (port_state_in_14_1_7   ), //i
    .port_byte_out_0 (mul3_61_port_byte_out_0), //o
    .port_byte_out_1 (mul3_61_port_byte_out_1), //o
    .port_byte_out_2 (mul3_61_port_byte_out_2), //o
    .port_byte_out_3 (mul3_61_port_byte_out_3), //o
    .port_byte_out_4 (mul3_61_port_byte_out_4), //o
    .port_byte_out_5 (mul3_61_port_byte_out_5), //o
    .port_byte_out_6 (mul3_61_port_byte_out_6), //o
    .port_byte_out_7 (mul3_61_port_byte_out_7)  //o
  );
  Mul2 mul2_62 (
    .port_byte_in_0  (port_state_in_14_1_0   ), //i
    .port_byte_in_1  (port_state_in_14_1_1   ), //i
    .port_byte_in_2  (port_state_in_14_1_2   ), //i
    .port_byte_in_3  (port_state_in_14_1_3   ), //i
    .port_byte_in_4  (port_state_in_14_1_4   ), //i
    .port_byte_in_5  (port_state_in_14_1_5   ), //i
    .port_byte_in_6  (port_state_in_14_1_6   ), //i
    .port_byte_in_7  (port_state_in_14_1_7   ), //i
    .port_byte_out_0 (mul2_62_port_byte_out_0), //o
    .port_byte_out_1 (mul2_62_port_byte_out_1), //o
    .port_byte_out_2 (mul2_62_port_byte_out_2), //o
    .port_byte_out_3 (mul2_62_port_byte_out_3), //o
    .port_byte_out_4 (mul2_62_port_byte_out_4), //o
    .port_byte_out_5 (mul2_62_port_byte_out_5), //o
    .port_byte_out_6 (mul2_62_port_byte_out_6), //o
    .port_byte_out_7 (mul2_62_port_byte_out_7)  //o
  );
  Mul3 mul3_62 (
    .port_byte_in_0  (port_state_in_15_1_0   ), //i
    .port_byte_in_1  (port_state_in_15_1_1   ), //i
    .port_byte_in_2  (port_state_in_15_1_2   ), //i
    .port_byte_in_3  (port_state_in_15_1_3   ), //i
    .port_byte_in_4  (port_state_in_15_1_4   ), //i
    .port_byte_in_5  (port_state_in_15_1_5   ), //i
    .port_byte_in_6  (port_state_in_15_1_6   ), //i
    .port_byte_in_7  (port_state_in_15_1_7   ), //i
    .port_byte_out_0 (mul3_62_port_byte_out_0), //o
    .port_byte_out_1 (mul3_62_port_byte_out_1), //o
    .port_byte_out_2 (mul3_62_port_byte_out_2), //o
    .port_byte_out_3 (mul3_62_port_byte_out_3), //o
    .port_byte_out_4 (mul3_62_port_byte_out_4), //o
    .port_byte_out_5 (mul3_62_port_byte_out_5), //o
    .port_byte_out_6 (mul3_62_port_byte_out_6), //o
    .port_byte_out_7 (mul3_62_port_byte_out_7)  //o
  );
  Mul2 mul2_63 (
    .port_byte_in_0  (port_state_in_15_1_0   ), //i
    .port_byte_in_1  (port_state_in_15_1_1   ), //i
    .port_byte_in_2  (port_state_in_15_1_2   ), //i
    .port_byte_in_3  (port_state_in_15_1_3   ), //i
    .port_byte_in_4  (port_state_in_15_1_4   ), //i
    .port_byte_in_5  (port_state_in_15_1_5   ), //i
    .port_byte_in_6  (port_state_in_15_1_6   ), //i
    .port_byte_in_7  (port_state_in_15_1_7   ), //i
    .port_byte_out_0 (mul2_63_port_byte_out_0), //o
    .port_byte_out_1 (mul2_63_port_byte_out_1), //o
    .port_byte_out_2 (mul2_63_port_byte_out_2), //o
    .port_byte_out_3 (mul2_63_port_byte_out_3), //o
    .port_byte_out_4 (mul2_63_port_byte_out_4), //o
    .port_byte_out_5 (mul2_63_port_byte_out_5), //o
    .port_byte_out_6 (mul2_63_port_byte_out_6), //o
    .port_byte_out_7 (mul2_63_port_byte_out_7)  //o
  );
  Mul3 mul3_63 (
    .port_byte_in_0  (port_state_in_12_1_0   ), //i
    .port_byte_in_1  (port_state_in_12_1_1   ), //i
    .port_byte_in_2  (port_state_in_12_1_2   ), //i
    .port_byte_in_3  (port_state_in_12_1_3   ), //i
    .port_byte_in_4  (port_state_in_12_1_4   ), //i
    .port_byte_in_5  (port_state_in_12_1_5   ), //i
    .port_byte_in_6  (port_state_in_12_1_6   ), //i
    .port_byte_in_7  (port_state_in_12_1_7   ), //i
    .port_byte_out_0 (mul3_63_port_byte_out_0), //o
    .port_byte_out_1 (mul3_63_port_byte_out_1), //o
    .port_byte_out_2 (mul3_63_port_byte_out_2), //o
    .port_byte_out_3 (mul3_63_port_byte_out_3), //o
    .port_byte_out_4 (mul3_63_port_byte_out_4), //o
    .port_byte_out_5 (mul3_63_port_byte_out_5), //o
    .port_byte_out_6 (mul3_63_port_byte_out_6), //o
    .port_byte_out_7 (mul3_63_port_byte_out_7)  //o
  );
  assign state_out_0_0_0 = (((mul2_32_port_byte_out_0 ^ mul3_32_port_byte_out_0) ^ port_state_in_2_0_0) ^ port_state_in_3_0_0);
  assign state_out_1_0_0 = (((mul2_33_port_byte_out_0 ^ mul3_33_port_byte_out_0) ^ port_state_in_0_0_0) ^ port_state_in_3_0_0);
  assign state_out_2_0_0 = (((mul2_34_port_byte_out_0 ^ mul3_34_port_byte_out_0) ^ port_state_in_0_0_0) ^ port_state_in_1_0_0);
  assign state_out_3_0_0 = (((mul2_35_port_byte_out_0 ^ mul3_35_port_byte_out_0) ^ port_state_in_1_0_0) ^ port_state_in_2_0_0);
  assign state_out_0_0_1 = (((mul2_32_port_byte_out_1 ^ mul3_32_port_byte_out_1) ^ port_state_in_2_0_1) ^ port_state_in_3_0_1);
  assign state_out_1_0_1 = (((mul2_33_port_byte_out_1 ^ mul3_33_port_byte_out_1) ^ port_state_in_0_0_1) ^ port_state_in_3_0_1);
  assign state_out_2_0_1 = (((mul2_34_port_byte_out_1 ^ mul3_34_port_byte_out_1) ^ port_state_in_0_0_1) ^ port_state_in_1_0_1);
  assign state_out_3_0_1 = (((mul2_35_port_byte_out_1 ^ mul3_35_port_byte_out_1) ^ port_state_in_1_0_1) ^ port_state_in_2_0_1);
  assign state_out_0_0_2 = (((mul2_32_port_byte_out_2 ^ mul3_32_port_byte_out_2) ^ port_state_in_2_0_2) ^ port_state_in_3_0_2);
  assign state_out_1_0_2 = (((mul2_33_port_byte_out_2 ^ mul3_33_port_byte_out_2) ^ port_state_in_0_0_2) ^ port_state_in_3_0_2);
  assign state_out_2_0_2 = (((mul2_34_port_byte_out_2 ^ mul3_34_port_byte_out_2) ^ port_state_in_0_0_2) ^ port_state_in_1_0_2);
  assign state_out_3_0_2 = (((mul2_35_port_byte_out_2 ^ mul3_35_port_byte_out_2) ^ port_state_in_1_0_2) ^ port_state_in_2_0_2);
  assign state_out_0_0_3 = (((mul2_32_port_byte_out_3 ^ mul3_32_port_byte_out_3) ^ port_state_in_2_0_3) ^ port_state_in_3_0_3);
  assign state_out_1_0_3 = (((mul2_33_port_byte_out_3 ^ mul3_33_port_byte_out_3) ^ port_state_in_0_0_3) ^ port_state_in_3_0_3);
  assign state_out_2_0_3 = (((mul2_34_port_byte_out_3 ^ mul3_34_port_byte_out_3) ^ port_state_in_0_0_3) ^ port_state_in_1_0_3);
  assign state_out_3_0_3 = (((mul2_35_port_byte_out_3 ^ mul3_35_port_byte_out_3) ^ port_state_in_1_0_3) ^ port_state_in_2_0_3);
  assign state_out_0_0_4 = (((mul2_32_port_byte_out_4 ^ mul3_32_port_byte_out_4) ^ port_state_in_2_0_4) ^ port_state_in_3_0_4);
  assign state_out_1_0_4 = (((mul2_33_port_byte_out_4 ^ mul3_33_port_byte_out_4) ^ port_state_in_0_0_4) ^ port_state_in_3_0_4);
  assign state_out_2_0_4 = (((mul2_34_port_byte_out_4 ^ mul3_34_port_byte_out_4) ^ port_state_in_0_0_4) ^ port_state_in_1_0_4);
  assign state_out_3_0_4 = (((mul2_35_port_byte_out_4 ^ mul3_35_port_byte_out_4) ^ port_state_in_1_0_4) ^ port_state_in_2_0_4);
  assign state_out_0_0_5 = (((mul2_32_port_byte_out_5 ^ mul3_32_port_byte_out_5) ^ port_state_in_2_0_5) ^ port_state_in_3_0_5);
  assign state_out_1_0_5 = (((mul2_33_port_byte_out_5 ^ mul3_33_port_byte_out_5) ^ port_state_in_0_0_5) ^ port_state_in_3_0_5);
  assign state_out_2_0_5 = (((mul2_34_port_byte_out_5 ^ mul3_34_port_byte_out_5) ^ port_state_in_0_0_5) ^ port_state_in_1_0_5);
  assign state_out_3_0_5 = (((mul2_35_port_byte_out_5 ^ mul3_35_port_byte_out_5) ^ port_state_in_1_0_5) ^ port_state_in_2_0_5);
  assign state_out_0_0_6 = (((mul2_32_port_byte_out_6 ^ mul3_32_port_byte_out_6) ^ port_state_in_2_0_6) ^ port_state_in_3_0_6);
  assign state_out_1_0_6 = (((mul2_33_port_byte_out_6 ^ mul3_33_port_byte_out_6) ^ port_state_in_0_0_6) ^ port_state_in_3_0_6);
  assign state_out_2_0_6 = (((mul2_34_port_byte_out_6 ^ mul3_34_port_byte_out_6) ^ port_state_in_0_0_6) ^ port_state_in_1_0_6);
  assign state_out_3_0_6 = (((mul2_35_port_byte_out_6 ^ mul3_35_port_byte_out_6) ^ port_state_in_1_0_6) ^ port_state_in_2_0_6);
  assign state_out_0_0_7 = (((mul2_32_port_byte_out_7 ^ mul3_32_port_byte_out_7) ^ port_state_in_2_0_7) ^ port_state_in_3_0_7);
  assign state_out_1_0_7 = (((mul2_33_port_byte_out_7 ^ mul3_33_port_byte_out_7) ^ port_state_in_0_0_7) ^ port_state_in_3_0_7);
  assign state_out_2_0_7 = (((mul2_34_port_byte_out_7 ^ mul3_34_port_byte_out_7) ^ port_state_in_0_0_7) ^ port_state_in_1_0_7);
  assign state_out_3_0_7 = (((mul2_35_port_byte_out_7 ^ mul3_35_port_byte_out_7) ^ port_state_in_1_0_7) ^ port_state_in_2_0_7);
  assign state_out_0_1_0 = (((mul2_36_port_byte_out_0 ^ mul3_36_port_byte_out_0) ^ port_state_in_2_1_0) ^ port_state_in_3_1_0);
  assign state_out_1_1_0 = (((mul2_37_port_byte_out_0 ^ mul3_37_port_byte_out_0) ^ port_state_in_0_1_0) ^ port_state_in_3_1_0);
  assign state_out_2_1_0 = (((mul2_38_port_byte_out_0 ^ mul3_38_port_byte_out_0) ^ port_state_in_0_1_0) ^ port_state_in_1_1_0);
  assign state_out_3_1_0 = (((mul2_39_port_byte_out_0 ^ mul3_39_port_byte_out_0) ^ port_state_in_1_1_0) ^ port_state_in_2_1_0);
  assign state_out_0_1_1 = (((mul2_36_port_byte_out_1 ^ mul3_36_port_byte_out_1) ^ port_state_in_2_1_1) ^ port_state_in_3_1_1);
  assign state_out_1_1_1 = (((mul2_37_port_byte_out_1 ^ mul3_37_port_byte_out_1) ^ port_state_in_0_1_1) ^ port_state_in_3_1_1);
  assign state_out_2_1_1 = (((mul2_38_port_byte_out_1 ^ mul3_38_port_byte_out_1) ^ port_state_in_0_1_1) ^ port_state_in_1_1_1);
  assign state_out_3_1_1 = (((mul2_39_port_byte_out_1 ^ mul3_39_port_byte_out_1) ^ port_state_in_1_1_1) ^ port_state_in_2_1_1);
  assign state_out_0_1_2 = (((mul2_36_port_byte_out_2 ^ mul3_36_port_byte_out_2) ^ port_state_in_2_1_2) ^ port_state_in_3_1_2);
  assign state_out_1_1_2 = (((mul2_37_port_byte_out_2 ^ mul3_37_port_byte_out_2) ^ port_state_in_0_1_2) ^ port_state_in_3_1_2);
  assign state_out_2_1_2 = (((mul2_38_port_byte_out_2 ^ mul3_38_port_byte_out_2) ^ port_state_in_0_1_2) ^ port_state_in_1_1_2);
  assign state_out_3_1_2 = (((mul2_39_port_byte_out_2 ^ mul3_39_port_byte_out_2) ^ port_state_in_1_1_2) ^ port_state_in_2_1_2);
  assign state_out_0_1_3 = (((mul2_36_port_byte_out_3 ^ mul3_36_port_byte_out_3) ^ port_state_in_2_1_3) ^ port_state_in_3_1_3);
  assign state_out_1_1_3 = (((mul2_37_port_byte_out_3 ^ mul3_37_port_byte_out_3) ^ port_state_in_0_1_3) ^ port_state_in_3_1_3);
  assign state_out_2_1_3 = (((mul2_38_port_byte_out_3 ^ mul3_38_port_byte_out_3) ^ port_state_in_0_1_3) ^ port_state_in_1_1_3);
  assign state_out_3_1_3 = (((mul2_39_port_byte_out_3 ^ mul3_39_port_byte_out_3) ^ port_state_in_1_1_3) ^ port_state_in_2_1_3);
  assign state_out_0_1_4 = (((mul2_36_port_byte_out_4 ^ mul3_36_port_byte_out_4) ^ port_state_in_2_1_4) ^ port_state_in_3_1_4);
  assign state_out_1_1_4 = (((mul2_37_port_byte_out_4 ^ mul3_37_port_byte_out_4) ^ port_state_in_0_1_4) ^ port_state_in_3_1_4);
  assign state_out_2_1_4 = (((mul2_38_port_byte_out_4 ^ mul3_38_port_byte_out_4) ^ port_state_in_0_1_4) ^ port_state_in_1_1_4);
  assign state_out_3_1_4 = (((mul2_39_port_byte_out_4 ^ mul3_39_port_byte_out_4) ^ port_state_in_1_1_4) ^ port_state_in_2_1_4);
  assign state_out_0_1_5 = (((mul2_36_port_byte_out_5 ^ mul3_36_port_byte_out_5) ^ port_state_in_2_1_5) ^ port_state_in_3_1_5);
  assign state_out_1_1_5 = (((mul2_37_port_byte_out_5 ^ mul3_37_port_byte_out_5) ^ port_state_in_0_1_5) ^ port_state_in_3_1_5);
  assign state_out_2_1_5 = (((mul2_38_port_byte_out_5 ^ mul3_38_port_byte_out_5) ^ port_state_in_0_1_5) ^ port_state_in_1_1_5);
  assign state_out_3_1_5 = (((mul2_39_port_byte_out_5 ^ mul3_39_port_byte_out_5) ^ port_state_in_1_1_5) ^ port_state_in_2_1_5);
  assign state_out_0_1_6 = (((mul2_36_port_byte_out_6 ^ mul3_36_port_byte_out_6) ^ port_state_in_2_1_6) ^ port_state_in_3_1_6);
  assign state_out_1_1_6 = (((mul2_37_port_byte_out_6 ^ mul3_37_port_byte_out_6) ^ port_state_in_0_1_6) ^ port_state_in_3_1_6);
  assign state_out_2_1_6 = (((mul2_38_port_byte_out_6 ^ mul3_38_port_byte_out_6) ^ port_state_in_0_1_6) ^ port_state_in_1_1_6);
  assign state_out_3_1_6 = (((mul2_39_port_byte_out_6 ^ mul3_39_port_byte_out_6) ^ port_state_in_1_1_6) ^ port_state_in_2_1_6);
  assign state_out_0_1_7 = (((mul2_36_port_byte_out_7 ^ mul3_36_port_byte_out_7) ^ port_state_in_2_1_7) ^ port_state_in_3_1_7);
  assign state_out_1_1_7 = (((mul2_37_port_byte_out_7 ^ mul3_37_port_byte_out_7) ^ port_state_in_0_1_7) ^ port_state_in_3_1_7);
  assign state_out_2_1_7 = (((mul2_38_port_byte_out_7 ^ mul3_38_port_byte_out_7) ^ port_state_in_0_1_7) ^ port_state_in_1_1_7);
  assign state_out_3_1_7 = (((mul2_39_port_byte_out_7 ^ mul3_39_port_byte_out_7) ^ port_state_in_1_1_7) ^ port_state_in_2_1_7);
  assign state_out_4_0_0 = (((mul2_40_port_byte_out_0 ^ mul3_40_port_byte_out_0) ^ port_state_in_6_0_0) ^ port_state_in_7_0_0);
  assign state_out_5_0_0 = (((mul2_41_port_byte_out_0 ^ mul3_41_port_byte_out_0) ^ port_state_in_4_0_0) ^ port_state_in_7_0_0);
  assign state_out_6_0_0 = (((mul2_42_port_byte_out_0 ^ mul3_42_port_byte_out_0) ^ port_state_in_4_0_0) ^ port_state_in_5_0_0);
  assign state_out_7_0_0 = (((mul2_43_port_byte_out_0 ^ mul3_43_port_byte_out_0) ^ port_state_in_5_0_0) ^ port_state_in_6_0_0);
  assign state_out_4_0_1 = (((mul2_40_port_byte_out_1 ^ mul3_40_port_byte_out_1) ^ port_state_in_6_0_1) ^ port_state_in_7_0_1);
  assign state_out_5_0_1 = (((mul2_41_port_byte_out_1 ^ mul3_41_port_byte_out_1) ^ port_state_in_4_0_1) ^ port_state_in_7_0_1);
  assign state_out_6_0_1 = (((mul2_42_port_byte_out_1 ^ mul3_42_port_byte_out_1) ^ port_state_in_4_0_1) ^ port_state_in_5_0_1);
  assign state_out_7_0_1 = (((mul2_43_port_byte_out_1 ^ mul3_43_port_byte_out_1) ^ port_state_in_5_0_1) ^ port_state_in_6_0_1);
  assign state_out_4_0_2 = (((mul2_40_port_byte_out_2 ^ mul3_40_port_byte_out_2) ^ port_state_in_6_0_2) ^ port_state_in_7_0_2);
  assign state_out_5_0_2 = (((mul2_41_port_byte_out_2 ^ mul3_41_port_byte_out_2) ^ port_state_in_4_0_2) ^ port_state_in_7_0_2);
  assign state_out_6_0_2 = (((mul2_42_port_byte_out_2 ^ mul3_42_port_byte_out_2) ^ port_state_in_4_0_2) ^ port_state_in_5_0_2);
  assign state_out_7_0_2 = (((mul2_43_port_byte_out_2 ^ mul3_43_port_byte_out_2) ^ port_state_in_5_0_2) ^ port_state_in_6_0_2);
  assign state_out_4_0_3 = (((mul2_40_port_byte_out_3 ^ mul3_40_port_byte_out_3) ^ port_state_in_6_0_3) ^ port_state_in_7_0_3);
  assign state_out_5_0_3 = (((mul2_41_port_byte_out_3 ^ mul3_41_port_byte_out_3) ^ port_state_in_4_0_3) ^ port_state_in_7_0_3);
  assign state_out_6_0_3 = (((mul2_42_port_byte_out_3 ^ mul3_42_port_byte_out_3) ^ port_state_in_4_0_3) ^ port_state_in_5_0_3);
  assign state_out_7_0_3 = (((mul2_43_port_byte_out_3 ^ mul3_43_port_byte_out_3) ^ port_state_in_5_0_3) ^ port_state_in_6_0_3);
  assign state_out_4_0_4 = (((mul2_40_port_byte_out_4 ^ mul3_40_port_byte_out_4) ^ port_state_in_6_0_4) ^ port_state_in_7_0_4);
  assign state_out_5_0_4 = (((mul2_41_port_byte_out_4 ^ mul3_41_port_byte_out_4) ^ port_state_in_4_0_4) ^ port_state_in_7_0_4);
  assign state_out_6_0_4 = (((mul2_42_port_byte_out_4 ^ mul3_42_port_byte_out_4) ^ port_state_in_4_0_4) ^ port_state_in_5_0_4);
  assign state_out_7_0_4 = (((mul2_43_port_byte_out_4 ^ mul3_43_port_byte_out_4) ^ port_state_in_5_0_4) ^ port_state_in_6_0_4);
  assign state_out_4_0_5 = (((mul2_40_port_byte_out_5 ^ mul3_40_port_byte_out_5) ^ port_state_in_6_0_5) ^ port_state_in_7_0_5);
  assign state_out_5_0_5 = (((mul2_41_port_byte_out_5 ^ mul3_41_port_byte_out_5) ^ port_state_in_4_0_5) ^ port_state_in_7_0_5);
  assign state_out_6_0_5 = (((mul2_42_port_byte_out_5 ^ mul3_42_port_byte_out_5) ^ port_state_in_4_0_5) ^ port_state_in_5_0_5);
  assign state_out_7_0_5 = (((mul2_43_port_byte_out_5 ^ mul3_43_port_byte_out_5) ^ port_state_in_5_0_5) ^ port_state_in_6_0_5);
  assign state_out_4_0_6 = (((mul2_40_port_byte_out_6 ^ mul3_40_port_byte_out_6) ^ port_state_in_6_0_6) ^ port_state_in_7_0_6);
  assign state_out_5_0_6 = (((mul2_41_port_byte_out_6 ^ mul3_41_port_byte_out_6) ^ port_state_in_4_0_6) ^ port_state_in_7_0_6);
  assign state_out_6_0_6 = (((mul2_42_port_byte_out_6 ^ mul3_42_port_byte_out_6) ^ port_state_in_4_0_6) ^ port_state_in_5_0_6);
  assign state_out_7_0_6 = (((mul2_43_port_byte_out_6 ^ mul3_43_port_byte_out_6) ^ port_state_in_5_0_6) ^ port_state_in_6_0_6);
  assign state_out_4_0_7 = (((mul2_40_port_byte_out_7 ^ mul3_40_port_byte_out_7) ^ port_state_in_6_0_7) ^ port_state_in_7_0_7);
  assign state_out_5_0_7 = (((mul2_41_port_byte_out_7 ^ mul3_41_port_byte_out_7) ^ port_state_in_4_0_7) ^ port_state_in_7_0_7);
  assign state_out_6_0_7 = (((mul2_42_port_byte_out_7 ^ mul3_42_port_byte_out_7) ^ port_state_in_4_0_7) ^ port_state_in_5_0_7);
  assign state_out_7_0_7 = (((mul2_43_port_byte_out_7 ^ mul3_43_port_byte_out_7) ^ port_state_in_5_0_7) ^ port_state_in_6_0_7);
  assign state_out_4_1_0 = (((mul2_44_port_byte_out_0 ^ mul3_44_port_byte_out_0) ^ port_state_in_6_1_0) ^ port_state_in_7_1_0);
  assign state_out_5_1_0 = (((mul2_45_port_byte_out_0 ^ mul3_45_port_byte_out_0) ^ port_state_in_4_1_0) ^ port_state_in_7_1_0);
  assign state_out_6_1_0 = (((mul2_46_port_byte_out_0 ^ mul3_46_port_byte_out_0) ^ port_state_in_4_1_0) ^ port_state_in_5_1_0);
  assign state_out_7_1_0 = (((mul2_47_port_byte_out_0 ^ mul3_47_port_byte_out_0) ^ port_state_in_5_1_0) ^ port_state_in_6_1_0);
  assign state_out_4_1_1 = (((mul2_44_port_byte_out_1 ^ mul3_44_port_byte_out_1) ^ port_state_in_6_1_1) ^ port_state_in_7_1_1);
  assign state_out_5_1_1 = (((mul2_45_port_byte_out_1 ^ mul3_45_port_byte_out_1) ^ port_state_in_4_1_1) ^ port_state_in_7_1_1);
  assign state_out_6_1_1 = (((mul2_46_port_byte_out_1 ^ mul3_46_port_byte_out_1) ^ port_state_in_4_1_1) ^ port_state_in_5_1_1);
  assign state_out_7_1_1 = (((mul2_47_port_byte_out_1 ^ mul3_47_port_byte_out_1) ^ port_state_in_5_1_1) ^ port_state_in_6_1_1);
  assign state_out_4_1_2 = (((mul2_44_port_byte_out_2 ^ mul3_44_port_byte_out_2) ^ port_state_in_6_1_2) ^ port_state_in_7_1_2);
  assign state_out_5_1_2 = (((mul2_45_port_byte_out_2 ^ mul3_45_port_byte_out_2) ^ port_state_in_4_1_2) ^ port_state_in_7_1_2);
  assign state_out_6_1_2 = (((mul2_46_port_byte_out_2 ^ mul3_46_port_byte_out_2) ^ port_state_in_4_1_2) ^ port_state_in_5_1_2);
  assign state_out_7_1_2 = (((mul2_47_port_byte_out_2 ^ mul3_47_port_byte_out_2) ^ port_state_in_5_1_2) ^ port_state_in_6_1_2);
  assign state_out_4_1_3 = (((mul2_44_port_byte_out_3 ^ mul3_44_port_byte_out_3) ^ port_state_in_6_1_3) ^ port_state_in_7_1_3);
  assign state_out_5_1_3 = (((mul2_45_port_byte_out_3 ^ mul3_45_port_byte_out_3) ^ port_state_in_4_1_3) ^ port_state_in_7_1_3);
  assign state_out_6_1_3 = (((mul2_46_port_byte_out_3 ^ mul3_46_port_byte_out_3) ^ port_state_in_4_1_3) ^ port_state_in_5_1_3);
  assign state_out_7_1_3 = (((mul2_47_port_byte_out_3 ^ mul3_47_port_byte_out_3) ^ port_state_in_5_1_3) ^ port_state_in_6_1_3);
  assign state_out_4_1_4 = (((mul2_44_port_byte_out_4 ^ mul3_44_port_byte_out_4) ^ port_state_in_6_1_4) ^ port_state_in_7_1_4);
  assign state_out_5_1_4 = (((mul2_45_port_byte_out_4 ^ mul3_45_port_byte_out_4) ^ port_state_in_4_1_4) ^ port_state_in_7_1_4);
  assign state_out_6_1_4 = (((mul2_46_port_byte_out_4 ^ mul3_46_port_byte_out_4) ^ port_state_in_4_1_4) ^ port_state_in_5_1_4);
  assign state_out_7_1_4 = (((mul2_47_port_byte_out_4 ^ mul3_47_port_byte_out_4) ^ port_state_in_5_1_4) ^ port_state_in_6_1_4);
  assign state_out_4_1_5 = (((mul2_44_port_byte_out_5 ^ mul3_44_port_byte_out_5) ^ port_state_in_6_1_5) ^ port_state_in_7_1_5);
  assign state_out_5_1_5 = (((mul2_45_port_byte_out_5 ^ mul3_45_port_byte_out_5) ^ port_state_in_4_1_5) ^ port_state_in_7_1_5);
  assign state_out_6_1_5 = (((mul2_46_port_byte_out_5 ^ mul3_46_port_byte_out_5) ^ port_state_in_4_1_5) ^ port_state_in_5_1_5);
  assign state_out_7_1_5 = (((mul2_47_port_byte_out_5 ^ mul3_47_port_byte_out_5) ^ port_state_in_5_1_5) ^ port_state_in_6_1_5);
  assign state_out_4_1_6 = (((mul2_44_port_byte_out_6 ^ mul3_44_port_byte_out_6) ^ port_state_in_6_1_6) ^ port_state_in_7_1_6);
  assign state_out_5_1_6 = (((mul2_45_port_byte_out_6 ^ mul3_45_port_byte_out_6) ^ port_state_in_4_1_6) ^ port_state_in_7_1_6);
  assign state_out_6_1_6 = (((mul2_46_port_byte_out_6 ^ mul3_46_port_byte_out_6) ^ port_state_in_4_1_6) ^ port_state_in_5_1_6);
  assign state_out_7_1_6 = (((mul2_47_port_byte_out_6 ^ mul3_47_port_byte_out_6) ^ port_state_in_5_1_6) ^ port_state_in_6_1_6);
  assign state_out_4_1_7 = (((mul2_44_port_byte_out_7 ^ mul3_44_port_byte_out_7) ^ port_state_in_6_1_7) ^ port_state_in_7_1_7);
  assign state_out_5_1_7 = (((mul2_45_port_byte_out_7 ^ mul3_45_port_byte_out_7) ^ port_state_in_4_1_7) ^ port_state_in_7_1_7);
  assign state_out_6_1_7 = (((mul2_46_port_byte_out_7 ^ mul3_46_port_byte_out_7) ^ port_state_in_4_1_7) ^ port_state_in_5_1_7);
  assign state_out_7_1_7 = (((mul2_47_port_byte_out_7 ^ mul3_47_port_byte_out_7) ^ port_state_in_5_1_7) ^ port_state_in_6_1_7);
  assign state_out_8_0_0 = (((mul2_48_port_byte_out_0 ^ mul3_48_port_byte_out_0) ^ port_state_in_10_0_0) ^ port_state_in_11_0_0);
  assign state_out_9_0_0 = (((mul2_49_port_byte_out_0 ^ mul3_49_port_byte_out_0) ^ port_state_in_8_0_0) ^ port_state_in_11_0_0);
  assign state_out_10_0_0 = (((mul2_50_port_byte_out_0 ^ mul3_50_port_byte_out_0) ^ port_state_in_8_0_0) ^ port_state_in_9_0_0);
  assign state_out_11_0_0 = (((mul2_51_port_byte_out_0 ^ mul3_51_port_byte_out_0) ^ port_state_in_9_0_0) ^ port_state_in_10_0_0);
  assign state_out_8_0_1 = (((mul2_48_port_byte_out_1 ^ mul3_48_port_byte_out_1) ^ port_state_in_10_0_1) ^ port_state_in_11_0_1);
  assign state_out_9_0_1 = (((mul2_49_port_byte_out_1 ^ mul3_49_port_byte_out_1) ^ port_state_in_8_0_1) ^ port_state_in_11_0_1);
  assign state_out_10_0_1 = (((mul2_50_port_byte_out_1 ^ mul3_50_port_byte_out_1) ^ port_state_in_8_0_1) ^ port_state_in_9_0_1);
  assign state_out_11_0_1 = (((mul2_51_port_byte_out_1 ^ mul3_51_port_byte_out_1) ^ port_state_in_9_0_1) ^ port_state_in_10_0_1);
  assign state_out_8_0_2 = (((mul2_48_port_byte_out_2 ^ mul3_48_port_byte_out_2) ^ port_state_in_10_0_2) ^ port_state_in_11_0_2);
  assign state_out_9_0_2 = (((mul2_49_port_byte_out_2 ^ mul3_49_port_byte_out_2) ^ port_state_in_8_0_2) ^ port_state_in_11_0_2);
  assign state_out_10_0_2 = (((mul2_50_port_byte_out_2 ^ mul3_50_port_byte_out_2) ^ port_state_in_8_0_2) ^ port_state_in_9_0_2);
  assign state_out_11_0_2 = (((mul2_51_port_byte_out_2 ^ mul3_51_port_byte_out_2) ^ port_state_in_9_0_2) ^ port_state_in_10_0_2);
  assign state_out_8_0_3 = (((mul2_48_port_byte_out_3 ^ mul3_48_port_byte_out_3) ^ port_state_in_10_0_3) ^ port_state_in_11_0_3);
  assign state_out_9_0_3 = (((mul2_49_port_byte_out_3 ^ mul3_49_port_byte_out_3) ^ port_state_in_8_0_3) ^ port_state_in_11_0_3);
  assign state_out_10_0_3 = (((mul2_50_port_byte_out_3 ^ mul3_50_port_byte_out_3) ^ port_state_in_8_0_3) ^ port_state_in_9_0_3);
  assign state_out_11_0_3 = (((mul2_51_port_byte_out_3 ^ mul3_51_port_byte_out_3) ^ port_state_in_9_0_3) ^ port_state_in_10_0_3);
  assign state_out_8_0_4 = (((mul2_48_port_byte_out_4 ^ mul3_48_port_byte_out_4) ^ port_state_in_10_0_4) ^ port_state_in_11_0_4);
  assign state_out_9_0_4 = (((mul2_49_port_byte_out_4 ^ mul3_49_port_byte_out_4) ^ port_state_in_8_0_4) ^ port_state_in_11_0_4);
  assign state_out_10_0_4 = (((mul2_50_port_byte_out_4 ^ mul3_50_port_byte_out_4) ^ port_state_in_8_0_4) ^ port_state_in_9_0_4);
  assign state_out_11_0_4 = (((mul2_51_port_byte_out_4 ^ mul3_51_port_byte_out_4) ^ port_state_in_9_0_4) ^ port_state_in_10_0_4);
  assign state_out_8_0_5 = (((mul2_48_port_byte_out_5 ^ mul3_48_port_byte_out_5) ^ port_state_in_10_0_5) ^ port_state_in_11_0_5);
  assign state_out_9_0_5 = (((mul2_49_port_byte_out_5 ^ mul3_49_port_byte_out_5) ^ port_state_in_8_0_5) ^ port_state_in_11_0_5);
  assign state_out_10_0_5 = (((mul2_50_port_byte_out_5 ^ mul3_50_port_byte_out_5) ^ port_state_in_8_0_5) ^ port_state_in_9_0_5);
  assign state_out_11_0_5 = (((mul2_51_port_byte_out_5 ^ mul3_51_port_byte_out_5) ^ port_state_in_9_0_5) ^ port_state_in_10_0_5);
  assign state_out_8_0_6 = (((mul2_48_port_byte_out_6 ^ mul3_48_port_byte_out_6) ^ port_state_in_10_0_6) ^ port_state_in_11_0_6);
  assign state_out_9_0_6 = (((mul2_49_port_byte_out_6 ^ mul3_49_port_byte_out_6) ^ port_state_in_8_0_6) ^ port_state_in_11_0_6);
  assign state_out_10_0_6 = (((mul2_50_port_byte_out_6 ^ mul3_50_port_byte_out_6) ^ port_state_in_8_0_6) ^ port_state_in_9_0_6);
  assign state_out_11_0_6 = (((mul2_51_port_byte_out_6 ^ mul3_51_port_byte_out_6) ^ port_state_in_9_0_6) ^ port_state_in_10_0_6);
  assign state_out_8_0_7 = (((mul2_48_port_byte_out_7 ^ mul3_48_port_byte_out_7) ^ port_state_in_10_0_7) ^ port_state_in_11_0_7);
  assign state_out_9_0_7 = (((mul2_49_port_byte_out_7 ^ mul3_49_port_byte_out_7) ^ port_state_in_8_0_7) ^ port_state_in_11_0_7);
  assign state_out_10_0_7 = (((mul2_50_port_byte_out_7 ^ mul3_50_port_byte_out_7) ^ port_state_in_8_0_7) ^ port_state_in_9_0_7);
  assign state_out_11_0_7 = (((mul2_51_port_byte_out_7 ^ mul3_51_port_byte_out_7) ^ port_state_in_9_0_7) ^ port_state_in_10_0_7);
  assign state_out_8_1_0 = (((mul2_52_port_byte_out_0 ^ mul3_52_port_byte_out_0) ^ port_state_in_10_1_0) ^ port_state_in_11_1_0);
  assign state_out_9_1_0 = (((mul2_53_port_byte_out_0 ^ mul3_53_port_byte_out_0) ^ port_state_in_8_1_0) ^ port_state_in_11_1_0);
  assign state_out_10_1_0 = (((mul2_54_port_byte_out_0 ^ mul3_54_port_byte_out_0) ^ port_state_in_8_1_0) ^ port_state_in_9_1_0);
  assign state_out_11_1_0 = (((mul2_55_port_byte_out_0 ^ mul3_55_port_byte_out_0) ^ port_state_in_9_1_0) ^ port_state_in_10_1_0);
  assign state_out_8_1_1 = (((mul2_52_port_byte_out_1 ^ mul3_52_port_byte_out_1) ^ port_state_in_10_1_1) ^ port_state_in_11_1_1);
  assign state_out_9_1_1 = (((mul2_53_port_byte_out_1 ^ mul3_53_port_byte_out_1) ^ port_state_in_8_1_1) ^ port_state_in_11_1_1);
  assign state_out_10_1_1 = (((mul2_54_port_byte_out_1 ^ mul3_54_port_byte_out_1) ^ port_state_in_8_1_1) ^ port_state_in_9_1_1);
  assign state_out_11_1_1 = (((mul2_55_port_byte_out_1 ^ mul3_55_port_byte_out_1) ^ port_state_in_9_1_1) ^ port_state_in_10_1_1);
  assign state_out_8_1_2 = (((mul2_52_port_byte_out_2 ^ mul3_52_port_byte_out_2) ^ port_state_in_10_1_2) ^ port_state_in_11_1_2);
  assign state_out_9_1_2 = (((mul2_53_port_byte_out_2 ^ mul3_53_port_byte_out_2) ^ port_state_in_8_1_2) ^ port_state_in_11_1_2);
  assign state_out_10_1_2 = (((mul2_54_port_byte_out_2 ^ mul3_54_port_byte_out_2) ^ port_state_in_8_1_2) ^ port_state_in_9_1_2);
  assign state_out_11_1_2 = (((mul2_55_port_byte_out_2 ^ mul3_55_port_byte_out_2) ^ port_state_in_9_1_2) ^ port_state_in_10_1_2);
  assign state_out_8_1_3 = (((mul2_52_port_byte_out_3 ^ mul3_52_port_byte_out_3) ^ port_state_in_10_1_3) ^ port_state_in_11_1_3);
  assign state_out_9_1_3 = (((mul2_53_port_byte_out_3 ^ mul3_53_port_byte_out_3) ^ port_state_in_8_1_3) ^ port_state_in_11_1_3);
  assign state_out_10_1_3 = (((mul2_54_port_byte_out_3 ^ mul3_54_port_byte_out_3) ^ port_state_in_8_1_3) ^ port_state_in_9_1_3);
  assign state_out_11_1_3 = (((mul2_55_port_byte_out_3 ^ mul3_55_port_byte_out_3) ^ port_state_in_9_1_3) ^ port_state_in_10_1_3);
  assign state_out_8_1_4 = (((mul2_52_port_byte_out_4 ^ mul3_52_port_byte_out_4) ^ port_state_in_10_1_4) ^ port_state_in_11_1_4);
  assign state_out_9_1_4 = (((mul2_53_port_byte_out_4 ^ mul3_53_port_byte_out_4) ^ port_state_in_8_1_4) ^ port_state_in_11_1_4);
  assign state_out_10_1_4 = (((mul2_54_port_byte_out_4 ^ mul3_54_port_byte_out_4) ^ port_state_in_8_1_4) ^ port_state_in_9_1_4);
  assign state_out_11_1_4 = (((mul2_55_port_byte_out_4 ^ mul3_55_port_byte_out_4) ^ port_state_in_9_1_4) ^ port_state_in_10_1_4);
  assign state_out_8_1_5 = (((mul2_52_port_byte_out_5 ^ mul3_52_port_byte_out_5) ^ port_state_in_10_1_5) ^ port_state_in_11_1_5);
  assign state_out_9_1_5 = (((mul2_53_port_byte_out_5 ^ mul3_53_port_byte_out_5) ^ port_state_in_8_1_5) ^ port_state_in_11_1_5);
  assign state_out_10_1_5 = (((mul2_54_port_byte_out_5 ^ mul3_54_port_byte_out_5) ^ port_state_in_8_1_5) ^ port_state_in_9_1_5);
  assign state_out_11_1_5 = (((mul2_55_port_byte_out_5 ^ mul3_55_port_byte_out_5) ^ port_state_in_9_1_5) ^ port_state_in_10_1_5);
  assign state_out_8_1_6 = (((mul2_52_port_byte_out_6 ^ mul3_52_port_byte_out_6) ^ port_state_in_10_1_6) ^ port_state_in_11_1_6);
  assign state_out_9_1_6 = (((mul2_53_port_byte_out_6 ^ mul3_53_port_byte_out_6) ^ port_state_in_8_1_6) ^ port_state_in_11_1_6);
  assign state_out_10_1_6 = (((mul2_54_port_byte_out_6 ^ mul3_54_port_byte_out_6) ^ port_state_in_8_1_6) ^ port_state_in_9_1_6);
  assign state_out_11_1_6 = (((mul2_55_port_byte_out_6 ^ mul3_55_port_byte_out_6) ^ port_state_in_9_1_6) ^ port_state_in_10_1_6);
  assign state_out_8_1_7 = (((mul2_52_port_byte_out_7 ^ mul3_52_port_byte_out_7) ^ port_state_in_10_1_7) ^ port_state_in_11_1_7);
  assign state_out_9_1_7 = (((mul2_53_port_byte_out_7 ^ mul3_53_port_byte_out_7) ^ port_state_in_8_1_7) ^ port_state_in_11_1_7);
  assign state_out_10_1_7 = (((mul2_54_port_byte_out_7 ^ mul3_54_port_byte_out_7) ^ port_state_in_8_1_7) ^ port_state_in_9_1_7);
  assign state_out_11_1_7 = (((mul2_55_port_byte_out_7 ^ mul3_55_port_byte_out_7) ^ port_state_in_9_1_7) ^ port_state_in_10_1_7);
  assign state_out_12_0_0 = (((mul2_56_port_byte_out_0 ^ mul3_56_port_byte_out_0) ^ port_state_in_14_0_0) ^ port_state_in_15_0_0);
  assign state_out_13_0_0 = (((mul2_57_port_byte_out_0 ^ mul3_57_port_byte_out_0) ^ port_state_in_12_0_0) ^ port_state_in_15_0_0);
  assign state_out_14_0_0 = (((mul2_58_port_byte_out_0 ^ mul3_58_port_byte_out_0) ^ port_state_in_12_0_0) ^ port_state_in_13_0_0);
  assign state_out_15_0_0 = (((mul2_59_port_byte_out_0 ^ mul3_59_port_byte_out_0) ^ port_state_in_13_0_0) ^ port_state_in_14_0_0);
  assign state_out_12_0_1 = (((mul2_56_port_byte_out_1 ^ mul3_56_port_byte_out_1) ^ port_state_in_14_0_1) ^ port_state_in_15_0_1);
  assign state_out_13_0_1 = (((mul2_57_port_byte_out_1 ^ mul3_57_port_byte_out_1) ^ port_state_in_12_0_1) ^ port_state_in_15_0_1);
  assign state_out_14_0_1 = (((mul2_58_port_byte_out_1 ^ mul3_58_port_byte_out_1) ^ port_state_in_12_0_1) ^ port_state_in_13_0_1);
  assign state_out_15_0_1 = (((mul2_59_port_byte_out_1 ^ mul3_59_port_byte_out_1) ^ port_state_in_13_0_1) ^ port_state_in_14_0_1);
  assign state_out_12_0_2 = (((mul2_56_port_byte_out_2 ^ mul3_56_port_byte_out_2) ^ port_state_in_14_0_2) ^ port_state_in_15_0_2);
  assign state_out_13_0_2 = (((mul2_57_port_byte_out_2 ^ mul3_57_port_byte_out_2) ^ port_state_in_12_0_2) ^ port_state_in_15_0_2);
  assign state_out_14_0_2 = (((mul2_58_port_byte_out_2 ^ mul3_58_port_byte_out_2) ^ port_state_in_12_0_2) ^ port_state_in_13_0_2);
  assign state_out_15_0_2 = (((mul2_59_port_byte_out_2 ^ mul3_59_port_byte_out_2) ^ port_state_in_13_0_2) ^ port_state_in_14_0_2);
  assign state_out_12_0_3 = (((mul2_56_port_byte_out_3 ^ mul3_56_port_byte_out_3) ^ port_state_in_14_0_3) ^ port_state_in_15_0_3);
  assign state_out_13_0_3 = (((mul2_57_port_byte_out_3 ^ mul3_57_port_byte_out_3) ^ port_state_in_12_0_3) ^ port_state_in_15_0_3);
  assign state_out_14_0_3 = (((mul2_58_port_byte_out_3 ^ mul3_58_port_byte_out_3) ^ port_state_in_12_0_3) ^ port_state_in_13_0_3);
  assign state_out_15_0_3 = (((mul2_59_port_byte_out_3 ^ mul3_59_port_byte_out_3) ^ port_state_in_13_0_3) ^ port_state_in_14_0_3);
  assign state_out_12_0_4 = (((mul2_56_port_byte_out_4 ^ mul3_56_port_byte_out_4) ^ port_state_in_14_0_4) ^ port_state_in_15_0_4);
  assign state_out_13_0_4 = (((mul2_57_port_byte_out_4 ^ mul3_57_port_byte_out_4) ^ port_state_in_12_0_4) ^ port_state_in_15_0_4);
  assign state_out_14_0_4 = (((mul2_58_port_byte_out_4 ^ mul3_58_port_byte_out_4) ^ port_state_in_12_0_4) ^ port_state_in_13_0_4);
  assign state_out_15_0_4 = (((mul2_59_port_byte_out_4 ^ mul3_59_port_byte_out_4) ^ port_state_in_13_0_4) ^ port_state_in_14_0_4);
  assign state_out_12_0_5 = (((mul2_56_port_byte_out_5 ^ mul3_56_port_byte_out_5) ^ port_state_in_14_0_5) ^ port_state_in_15_0_5);
  assign state_out_13_0_5 = (((mul2_57_port_byte_out_5 ^ mul3_57_port_byte_out_5) ^ port_state_in_12_0_5) ^ port_state_in_15_0_5);
  assign state_out_14_0_5 = (((mul2_58_port_byte_out_5 ^ mul3_58_port_byte_out_5) ^ port_state_in_12_0_5) ^ port_state_in_13_0_5);
  assign state_out_15_0_5 = (((mul2_59_port_byte_out_5 ^ mul3_59_port_byte_out_5) ^ port_state_in_13_0_5) ^ port_state_in_14_0_5);
  assign state_out_12_0_6 = (((mul2_56_port_byte_out_6 ^ mul3_56_port_byte_out_6) ^ port_state_in_14_0_6) ^ port_state_in_15_0_6);
  assign state_out_13_0_6 = (((mul2_57_port_byte_out_6 ^ mul3_57_port_byte_out_6) ^ port_state_in_12_0_6) ^ port_state_in_15_0_6);
  assign state_out_14_0_6 = (((mul2_58_port_byte_out_6 ^ mul3_58_port_byte_out_6) ^ port_state_in_12_0_6) ^ port_state_in_13_0_6);
  assign state_out_15_0_6 = (((mul2_59_port_byte_out_6 ^ mul3_59_port_byte_out_6) ^ port_state_in_13_0_6) ^ port_state_in_14_0_6);
  assign state_out_12_0_7 = (((mul2_56_port_byte_out_7 ^ mul3_56_port_byte_out_7) ^ port_state_in_14_0_7) ^ port_state_in_15_0_7);
  assign state_out_13_0_7 = (((mul2_57_port_byte_out_7 ^ mul3_57_port_byte_out_7) ^ port_state_in_12_0_7) ^ port_state_in_15_0_7);
  assign state_out_14_0_7 = (((mul2_58_port_byte_out_7 ^ mul3_58_port_byte_out_7) ^ port_state_in_12_0_7) ^ port_state_in_13_0_7);
  assign state_out_15_0_7 = (((mul2_59_port_byte_out_7 ^ mul3_59_port_byte_out_7) ^ port_state_in_13_0_7) ^ port_state_in_14_0_7);
  assign state_out_12_1_0 = (((mul2_60_port_byte_out_0 ^ mul3_60_port_byte_out_0) ^ port_state_in_14_1_0) ^ port_state_in_15_1_0);
  assign state_out_13_1_0 = (((mul2_61_port_byte_out_0 ^ mul3_61_port_byte_out_0) ^ port_state_in_12_1_0) ^ port_state_in_15_1_0);
  assign state_out_14_1_0 = (((mul2_62_port_byte_out_0 ^ mul3_62_port_byte_out_0) ^ port_state_in_12_1_0) ^ port_state_in_13_1_0);
  assign state_out_15_1_0 = (((mul2_63_port_byte_out_0 ^ mul3_63_port_byte_out_0) ^ port_state_in_13_1_0) ^ port_state_in_14_1_0);
  assign state_out_12_1_1 = (((mul2_60_port_byte_out_1 ^ mul3_60_port_byte_out_1) ^ port_state_in_14_1_1) ^ port_state_in_15_1_1);
  assign state_out_13_1_1 = (((mul2_61_port_byte_out_1 ^ mul3_61_port_byte_out_1) ^ port_state_in_12_1_1) ^ port_state_in_15_1_1);
  assign state_out_14_1_1 = (((mul2_62_port_byte_out_1 ^ mul3_62_port_byte_out_1) ^ port_state_in_12_1_1) ^ port_state_in_13_1_1);
  assign state_out_15_1_1 = (((mul2_63_port_byte_out_1 ^ mul3_63_port_byte_out_1) ^ port_state_in_13_1_1) ^ port_state_in_14_1_1);
  assign state_out_12_1_2 = (((mul2_60_port_byte_out_2 ^ mul3_60_port_byte_out_2) ^ port_state_in_14_1_2) ^ port_state_in_15_1_2);
  assign state_out_13_1_2 = (((mul2_61_port_byte_out_2 ^ mul3_61_port_byte_out_2) ^ port_state_in_12_1_2) ^ port_state_in_15_1_2);
  assign state_out_14_1_2 = (((mul2_62_port_byte_out_2 ^ mul3_62_port_byte_out_2) ^ port_state_in_12_1_2) ^ port_state_in_13_1_2);
  assign state_out_15_1_2 = (((mul2_63_port_byte_out_2 ^ mul3_63_port_byte_out_2) ^ port_state_in_13_1_2) ^ port_state_in_14_1_2);
  assign state_out_12_1_3 = (((mul2_60_port_byte_out_3 ^ mul3_60_port_byte_out_3) ^ port_state_in_14_1_3) ^ port_state_in_15_1_3);
  assign state_out_13_1_3 = (((mul2_61_port_byte_out_3 ^ mul3_61_port_byte_out_3) ^ port_state_in_12_1_3) ^ port_state_in_15_1_3);
  assign state_out_14_1_3 = (((mul2_62_port_byte_out_3 ^ mul3_62_port_byte_out_3) ^ port_state_in_12_1_3) ^ port_state_in_13_1_3);
  assign state_out_15_1_3 = (((mul2_63_port_byte_out_3 ^ mul3_63_port_byte_out_3) ^ port_state_in_13_1_3) ^ port_state_in_14_1_3);
  assign state_out_12_1_4 = (((mul2_60_port_byte_out_4 ^ mul3_60_port_byte_out_4) ^ port_state_in_14_1_4) ^ port_state_in_15_1_4);
  assign state_out_13_1_4 = (((mul2_61_port_byte_out_4 ^ mul3_61_port_byte_out_4) ^ port_state_in_12_1_4) ^ port_state_in_15_1_4);
  assign state_out_14_1_4 = (((mul2_62_port_byte_out_4 ^ mul3_62_port_byte_out_4) ^ port_state_in_12_1_4) ^ port_state_in_13_1_4);
  assign state_out_15_1_4 = (((mul2_63_port_byte_out_4 ^ mul3_63_port_byte_out_4) ^ port_state_in_13_1_4) ^ port_state_in_14_1_4);
  assign state_out_12_1_5 = (((mul2_60_port_byte_out_5 ^ mul3_60_port_byte_out_5) ^ port_state_in_14_1_5) ^ port_state_in_15_1_5);
  assign state_out_13_1_5 = (((mul2_61_port_byte_out_5 ^ mul3_61_port_byte_out_5) ^ port_state_in_12_1_5) ^ port_state_in_15_1_5);
  assign state_out_14_1_5 = (((mul2_62_port_byte_out_5 ^ mul3_62_port_byte_out_5) ^ port_state_in_12_1_5) ^ port_state_in_13_1_5);
  assign state_out_15_1_5 = (((mul2_63_port_byte_out_5 ^ mul3_63_port_byte_out_5) ^ port_state_in_13_1_5) ^ port_state_in_14_1_5);
  assign state_out_12_1_6 = (((mul2_60_port_byte_out_6 ^ mul3_60_port_byte_out_6) ^ port_state_in_14_1_6) ^ port_state_in_15_1_6);
  assign state_out_13_1_6 = (((mul2_61_port_byte_out_6 ^ mul3_61_port_byte_out_6) ^ port_state_in_12_1_6) ^ port_state_in_15_1_6);
  assign state_out_14_1_6 = (((mul2_62_port_byte_out_6 ^ mul3_62_port_byte_out_6) ^ port_state_in_12_1_6) ^ port_state_in_13_1_6);
  assign state_out_15_1_6 = (((mul2_63_port_byte_out_6 ^ mul3_63_port_byte_out_6) ^ port_state_in_13_1_6) ^ port_state_in_14_1_6);
  assign state_out_12_1_7 = (((mul2_60_port_byte_out_7 ^ mul3_60_port_byte_out_7) ^ port_state_in_14_1_7) ^ port_state_in_15_1_7);
  assign state_out_13_1_7 = (((mul2_61_port_byte_out_7 ^ mul3_61_port_byte_out_7) ^ port_state_in_12_1_7) ^ port_state_in_15_1_7);
  assign state_out_14_1_7 = (((mul2_62_port_byte_out_7 ^ mul3_62_port_byte_out_7) ^ port_state_in_12_1_7) ^ port_state_in_13_1_7);
  assign state_out_15_1_7 = (((mul2_63_port_byte_out_7 ^ mul3_63_port_byte_out_7) ^ port_state_in_13_1_7) ^ port_state_in_14_1_7);
  assign port_state_out_0_0_0 = state_out_0_0_0;
  assign port_state_out_0_0_1 = state_out_0_0_1;
  assign port_state_out_0_0_2 = state_out_0_0_2;
  assign port_state_out_0_0_3 = state_out_0_0_3;
  assign port_state_out_0_0_4 = state_out_0_0_4;
  assign port_state_out_0_0_5 = state_out_0_0_5;
  assign port_state_out_0_0_6 = state_out_0_0_6;
  assign port_state_out_0_0_7 = state_out_0_0_7;
  assign port_state_out_0_1_0 = state_out_0_1_0;
  assign port_state_out_0_1_1 = state_out_0_1_1;
  assign port_state_out_0_1_2 = state_out_0_1_2;
  assign port_state_out_0_1_3 = state_out_0_1_3;
  assign port_state_out_0_1_4 = state_out_0_1_4;
  assign port_state_out_0_1_5 = state_out_0_1_5;
  assign port_state_out_0_1_6 = state_out_0_1_6;
  assign port_state_out_0_1_7 = state_out_0_1_7;
  assign port_state_out_1_0_0 = state_out_1_0_0;
  assign port_state_out_1_0_1 = state_out_1_0_1;
  assign port_state_out_1_0_2 = state_out_1_0_2;
  assign port_state_out_1_0_3 = state_out_1_0_3;
  assign port_state_out_1_0_4 = state_out_1_0_4;
  assign port_state_out_1_0_5 = state_out_1_0_5;
  assign port_state_out_1_0_6 = state_out_1_0_6;
  assign port_state_out_1_0_7 = state_out_1_0_7;
  assign port_state_out_1_1_0 = state_out_1_1_0;
  assign port_state_out_1_1_1 = state_out_1_1_1;
  assign port_state_out_1_1_2 = state_out_1_1_2;
  assign port_state_out_1_1_3 = state_out_1_1_3;
  assign port_state_out_1_1_4 = state_out_1_1_4;
  assign port_state_out_1_1_5 = state_out_1_1_5;
  assign port_state_out_1_1_6 = state_out_1_1_6;
  assign port_state_out_1_1_7 = state_out_1_1_7;
  assign port_state_out_2_0_0 = state_out_2_0_0;
  assign port_state_out_2_0_1 = state_out_2_0_1;
  assign port_state_out_2_0_2 = state_out_2_0_2;
  assign port_state_out_2_0_3 = state_out_2_0_3;
  assign port_state_out_2_0_4 = state_out_2_0_4;
  assign port_state_out_2_0_5 = state_out_2_0_5;
  assign port_state_out_2_0_6 = state_out_2_0_6;
  assign port_state_out_2_0_7 = state_out_2_0_7;
  assign port_state_out_2_1_0 = state_out_2_1_0;
  assign port_state_out_2_1_1 = state_out_2_1_1;
  assign port_state_out_2_1_2 = state_out_2_1_2;
  assign port_state_out_2_1_3 = state_out_2_1_3;
  assign port_state_out_2_1_4 = state_out_2_1_4;
  assign port_state_out_2_1_5 = state_out_2_1_5;
  assign port_state_out_2_1_6 = state_out_2_1_6;
  assign port_state_out_2_1_7 = state_out_2_1_7;
  assign port_state_out_3_0_0 = state_out_3_0_0;
  assign port_state_out_3_0_1 = state_out_3_0_1;
  assign port_state_out_3_0_2 = state_out_3_0_2;
  assign port_state_out_3_0_3 = state_out_3_0_3;
  assign port_state_out_3_0_4 = state_out_3_0_4;
  assign port_state_out_3_0_5 = state_out_3_0_5;
  assign port_state_out_3_0_6 = state_out_3_0_6;
  assign port_state_out_3_0_7 = state_out_3_0_7;
  assign port_state_out_3_1_0 = state_out_3_1_0;
  assign port_state_out_3_1_1 = state_out_3_1_1;
  assign port_state_out_3_1_2 = state_out_3_1_2;
  assign port_state_out_3_1_3 = state_out_3_1_3;
  assign port_state_out_3_1_4 = state_out_3_1_4;
  assign port_state_out_3_1_5 = state_out_3_1_5;
  assign port_state_out_3_1_6 = state_out_3_1_6;
  assign port_state_out_3_1_7 = state_out_3_1_7;
  assign port_state_out_4_0_0 = state_out_4_0_0;
  assign port_state_out_4_0_1 = state_out_4_0_1;
  assign port_state_out_4_0_2 = state_out_4_0_2;
  assign port_state_out_4_0_3 = state_out_4_0_3;
  assign port_state_out_4_0_4 = state_out_4_0_4;
  assign port_state_out_4_0_5 = state_out_4_0_5;
  assign port_state_out_4_0_6 = state_out_4_0_6;
  assign port_state_out_4_0_7 = state_out_4_0_7;
  assign port_state_out_4_1_0 = state_out_4_1_0;
  assign port_state_out_4_1_1 = state_out_4_1_1;
  assign port_state_out_4_1_2 = state_out_4_1_2;
  assign port_state_out_4_1_3 = state_out_4_1_3;
  assign port_state_out_4_1_4 = state_out_4_1_4;
  assign port_state_out_4_1_5 = state_out_4_1_5;
  assign port_state_out_4_1_6 = state_out_4_1_6;
  assign port_state_out_4_1_7 = state_out_4_1_7;
  assign port_state_out_5_0_0 = state_out_5_0_0;
  assign port_state_out_5_0_1 = state_out_5_0_1;
  assign port_state_out_5_0_2 = state_out_5_0_2;
  assign port_state_out_5_0_3 = state_out_5_0_3;
  assign port_state_out_5_0_4 = state_out_5_0_4;
  assign port_state_out_5_0_5 = state_out_5_0_5;
  assign port_state_out_5_0_6 = state_out_5_0_6;
  assign port_state_out_5_0_7 = state_out_5_0_7;
  assign port_state_out_5_1_0 = state_out_5_1_0;
  assign port_state_out_5_1_1 = state_out_5_1_1;
  assign port_state_out_5_1_2 = state_out_5_1_2;
  assign port_state_out_5_1_3 = state_out_5_1_3;
  assign port_state_out_5_1_4 = state_out_5_1_4;
  assign port_state_out_5_1_5 = state_out_5_1_5;
  assign port_state_out_5_1_6 = state_out_5_1_6;
  assign port_state_out_5_1_7 = state_out_5_1_7;
  assign port_state_out_6_0_0 = state_out_6_0_0;
  assign port_state_out_6_0_1 = state_out_6_0_1;
  assign port_state_out_6_0_2 = state_out_6_0_2;
  assign port_state_out_6_0_3 = state_out_6_0_3;
  assign port_state_out_6_0_4 = state_out_6_0_4;
  assign port_state_out_6_0_5 = state_out_6_0_5;
  assign port_state_out_6_0_6 = state_out_6_0_6;
  assign port_state_out_6_0_7 = state_out_6_0_7;
  assign port_state_out_6_1_0 = state_out_6_1_0;
  assign port_state_out_6_1_1 = state_out_6_1_1;
  assign port_state_out_6_1_2 = state_out_6_1_2;
  assign port_state_out_6_1_3 = state_out_6_1_3;
  assign port_state_out_6_1_4 = state_out_6_1_4;
  assign port_state_out_6_1_5 = state_out_6_1_5;
  assign port_state_out_6_1_6 = state_out_6_1_6;
  assign port_state_out_6_1_7 = state_out_6_1_7;
  assign port_state_out_7_0_0 = state_out_7_0_0;
  assign port_state_out_7_0_1 = state_out_7_0_1;
  assign port_state_out_7_0_2 = state_out_7_0_2;
  assign port_state_out_7_0_3 = state_out_7_0_3;
  assign port_state_out_7_0_4 = state_out_7_0_4;
  assign port_state_out_7_0_5 = state_out_7_0_5;
  assign port_state_out_7_0_6 = state_out_7_0_6;
  assign port_state_out_7_0_7 = state_out_7_0_7;
  assign port_state_out_7_1_0 = state_out_7_1_0;
  assign port_state_out_7_1_1 = state_out_7_1_1;
  assign port_state_out_7_1_2 = state_out_7_1_2;
  assign port_state_out_7_1_3 = state_out_7_1_3;
  assign port_state_out_7_1_4 = state_out_7_1_4;
  assign port_state_out_7_1_5 = state_out_7_1_5;
  assign port_state_out_7_1_6 = state_out_7_1_6;
  assign port_state_out_7_1_7 = state_out_7_1_7;
  assign port_state_out_8_0_0 = state_out_8_0_0;
  assign port_state_out_8_0_1 = state_out_8_0_1;
  assign port_state_out_8_0_2 = state_out_8_0_2;
  assign port_state_out_8_0_3 = state_out_8_0_3;
  assign port_state_out_8_0_4 = state_out_8_0_4;
  assign port_state_out_8_0_5 = state_out_8_0_5;
  assign port_state_out_8_0_6 = state_out_8_0_6;
  assign port_state_out_8_0_7 = state_out_8_0_7;
  assign port_state_out_8_1_0 = state_out_8_1_0;
  assign port_state_out_8_1_1 = state_out_8_1_1;
  assign port_state_out_8_1_2 = state_out_8_1_2;
  assign port_state_out_8_1_3 = state_out_8_1_3;
  assign port_state_out_8_1_4 = state_out_8_1_4;
  assign port_state_out_8_1_5 = state_out_8_1_5;
  assign port_state_out_8_1_6 = state_out_8_1_6;
  assign port_state_out_8_1_7 = state_out_8_1_7;
  assign port_state_out_9_0_0 = state_out_9_0_0;
  assign port_state_out_9_0_1 = state_out_9_0_1;
  assign port_state_out_9_0_2 = state_out_9_0_2;
  assign port_state_out_9_0_3 = state_out_9_0_3;
  assign port_state_out_9_0_4 = state_out_9_0_4;
  assign port_state_out_9_0_5 = state_out_9_0_5;
  assign port_state_out_9_0_6 = state_out_9_0_6;
  assign port_state_out_9_0_7 = state_out_9_0_7;
  assign port_state_out_9_1_0 = state_out_9_1_0;
  assign port_state_out_9_1_1 = state_out_9_1_1;
  assign port_state_out_9_1_2 = state_out_9_1_2;
  assign port_state_out_9_1_3 = state_out_9_1_3;
  assign port_state_out_9_1_4 = state_out_9_1_4;
  assign port_state_out_9_1_5 = state_out_9_1_5;
  assign port_state_out_9_1_6 = state_out_9_1_6;
  assign port_state_out_9_1_7 = state_out_9_1_7;
  assign port_state_out_10_0_0 = state_out_10_0_0;
  assign port_state_out_10_0_1 = state_out_10_0_1;
  assign port_state_out_10_0_2 = state_out_10_0_2;
  assign port_state_out_10_0_3 = state_out_10_0_3;
  assign port_state_out_10_0_4 = state_out_10_0_4;
  assign port_state_out_10_0_5 = state_out_10_0_5;
  assign port_state_out_10_0_6 = state_out_10_0_6;
  assign port_state_out_10_0_7 = state_out_10_0_7;
  assign port_state_out_10_1_0 = state_out_10_1_0;
  assign port_state_out_10_1_1 = state_out_10_1_1;
  assign port_state_out_10_1_2 = state_out_10_1_2;
  assign port_state_out_10_1_3 = state_out_10_1_3;
  assign port_state_out_10_1_4 = state_out_10_1_4;
  assign port_state_out_10_1_5 = state_out_10_1_5;
  assign port_state_out_10_1_6 = state_out_10_1_6;
  assign port_state_out_10_1_7 = state_out_10_1_7;
  assign port_state_out_11_0_0 = state_out_11_0_0;
  assign port_state_out_11_0_1 = state_out_11_0_1;
  assign port_state_out_11_0_2 = state_out_11_0_2;
  assign port_state_out_11_0_3 = state_out_11_0_3;
  assign port_state_out_11_0_4 = state_out_11_0_4;
  assign port_state_out_11_0_5 = state_out_11_0_5;
  assign port_state_out_11_0_6 = state_out_11_0_6;
  assign port_state_out_11_0_7 = state_out_11_0_7;
  assign port_state_out_11_1_0 = state_out_11_1_0;
  assign port_state_out_11_1_1 = state_out_11_1_1;
  assign port_state_out_11_1_2 = state_out_11_1_2;
  assign port_state_out_11_1_3 = state_out_11_1_3;
  assign port_state_out_11_1_4 = state_out_11_1_4;
  assign port_state_out_11_1_5 = state_out_11_1_5;
  assign port_state_out_11_1_6 = state_out_11_1_6;
  assign port_state_out_11_1_7 = state_out_11_1_7;
  assign port_state_out_12_0_0 = state_out_12_0_0;
  assign port_state_out_12_0_1 = state_out_12_0_1;
  assign port_state_out_12_0_2 = state_out_12_0_2;
  assign port_state_out_12_0_3 = state_out_12_0_3;
  assign port_state_out_12_0_4 = state_out_12_0_4;
  assign port_state_out_12_0_5 = state_out_12_0_5;
  assign port_state_out_12_0_6 = state_out_12_0_6;
  assign port_state_out_12_0_7 = state_out_12_0_7;
  assign port_state_out_12_1_0 = state_out_12_1_0;
  assign port_state_out_12_1_1 = state_out_12_1_1;
  assign port_state_out_12_1_2 = state_out_12_1_2;
  assign port_state_out_12_1_3 = state_out_12_1_3;
  assign port_state_out_12_1_4 = state_out_12_1_4;
  assign port_state_out_12_1_5 = state_out_12_1_5;
  assign port_state_out_12_1_6 = state_out_12_1_6;
  assign port_state_out_12_1_7 = state_out_12_1_7;
  assign port_state_out_13_0_0 = state_out_13_0_0;
  assign port_state_out_13_0_1 = state_out_13_0_1;
  assign port_state_out_13_0_2 = state_out_13_0_2;
  assign port_state_out_13_0_3 = state_out_13_0_3;
  assign port_state_out_13_0_4 = state_out_13_0_4;
  assign port_state_out_13_0_5 = state_out_13_0_5;
  assign port_state_out_13_0_6 = state_out_13_0_6;
  assign port_state_out_13_0_7 = state_out_13_0_7;
  assign port_state_out_13_1_0 = state_out_13_1_0;
  assign port_state_out_13_1_1 = state_out_13_1_1;
  assign port_state_out_13_1_2 = state_out_13_1_2;
  assign port_state_out_13_1_3 = state_out_13_1_3;
  assign port_state_out_13_1_4 = state_out_13_1_4;
  assign port_state_out_13_1_5 = state_out_13_1_5;
  assign port_state_out_13_1_6 = state_out_13_1_6;
  assign port_state_out_13_1_7 = state_out_13_1_7;
  assign port_state_out_14_0_0 = state_out_14_0_0;
  assign port_state_out_14_0_1 = state_out_14_0_1;
  assign port_state_out_14_0_2 = state_out_14_0_2;
  assign port_state_out_14_0_3 = state_out_14_0_3;
  assign port_state_out_14_0_4 = state_out_14_0_4;
  assign port_state_out_14_0_5 = state_out_14_0_5;
  assign port_state_out_14_0_6 = state_out_14_0_6;
  assign port_state_out_14_0_7 = state_out_14_0_7;
  assign port_state_out_14_1_0 = state_out_14_1_0;
  assign port_state_out_14_1_1 = state_out_14_1_1;
  assign port_state_out_14_1_2 = state_out_14_1_2;
  assign port_state_out_14_1_3 = state_out_14_1_3;
  assign port_state_out_14_1_4 = state_out_14_1_4;
  assign port_state_out_14_1_5 = state_out_14_1_5;
  assign port_state_out_14_1_6 = state_out_14_1_6;
  assign port_state_out_14_1_7 = state_out_14_1_7;
  assign port_state_out_15_0_0 = state_out_15_0_0;
  assign port_state_out_15_0_1 = state_out_15_0_1;
  assign port_state_out_15_0_2 = state_out_15_0_2;
  assign port_state_out_15_0_3 = state_out_15_0_3;
  assign port_state_out_15_0_4 = state_out_15_0_4;
  assign port_state_out_15_0_5 = state_out_15_0_5;
  assign port_state_out_15_0_6 = state_out_15_0_6;
  assign port_state_out_15_0_7 = state_out_15_0_7;
  assign port_state_out_15_1_0 = state_out_15_1_0;
  assign port_state_out_15_1_1 = state_out_15_1_1;
  assign port_state_out_15_1_2 = state_out_15_1_2;
  assign port_state_out_15_1_3 = state_out_15_1_3;
  assign port_state_out_15_1_4 = state_out_15_1_4;
  assign port_state_out_15_1_5 = state_out_15_1_5;
  assign port_state_out_15_1_6 = state_out_15_1_6;
  assign port_state_out_15_1_7 = state_out_15_1_7;

endmodule

module AES_ShiftRows (
  input      [0:0]    port_state_in_0_0_0,
  input      [0:0]    port_state_in_0_0_1,
  input      [0:0]    port_state_in_0_0_2,
  input      [0:0]    port_state_in_0_0_3,
  input      [0:0]    port_state_in_0_0_4,
  input      [0:0]    port_state_in_0_0_5,
  input      [0:0]    port_state_in_0_0_6,
  input      [0:0]    port_state_in_0_0_7,
  input      [0:0]    port_state_in_0_1_0,
  input      [0:0]    port_state_in_0_1_1,
  input      [0:0]    port_state_in_0_1_2,
  input      [0:0]    port_state_in_0_1_3,
  input      [0:0]    port_state_in_0_1_4,
  input      [0:0]    port_state_in_0_1_5,
  input      [0:0]    port_state_in_0_1_6,
  input      [0:0]    port_state_in_0_1_7,
  input      [0:0]    port_state_in_1_0_0,
  input      [0:0]    port_state_in_1_0_1,
  input      [0:0]    port_state_in_1_0_2,
  input      [0:0]    port_state_in_1_0_3,
  input      [0:0]    port_state_in_1_0_4,
  input      [0:0]    port_state_in_1_0_5,
  input      [0:0]    port_state_in_1_0_6,
  input      [0:0]    port_state_in_1_0_7,
  input      [0:0]    port_state_in_1_1_0,
  input      [0:0]    port_state_in_1_1_1,
  input      [0:0]    port_state_in_1_1_2,
  input      [0:0]    port_state_in_1_1_3,
  input      [0:0]    port_state_in_1_1_4,
  input      [0:0]    port_state_in_1_1_5,
  input      [0:0]    port_state_in_1_1_6,
  input      [0:0]    port_state_in_1_1_7,
  input      [0:0]    port_state_in_2_0_0,
  input      [0:0]    port_state_in_2_0_1,
  input      [0:0]    port_state_in_2_0_2,
  input      [0:0]    port_state_in_2_0_3,
  input      [0:0]    port_state_in_2_0_4,
  input      [0:0]    port_state_in_2_0_5,
  input      [0:0]    port_state_in_2_0_6,
  input      [0:0]    port_state_in_2_0_7,
  input      [0:0]    port_state_in_2_1_0,
  input      [0:0]    port_state_in_2_1_1,
  input      [0:0]    port_state_in_2_1_2,
  input      [0:0]    port_state_in_2_1_3,
  input      [0:0]    port_state_in_2_1_4,
  input      [0:0]    port_state_in_2_1_5,
  input      [0:0]    port_state_in_2_1_6,
  input      [0:0]    port_state_in_2_1_7,
  input      [0:0]    port_state_in_3_0_0,
  input      [0:0]    port_state_in_3_0_1,
  input      [0:0]    port_state_in_3_0_2,
  input      [0:0]    port_state_in_3_0_3,
  input      [0:0]    port_state_in_3_0_4,
  input      [0:0]    port_state_in_3_0_5,
  input      [0:0]    port_state_in_3_0_6,
  input      [0:0]    port_state_in_3_0_7,
  input      [0:0]    port_state_in_3_1_0,
  input      [0:0]    port_state_in_3_1_1,
  input      [0:0]    port_state_in_3_1_2,
  input      [0:0]    port_state_in_3_1_3,
  input      [0:0]    port_state_in_3_1_4,
  input      [0:0]    port_state_in_3_1_5,
  input      [0:0]    port_state_in_3_1_6,
  input      [0:0]    port_state_in_3_1_7,
  input      [0:0]    port_state_in_4_0_0,
  input      [0:0]    port_state_in_4_0_1,
  input      [0:0]    port_state_in_4_0_2,
  input      [0:0]    port_state_in_4_0_3,
  input      [0:0]    port_state_in_4_0_4,
  input      [0:0]    port_state_in_4_0_5,
  input      [0:0]    port_state_in_4_0_6,
  input      [0:0]    port_state_in_4_0_7,
  input      [0:0]    port_state_in_4_1_0,
  input      [0:0]    port_state_in_4_1_1,
  input      [0:0]    port_state_in_4_1_2,
  input      [0:0]    port_state_in_4_1_3,
  input      [0:0]    port_state_in_4_1_4,
  input      [0:0]    port_state_in_4_1_5,
  input      [0:0]    port_state_in_4_1_6,
  input      [0:0]    port_state_in_4_1_7,
  input      [0:0]    port_state_in_5_0_0,
  input      [0:0]    port_state_in_5_0_1,
  input      [0:0]    port_state_in_5_0_2,
  input      [0:0]    port_state_in_5_0_3,
  input      [0:0]    port_state_in_5_0_4,
  input      [0:0]    port_state_in_5_0_5,
  input      [0:0]    port_state_in_5_0_6,
  input      [0:0]    port_state_in_5_0_7,
  input      [0:0]    port_state_in_5_1_0,
  input      [0:0]    port_state_in_5_1_1,
  input      [0:0]    port_state_in_5_1_2,
  input      [0:0]    port_state_in_5_1_3,
  input      [0:0]    port_state_in_5_1_4,
  input      [0:0]    port_state_in_5_1_5,
  input      [0:0]    port_state_in_5_1_6,
  input      [0:0]    port_state_in_5_1_7,
  input      [0:0]    port_state_in_6_0_0,
  input      [0:0]    port_state_in_6_0_1,
  input      [0:0]    port_state_in_6_0_2,
  input      [0:0]    port_state_in_6_0_3,
  input      [0:0]    port_state_in_6_0_4,
  input      [0:0]    port_state_in_6_0_5,
  input      [0:0]    port_state_in_6_0_6,
  input      [0:0]    port_state_in_6_0_7,
  input      [0:0]    port_state_in_6_1_0,
  input      [0:0]    port_state_in_6_1_1,
  input      [0:0]    port_state_in_6_1_2,
  input      [0:0]    port_state_in_6_1_3,
  input      [0:0]    port_state_in_6_1_4,
  input      [0:0]    port_state_in_6_1_5,
  input      [0:0]    port_state_in_6_1_6,
  input      [0:0]    port_state_in_6_1_7,
  input      [0:0]    port_state_in_7_0_0,
  input      [0:0]    port_state_in_7_0_1,
  input      [0:0]    port_state_in_7_0_2,
  input      [0:0]    port_state_in_7_0_3,
  input      [0:0]    port_state_in_7_0_4,
  input      [0:0]    port_state_in_7_0_5,
  input      [0:0]    port_state_in_7_0_6,
  input      [0:0]    port_state_in_7_0_7,
  input      [0:0]    port_state_in_7_1_0,
  input      [0:0]    port_state_in_7_1_1,
  input      [0:0]    port_state_in_7_1_2,
  input      [0:0]    port_state_in_7_1_3,
  input      [0:0]    port_state_in_7_1_4,
  input      [0:0]    port_state_in_7_1_5,
  input      [0:0]    port_state_in_7_1_6,
  input      [0:0]    port_state_in_7_1_7,
  input      [0:0]    port_state_in_8_0_0,
  input      [0:0]    port_state_in_8_0_1,
  input      [0:0]    port_state_in_8_0_2,
  input      [0:0]    port_state_in_8_0_3,
  input      [0:0]    port_state_in_8_0_4,
  input      [0:0]    port_state_in_8_0_5,
  input      [0:0]    port_state_in_8_0_6,
  input      [0:0]    port_state_in_8_0_7,
  input      [0:0]    port_state_in_8_1_0,
  input      [0:0]    port_state_in_8_1_1,
  input      [0:0]    port_state_in_8_1_2,
  input      [0:0]    port_state_in_8_1_3,
  input      [0:0]    port_state_in_8_1_4,
  input      [0:0]    port_state_in_8_1_5,
  input      [0:0]    port_state_in_8_1_6,
  input      [0:0]    port_state_in_8_1_7,
  input      [0:0]    port_state_in_9_0_0,
  input      [0:0]    port_state_in_9_0_1,
  input      [0:0]    port_state_in_9_0_2,
  input      [0:0]    port_state_in_9_0_3,
  input      [0:0]    port_state_in_9_0_4,
  input      [0:0]    port_state_in_9_0_5,
  input      [0:0]    port_state_in_9_0_6,
  input      [0:0]    port_state_in_9_0_7,
  input      [0:0]    port_state_in_9_1_0,
  input      [0:0]    port_state_in_9_1_1,
  input      [0:0]    port_state_in_9_1_2,
  input      [0:0]    port_state_in_9_1_3,
  input      [0:0]    port_state_in_9_1_4,
  input      [0:0]    port_state_in_9_1_5,
  input      [0:0]    port_state_in_9_1_6,
  input      [0:0]    port_state_in_9_1_7,
  input      [0:0]    port_state_in_10_0_0,
  input      [0:0]    port_state_in_10_0_1,
  input      [0:0]    port_state_in_10_0_2,
  input      [0:0]    port_state_in_10_0_3,
  input      [0:0]    port_state_in_10_0_4,
  input      [0:0]    port_state_in_10_0_5,
  input      [0:0]    port_state_in_10_0_6,
  input      [0:0]    port_state_in_10_0_7,
  input      [0:0]    port_state_in_10_1_0,
  input      [0:0]    port_state_in_10_1_1,
  input      [0:0]    port_state_in_10_1_2,
  input      [0:0]    port_state_in_10_1_3,
  input      [0:0]    port_state_in_10_1_4,
  input      [0:0]    port_state_in_10_1_5,
  input      [0:0]    port_state_in_10_1_6,
  input      [0:0]    port_state_in_10_1_7,
  input      [0:0]    port_state_in_11_0_0,
  input      [0:0]    port_state_in_11_0_1,
  input      [0:0]    port_state_in_11_0_2,
  input      [0:0]    port_state_in_11_0_3,
  input      [0:0]    port_state_in_11_0_4,
  input      [0:0]    port_state_in_11_0_5,
  input      [0:0]    port_state_in_11_0_6,
  input      [0:0]    port_state_in_11_0_7,
  input      [0:0]    port_state_in_11_1_0,
  input      [0:0]    port_state_in_11_1_1,
  input      [0:0]    port_state_in_11_1_2,
  input      [0:0]    port_state_in_11_1_3,
  input      [0:0]    port_state_in_11_1_4,
  input      [0:0]    port_state_in_11_1_5,
  input      [0:0]    port_state_in_11_1_6,
  input      [0:0]    port_state_in_11_1_7,
  input      [0:0]    port_state_in_12_0_0,
  input      [0:0]    port_state_in_12_0_1,
  input      [0:0]    port_state_in_12_0_2,
  input      [0:0]    port_state_in_12_0_3,
  input      [0:0]    port_state_in_12_0_4,
  input      [0:0]    port_state_in_12_0_5,
  input      [0:0]    port_state_in_12_0_6,
  input      [0:0]    port_state_in_12_0_7,
  input      [0:0]    port_state_in_12_1_0,
  input      [0:0]    port_state_in_12_1_1,
  input      [0:0]    port_state_in_12_1_2,
  input      [0:0]    port_state_in_12_1_3,
  input      [0:0]    port_state_in_12_1_4,
  input      [0:0]    port_state_in_12_1_5,
  input      [0:0]    port_state_in_12_1_6,
  input      [0:0]    port_state_in_12_1_7,
  input      [0:0]    port_state_in_13_0_0,
  input      [0:0]    port_state_in_13_0_1,
  input      [0:0]    port_state_in_13_0_2,
  input      [0:0]    port_state_in_13_0_3,
  input      [0:0]    port_state_in_13_0_4,
  input      [0:0]    port_state_in_13_0_5,
  input      [0:0]    port_state_in_13_0_6,
  input      [0:0]    port_state_in_13_0_7,
  input      [0:0]    port_state_in_13_1_0,
  input      [0:0]    port_state_in_13_1_1,
  input      [0:0]    port_state_in_13_1_2,
  input      [0:0]    port_state_in_13_1_3,
  input      [0:0]    port_state_in_13_1_4,
  input      [0:0]    port_state_in_13_1_5,
  input      [0:0]    port_state_in_13_1_6,
  input      [0:0]    port_state_in_13_1_7,
  input      [0:0]    port_state_in_14_0_0,
  input      [0:0]    port_state_in_14_0_1,
  input      [0:0]    port_state_in_14_0_2,
  input      [0:0]    port_state_in_14_0_3,
  input      [0:0]    port_state_in_14_0_4,
  input      [0:0]    port_state_in_14_0_5,
  input      [0:0]    port_state_in_14_0_6,
  input      [0:0]    port_state_in_14_0_7,
  input      [0:0]    port_state_in_14_1_0,
  input      [0:0]    port_state_in_14_1_1,
  input      [0:0]    port_state_in_14_1_2,
  input      [0:0]    port_state_in_14_1_3,
  input      [0:0]    port_state_in_14_1_4,
  input      [0:0]    port_state_in_14_1_5,
  input      [0:0]    port_state_in_14_1_6,
  input      [0:0]    port_state_in_14_1_7,
  input      [0:0]    port_state_in_15_0_0,
  input      [0:0]    port_state_in_15_0_1,
  input      [0:0]    port_state_in_15_0_2,
  input      [0:0]    port_state_in_15_0_3,
  input      [0:0]    port_state_in_15_0_4,
  input      [0:0]    port_state_in_15_0_5,
  input      [0:0]    port_state_in_15_0_6,
  input      [0:0]    port_state_in_15_0_7,
  input      [0:0]    port_state_in_15_1_0,
  input      [0:0]    port_state_in_15_1_1,
  input      [0:0]    port_state_in_15_1_2,
  input      [0:0]    port_state_in_15_1_3,
  input      [0:0]    port_state_in_15_1_4,
  input      [0:0]    port_state_in_15_1_5,
  input      [0:0]    port_state_in_15_1_6,
  input      [0:0]    port_state_in_15_1_7,
  output     [0:0]    port_state_out_0_0_0,
  output     [0:0]    port_state_out_0_0_1,
  output     [0:0]    port_state_out_0_0_2,
  output     [0:0]    port_state_out_0_0_3,
  output     [0:0]    port_state_out_0_0_4,
  output     [0:0]    port_state_out_0_0_5,
  output     [0:0]    port_state_out_0_0_6,
  output     [0:0]    port_state_out_0_0_7,
  output     [0:0]    port_state_out_0_1_0,
  output     [0:0]    port_state_out_0_1_1,
  output     [0:0]    port_state_out_0_1_2,
  output     [0:0]    port_state_out_0_1_3,
  output     [0:0]    port_state_out_0_1_4,
  output     [0:0]    port_state_out_0_1_5,
  output     [0:0]    port_state_out_0_1_6,
  output     [0:0]    port_state_out_0_1_7,
  output     [0:0]    port_state_out_1_0_0,
  output     [0:0]    port_state_out_1_0_1,
  output     [0:0]    port_state_out_1_0_2,
  output     [0:0]    port_state_out_1_0_3,
  output     [0:0]    port_state_out_1_0_4,
  output     [0:0]    port_state_out_1_0_5,
  output     [0:0]    port_state_out_1_0_6,
  output     [0:0]    port_state_out_1_0_7,
  output     [0:0]    port_state_out_1_1_0,
  output     [0:0]    port_state_out_1_1_1,
  output     [0:0]    port_state_out_1_1_2,
  output     [0:0]    port_state_out_1_1_3,
  output     [0:0]    port_state_out_1_1_4,
  output     [0:0]    port_state_out_1_1_5,
  output     [0:0]    port_state_out_1_1_6,
  output     [0:0]    port_state_out_1_1_7,
  output     [0:0]    port_state_out_2_0_0,
  output     [0:0]    port_state_out_2_0_1,
  output     [0:0]    port_state_out_2_0_2,
  output     [0:0]    port_state_out_2_0_3,
  output     [0:0]    port_state_out_2_0_4,
  output     [0:0]    port_state_out_2_0_5,
  output     [0:0]    port_state_out_2_0_6,
  output     [0:0]    port_state_out_2_0_7,
  output     [0:0]    port_state_out_2_1_0,
  output     [0:0]    port_state_out_2_1_1,
  output     [0:0]    port_state_out_2_1_2,
  output     [0:0]    port_state_out_2_1_3,
  output     [0:0]    port_state_out_2_1_4,
  output     [0:0]    port_state_out_2_1_5,
  output     [0:0]    port_state_out_2_1_6,
  output     [0:0]    port_state_out_2_1_7,
  output     [0:0]    port_state_out_3_0_0,
  output     [0:0]    port_state_out_3_0_1,
  output     [0:0]    port_state_out_3_0_2,
  output     [0:0]    port_state_out_3_0_3,
  output     [0:0]    port_state_out_3_0_4,
  output     [0:0]    port_state_out_3_0_5,
  output     [0:0]    port_state_out_3_0_6,
  output     [0:0]    port_state_out_3_0_7,
  output     [0:0]    port_state_out_3_1_0,
  output     [0:0]    port_state_out_3_1_1,
  output     [0:0]    port_state_out_3_1_2,
  output     [0:0]    port_state_out_3_1_3,
  output     [0:0]    port_state_out_3_1_4,
  output     [0:0]    port_state_out_3_1_5,
  output     [0:0]    port_state_out_3_1_6,
  output     [0:0]    port_state_out_3_1_7,
  output     [0:0]    port_state_out_4_0_0,
  output     [0:0]    port_state_out_4_0_1,
  output     [0:0]    port_state_out_4_0_2,
  output     [0:0]    port_state_out_4_0_3,
  output     [0:0]    port_state_out_4_0_4,
  output     [0:0]    port_state_out_4_0_5,
  output     [0:0]    port_state_out_4_0_6,
  output     [0:0]    port_state_out_4_0_7,
  output     [0:0]    port_state_out_4_1_0,
  output     [0:0]    port_state_out_4_1_1,
  output     [0:0]    port_state_out_4_1_2,
  output     [0:0]    port_state_out_4_1_3,
  output     [0:0]    port_state_out_4_1_4,
  output     [0:0]    port_state_out_4_1_5,
  output     [0:0]    port_state_out_4_1_6,
  output     [0:0]    port_state_out_4_1_7,
  output     [0:0]    port_state_out_5_0_0,
  output     [0:0]    port_state_out_5_0_1,
  output     [0:0]    port_state_out_5_0_2,
  output     [0:0]    port_state_out_5_0_3,
  output     [0:0]    port_state_out_5_0_4,
  output     [0:0]    port_state_out_5_0_5,
  output     [0:0]    port_state_out_5_0_6,
  output     [0:0]    port_state_out_5_0_7,
  output     [0:0]    port_state_out_5_1_0,
  output     [0:0]    port_state_out_5_1_1,
  output     [0:0]    port_state_out_5_1_2,
  output     [0:0]    port_state_out_5_1_3,
  output     [0:0]    port_state_out_5_1_4,
  output     [0:0]    port_state_out_5_1_5,
  output     [0:0]    port_state_out_5_1_6,
  output     [0:0]    port_state_out_5_1_7,
  output     [0:0]    port_state_out_6_0_0,
  output     [0:0]    port_state_out_6_0_1,
  output     [0:0]    port_state_out_6_0_2,
  output     [0:0]    port_state_out_6_0_3,
  output     [0:0]    port_state_out_6_0_4,
  output     [0:0]    port_state_out_6_0_5,
  output     [0:0]    port_state_out_6_0_6,
  output     [0:0]    port_state_out_6_0_7,
  output     [0:0]    port_state_out_6_1_0,
  output     [0:0]    port_state_out_6_1_1,
  output     [0:0]    port_state_out_6_1_2,
  output     [0:0]    port_state_out_6_1_3,
  output     [0:0]    port_state_out_6_1_4,
  output     [0:0]    port_state_out_6_1_5,
  output     [0:0]    port_state_out_6_1_6,
  output     [0:0]    port_state_out_6_1_7,
  output     [0:0]    port_state_out_7_0_0,
  output     [0:0]    port_state_out_7_0_1,
  output     [0:0]    port_state_out_7_0_2,
  output     [0:0]    port_state_out_7_0_3,
  output     [0:0]    port_state_out_7_0_4,
  output     [0:0]    port_state_out_7_0_5,
  output     [0:0]    port_state_out_7_0_6,
  output     [0:0]    port_state_out_7_0_7,
  output     [0:0]    port_state_out_7_1_0,
  output     [0:0]    port_state_out_7_1_1,
  output     [0:0]    port_state_out_7_1_2,
  output     [0:0]    port_state_out_7_1_3,
  output     [0:0]    port_state_out_7_1_4,
  output     [0:0]    port_state_out_7_1_5,
  output     [0:0]    port_state_out_7_1_6,
  output     [0:0]    port_state_out_7_1_7,
  output     [0:0]    port_state_out_8_0_0,
  output     [0:0]    port_state_out_8_0_1,
  output     [0:0]    port_state_out_8_0_2,
  output     [0:0]    port_state_out_8_0_3,
  output     [0:0]    port_state_out_8_0_4,
  output     [0:0]    port_state_out_8_0_5,
  output     [0:0]    port_state_out_8_0_6,
  output     [0:0]    port_state_out_8_0_7,
  output     [0:0]    port_state_out_8_1_0,
  output     [0:0]    port_state_out_8_1_1,
  output     [0:0]    port_state_out_8_1_2,
  output     [0:0]    port_state_out_8_1_3,
  output     [0:0]    port_state_out_8_1_4,
  output     [0:0]    port_state_out_8_1_5,
  output     [0:0]    port_state_out_8_1_6,
  output     [0:0]    port_state_out_8_1_7,
  output     [0:0]    port_state_out_9_0_0,
  output     [0:0]    port_state_out_9_0_1,
  output     [0:0]    port_state_out_9_0_2,
  output     [0:0]    port_state_out_9_0_3,
  output     [0:0]    port_state_out_9_0_4,
  output     [0:0]    port_state_out_9_0_5,
  output     [0:0]    port_state_out_9_0_6,
  output     [0:0]    port_state_out_9_0_7,
  output     [0:0]    port_state_out_9_1_0,
  output     [0:0]    port_state_out_9_1_1,
  output     [0:0]    port_state_out_9_1_2,
  output     [0:0]    port_state_out_9_1_3,
  output     [0:0]    port_state_out_9_1_4,
  output     [0:0]    port_state_out_9_1_5,
  output     [0:0]    port_state_out_9_1_6,
  output     [0:0]    port_state_out_9_1_7,
  output     [0:0]    port_state_out_10_0_0,
  output     [0:0]    port_state_out_10_0_1,
  output     [0:0]    port_state_out_10_0_2,
  output     [0:0]    port_state_out_10_0_3,
  output     [0:0]    port_state_out_10_0_4,
  output     [0:0]    port_state_out_10_0_5,
  output     [0:0]    port_state_out_10_0_6,
  output     [0:0]    port_state_out_10_0_7,
  output     [0:0]    port_state_out_10_1_0,
  output     [0:0]    port_state_out_10_1_1,
  output     [0:0]    port_state_out_10_1_2,
  output     [0:0]    port_state_out_10_1_3,
  output     [0:0]    port_state_out_10_1_4,
  output     [0:0]    port_state_out_10_1_5,
  output     [0:0]    port_state_out_10_1_6,
  output     [0:0]    port_state_out_10_1_7,
  output     [0:0]    port_state_out_11_0_0,
  output     [0:0]    port_state_out_11_0_1,
  output     [0:0]    port_state_out_11_0_2,
  output     [0:0]    port_state_out_11_0_3,
  output     [0:0]    port_state_out_11_0_4,
  output     [0:0]    port_state_out_11_0_5,
  output     [0:0]    port_state_out_11_0_6,
  output     [0:0]    port_state_out_11_0_7,
  output     [0:0]    port_state_out_11_1_0,
  output     [0:0]    port_state_out_11_1_1,
  output     [0:0]    port_state_out_11_1_2,
  output     [0:0]    port_state_out_11_1_3,
  output     [0:0]    port_state_out_11_1_4,
  output     [0:0]    port_state_out_11_1_5,
  output     [0:0]    port_state_out_11_1_6,
  output     [0:0]    port_state_out_11_1_7,
  output     [0:0]    port_state_out_12_0_0,
  output     [0:0]    port_state_out_12_0_1,
  output     [0:0]    port_state_out_12_0_2,
  output     [0:0]    port_state_out_12_0_3,
  output     [0:0]    port_state_out_12_0_4,
  output     [0:0]    port_state_out_12_0_5,
  output     [0:0]    port_state_out_12_0_6,
  output     [0:0]    port_state_out_12_0_7,
  output     [0:0]    port_state_out_12_1_0,
  output     [0:0]    port_state_out_12_1_1,
  output     [0:0]    port_state_out_12_1_2,
  output     [0:0]    port_state_out_12_1_3,
  output     [0:0]    port_state_out_12_1_4,
  output     [0:0]    port_state_out_12_1_5,
  output     [0:0]    port_state_out_12_1_6,
  output     [0:0]    port_state_out_12_1_7,
  output     [0:0]    port_state_out_13_0_0,
  output     [0:0]    port_state_out_13_0_1,
  output     [0:0]    port_state_out_13_0_2,
  output     [0:0]    port_state_out_13_0_3,
  output     [0:0]    port_state_out_13_0_4,
  output     [0:0]    port_state_out_13_0_5,
  output     [0:0]    port_state_out_13_0_6,
  output     [0:0]    port_state_out_13_0_7,
  output     [0:0]    port_state_out_13_1_0,
  output     [0:0]    port_state_out_13_1_1,
  output     [0:0]    port_state_out_13_1_2,
  output     [0:0]    port_state_out_13_1_3,
  output     [0:0]    port_state_out_13_1_4,
  output     [0:0]    port_state_out_13_1_5,
  output     [0:0]    port_state_out_13_1_6,
  output     [0:0]    port_state_out_13_1_7,
  output     [0:0]    port_state_out_14_0_0,
  output     [0:0]    port_state_out_14_0_1,
  output     [0:0]    port_state_out_14_0_2,
  output     [0:0]    port_state_out_14_0_3,
  output     [0:0]    port_state_out_14_0_4,
  output     [0:0]    port_state_out_14_0_5,
  output     [0:0]    port_state_out_14_0_6,
  output     [0:0]    port_state_out_14_0_7,
  output     [0:0]    port_state_out_14_1_0,
  output     [0:0]    port_state_out_14_1_1,
  output     [0:0]    port_state_out_14_1_2,
  output     [0:0]    port_state_out_14_1_3,
  output     [0:0]    port_state_out_14_1_4,
  output     [0:0]    port_state_out_14_1_5,
  output     [0:0]    port_state_out_14_1_6,
  output     [0:0]    port_state_out_14_1_7,
  output     [0:0]    port_state_out_15_0_0,
  output     [0:0]    port_state_out_15_0_1,
  output     [0:0]    port_state_out_15_0_2,
  output     [0:0]    port_state_out_15_0_3,
  output     [0:0]    port_state_out_15_0_4,
  output     [0:0]    port_state_out_15_0_5,
  output     [0:0]    port_state_out_15_0_6,
  output     [0:0]    port_state_out_15_0_7,
  output     [0:0]    port_state_out_15_1_0,
  output     [0:0]    port_state_out_15_1_1,
  output     [0:0]    port_state_out_15_1_2,
  output     [0:0]    port_state_out_15_1_3,
  output     [0:0]    port_state_out_15_1_4,
  output     [0:0]    port_state_out_15_1_5,
  output     [0:0]    port_state_out_15_1_6,
  output     [0:0]    port_state_out_15_1_7
);


  assign port_state_out_0_0_0 = port_state_in_0_0_0;
  assign port_state_out_0_0_1 = port_state_in_0_0_1;
  assign port_state_out_0_0_2 = port_state_in_0_0_2;
  assign port_state_out_0_0_3 = port_state_in_0_0_3;
  assign port_state_out_0_0_4 = port_state_in_0_0_4;
  assign port_state_out_0_0_5 = port_state_in_0_0_5;
  assign port_state_out_0_0_6 = port_state_in_0_0_6;
  assign port_state_out_0_0_7 = port_state_in_0_0_7;
  assign port_state_out_0_1_0 = port_state_in_0_1_0;
  assign port_state_out_0_1_1 = port_state_in_0_1_1;
  assign port_state_out_0_1_2 = port_state_in_0_1_2;
  assign port_state_out_0_1_3 = port_state_in_0_1_3;
  assign port_state_out_0_1_4 = port_state_in_0_1_4;
  assign port_state_out_0_1_5 = port_state_in_0_1_5;
  assign port_state_out_0_1_6 = port_state_in_0_1_6;
  assign port_state_out_0_1_7 = port_state_in_0_1_7;
  assign port_state_out_1_0_0 = port_state_in_5_0_0;
  assign port_state_out_1_0_1 = port_state_in_5_0_1;
  assign port_state_out_1_0_2 = port_state_in_5_0_2;
  assign port_state_out_1_0_3 = port_state_in_5_0_3;
  assign port_state_out_1_0_4 = port_state_in_5_0_4;
  assign port_state_out_1_0_5 = port_state_in_5_0_5;
  assign port_state_out_1_0_6 = port_state_in_5_0_6;
  assign port_state_out_1_0_7 = port_state_in_5_0_7;
  assign port_state_out_1_1_0 = port_state_in_5_1_0;
  assign port_state_out_1_1_1 = port_state_in_5_1_1;
  assign port_state_out_1_1_2 = port_state_in_5_1_2;
  assign port_state_out_1_1_3 = port_state_in_5_1_3;
  assign port_state_out_1_1_4 = port_state_in_5_1_4;
  assign port_state_out_1_1_5 = port_state_in_5_1_5;
  assign port_state_out_1_1_6 = port_state_in_5_1_6;
  assign port_state_out_1_1_7 = port_state_in_5_1_7;
  assign port_state_out_2_0_0 = port_state_in_10_0_0;
  assign port_state_out_2_0_1 = port_state_in_10_0_1;
  assign port_state_out_2_0_2 = port_state_in_10_0_2;
  assign port_state_out_2_0_3 = port_state_in_10_0_3;
  assign port_state_out_2_0_4 = port_state_in_10_0_4;
  assign port_state_out_2_0_5 = port_state_in_10_0_5;
  assign port_state_out_2_0_6 = port_state_in_10_0_6;
  assign port_state_out_2_0_7 = port_state_in_10_0_7;
  assign port_state_out_2_1_0 = port_state_in_10_1_0;
  assign port_state_out_2_1_1 = port_state_in_10_1_1;
  assign port_state_out_2_1_2 = port_state_in_10_1_2;
  assign port_state_out_2_1_3 = port_state_in_10_1_3;
  assign port_state_out_2_1_4 = port_state_in_10_1_4;
  assign port_state_out_2_1_5 = port_state_in_10_1_5;
  assign port_state_out_2_1_6 = port_state_in_10_1_6;
  assign port_state_out_2_1_7 = port_state_in_10_1_7;
  assign port_state_out_3_0_0 = port_state_in_15_0_0;
  assign port_state_out_3_0_1 = port_state_in_15_0_1;
  assign port_state_out_3_0_2 = port_state_in_15_0_2;
  assign port_state_out_3_0_3 = port_state_in_15_0_3;
  assign port_state_out_3_0_4 = port_state_in_15_0_4;
  assign port_state_out_3_0_5 = port_state_in_15_0_5;
  assign port_state_out_3_0_6 = port_state_in_15_0_6;
  assign port_state_out_3_0_7 = port_state_in_15_0_7;
  assign port_state_out_3_1_0 = port_state_in_15_1_0;
  assign port_state_out_3_1_1 = port_state_in_15_1_1;
  assign port_state_out_3_1_2 = port_state_in_15_1_2;
  assign port_state_out_3_1_3 = port_state_in_15_1_3;
  assign port_state_out_3_1_4 = port_state_in_15_1_4;
  assign port_state_out_3_1_5 = port_state_in_15_1_5;
  assign port_state_out_3_1_6 = port_state_in_15_1_6;
  assign port_state_out_3_1_7 = port_state_in_15_1_7;
  assign port_state_out_4_0_0 = port_state_in_4_0_0;
  assign port_state_out_4_0_1 = port_state_in_4_0_1;
  assign port_state_out_4_0_2 = port_state_in_4_0_2;
  assign port_state_out_4_0_3 = port_state_in_4_0_3;
  assign port_state_out_4_0_4 = port_state_in_4_0_4;
  assign port_state_out_4_0_5 = port_state_in_4_0_5;
  assign port_state_out_4_0_6 = port_state_in_4_0_6;
  assign port_state_out_4_0_7 = port_state_in_4_0_7;
  assign port_state_out_4_1_0 = port_state_in_4_1_0;
  assign port_state_out_4_1_1 = port_state_in_4_1_1;
  assign port_state_out_4_1_2 = port_state_in_4_1_2;
  assign port_state_out_4_1_3 = port_state_in_4_1_3;
  assign port_state_out_4_1_4 = port_state_in_4_1_4;
  assign port_state_out_4_1_5 = port_state_in_4_1_5;
  assign port_state_out_4_1_6 = port_state_in_4_1_6;
  assign port_state_out_4_1_7 = port_state_in_4_1_7;
  assign port_state_out_5_0_0 = port_state_in_9_0_0;
  assign port_state_out_5_0_1 = port_state_in_9_0_1;
  assign port_state_out_5_0_2 = port_state_in_9_0_2;
  assign port_state_out_5_0_3 = port_state_in_9_0_3;
  assign port_state_out_5_0_4 = port_state_in_9_0_4;
  assign port_state_out_5_0_5 = port_state_in_9_0_5;
  assign port_state_out_5_0_6 = port_state_in_9_0_6;
  assign port_state_out_5_0_7 = port_state_in_9_0_7;
  assign port_state_out_5_1_0 = port_state_in_9_1_0;
  assign port_state_out_5_1_1 = port_state_in_9_1_1;
  assign port_state_out_5_1_2 = port_state_in_9_1_2;
  assign port_state_out_5_1_3 = port_state_in_9_1_3;
  assign port_state_out_5_1_4 = port_state_in_9_1_4;
  assign port_state_out_5_1_5 = port_state_in_9_1_5;
  assign port_state_out_5_1_6 = port_state_in_9_1_6;
  assign port_state_out_5_1_7 = port_state_in_9_1_7;
  assign port_state_out_6_0_0 = port_state_in_14_0_0;
  assign port_state_out_6_0_1 = port_state_in_14_0_1;
  assign port_state_out_6_0_2 = port_state_in_14_0_2;
  assign port_state_out_6_0_3 = port_state_in_14_0_3;
  assign port_state_out_6_0_4 = port_state_in_14_0_4;
  assign port_state_out_6_0_5 = port_state_in_14_0_5;
  assign port_state_out_6_0_6 = port_state_in_14_0_6;
  assign port_state_out_6_0_7 = port_state_in_14_0_7;
  assign port_state_out_6_1_0 = port_state_in_14_1_0;
  assign port_state_out_6_1_1 = port_state_in_14_1_1;
  assign port_state_out_6_1_2 = port_state_in_14_1_2;
  assign port_state_out_6_1_3 = port_state_in_14_1_3;
  assign port_state_out_6_1_4 = port_state_in_14_1_4;
  assign port_state_out_6_1_5 = port_state_in_14_1_5;
  assign port_state_out_6_1_6 = port_state_in_14_1_6;
  assign port_state_out_6_1_7 = port_state_in_14_1_7;
  assign port_state_out_7_0_0 = port_state_in_3_0_0;
  assign port_state_out_7_0_1 = port_state_in_3_0_1;
  assign port_state_out_7_0_2 = port_state_in_3_0_2;
  assign port_state_out_7_0_3 = port_state_in_3_0_3;
  assign port_state_out_7_0_4 = port_state_in_3_0_4;
  assign port_state_out_7_0_5 = port_state_in_3_0_5;
  assign port_state_out_7_0_6 = port_state_in_3_0_6;
  assign port_state_out_7_0_7 = port_state_in_3_0_7;
  assign port_state_out_7_1_0 = port_state_in_3_1_0;
  assign port_state_out_7_1_1 = port_state_in_3_1_1;
  assign port_state_out_7_1_2 = port_state_in_3_1_2;
  assign port_state_out_7_1_3 = port_state_in_3_1_3;
  assign port_state_out_7_1_4 = port_state_in_3_1_4;
  assign port_state_out_7_1_5 = port_state_in_3_1_5;
  assign port_state_out_7_1_6 = port_state_in_3_1_6;
  assign port_state_out_7_1_7 = port_state_in_3_1_7;
  assign port_state_out_8_0_0 = port_state_in_8_0_0;
  assign port_state_out_8_0_1 = port_state_in_8_0_1;
  assign port_state_out_8_0_2 = port_state_in_8_0_2;
  assign port_state_out_8_0_3 = port_state_in_8_0_3;
  assign port_state_out_8_0_4 = port_state_in_8_0_4;
  assign port_state_out_8_0_5 = port_state_in_8_0_5;
  assign port_state_out_8_0_6 = port_state_in_8_0_6;
  assign port_state_out_8_0_7 = port_state_in_8_0_7;
  assign port_state_out_8_1_0 = port_state_in_8_1_0;
  assign port_state_out_8_1_1 = port_state_in_8_1_1;
  assign port_state_out_8_1_2 = port_state_in_8_1_2;
  assign port_state_out_8_1_3 = port_state_in_8_1_3;
  assign port_state_out_8_1_4 = port_state_in_8_1_4;
  assign port_state_out_8_1_5 = port_state_in_8_1_5;
  assign port_state_out_8_1_6 = port_state_in_8_1_6;
  assign port_state_out_8_1_7 = port_state_in_8_1_7;
  assign port_state_out_9_0_0 = port_state_in_13_0_0;
  assign port_state_out_9_0_1 = port_state_in_13_0_1;
  assign port_state_out_9_0_2 = port_state_in_13_0_2;
  assign port_state_out_9_0_3 = port_state_in_13_0_3;
  assign port_state_out_9_0_4 = port_state_in_13_0_4;
  assign port_state_out_9_0_5 = port_state_in_13_0_5;
  assign port_state_out_9_0_6 = port_state_in_13_0_6;
  assign port_state_out_9_0_7 = port_state_in_13_0_7;
  assign port_state_out_9_1_0 = port_state_in_13_1_0;
  assign port_state_out_9_1_1 = port_state_in_13_1_1;
  assign port_state_out_9_1_2 = port_state_in_13_1_2;
  assign port_state_out_9_1_3 = port_state_in_13_1_3;
  assign port_state_out_9_1_4 = port_state_in_13_1_4;
  assign port_state_out_9_1_5 = port_state_in_13_1_5;
  assign port_state_out_9_1_6 = port_state_in_13_1_6;
  assign port_state_out_9_1_7 = port_state_in_13_1_7;
  assign port_state_out_10_0_0 = port_state_in_2_0_0;
  assign port_state_out_10_0_1 = port_state_in_2_0_1;
  assign port_state_out_10_0_2 = port_state_in_2_0_2;
  assign port_state_out_10_0_3 = port_state_in_2_0_3;
  assign port_state_out_10_0_4 = port_state_in_2_0_4;
  assign port_state_out_10_0_5 = port_state_in_2_0_5;
  assign port_state_out_10_0_6 = port_state_in_2_0_6;
  assign port_state_out_10_0_7 = port_state_in_2_0_7;
  assign port_state_out_10_1_0 = port_state_in_2_1_0;
  assign port_state_out_10_1_1 = port_state_in_2_1_1;
  assign port_state_out_10_1_2 = port_state_in_2_1_2;
  assign port_state_out_10_1_3 = port_state_in_2_1_3;
  assign port_state_out_10_1_4 = port_state_in_2_1_4;
  assign port_state_out_10_1_5 = port_state_in_2_1_5;
  assign port_state_out_10_1_6 = port_state_in_2_1_6;
  assign port_state_out_10_1_7 = port_state_in_2_1_7;
  assign port_state_out_11_0_0 = port_state_in_7_0_0;
  assign port_state_out_11_0_1 = port_state_in_7_0_1;
  assign port_state_out_11_0_2 = port_state_in_7_0_2;
  assign port_state_out_11_0_3 = port_state_in_7_0_3;
  assign port_state_out_11_0_4 = port_state_in_7_0_4;
  assign port_state_out_11_0_5 = port_state_in_7_0_5;
  assign port_state_out_11_0_6 = port_state_in_7_0_6;
  assign port_state_out_11_0_7 = port_state_in_7_0_7;
  assign port_state_out_11_1_0 = port_state_in_7_1_0;
  assign port_state_out_11_1_1 = port_state_in_7_1_1;
  assign port_state_out_11_1_2 = port_state_in_7_1_2;
  assign port_state_out_11_1_3 = port_state_in_7_1_3;
  assign port_state_out_11_1_4 = port_state_in_7_1_4;
  assign port_state_out_11_1_5 = port_state_in_7_1_5;
  assign port_state_out_11_1_6 = port_state_in_7_1_6;
  assign port_state_out_11_1_7 = port_state_in_7_1_7;
  assign port_state_out_12_0_0 = port_state_in_12_0_0;
  assign port_state_out_12_0_1 = port_state_in_12_0_1;
  assign port_state_out_12_0_2 = port_state_in_12_0_2;
  assign port_state_out_12_0_3 = port_state_in_12_0_3;
  assign port_state_out_12_0_4 = port_state_in_12_0_4;
  assign port_state_out_12_0_5 = port_state_in_12_0_5;
  assign port_state_out_12_0_6 = port_state_in_12_0_6;
  assign port_state_out_12_0_7 = port_state_in_12_0_7;
  assign port_state_out_12_1_0 = port_state_in_12_1_0;
  assign port_state_out_12_1_1 = port_state_in_12_1_1;
  assign port_state_out_12_1_2 = port_state_in_12_1_2;
  assign port_state_out_12_1_3 = port_state_in_12_1_3;
  assign port_state_out_12_1_4 = port_state_in_12_1_4;
  assign port_state_out_12_1_5 = port_state_in_12_1_5;
  assign port_state_out_12_1_6 = port_state_in_12_1_6;
  assign port_state_out_12_1_7 = port_state_in_12_1_7;
  assign port_state_out_13_0_0 = port_state_in_1_0_0;
  assign port_state_out_13_0_1 = port_state_in_1_0_1;
  assign port_state_out_13_0_2 = port_state_in_1_0_2;
  assign port_state_out_13_0_3 = port_state_in_1_0_3;
  assign port_state_out_13_0_4 = port_state_in_1_0_4;
  assign port_state_out_13_0_5 = port_state_in_1_0_5;
  assign port_state_out_13_0_6 = port_state_in_1_0_6;
  assign port_state_out_13_0_7 = port_state_in_1_0_7;
  assign port_state_out_13_1_0 = port_state_in_1_1_0;
  assign port_state_out_13_1_1 = port_state_in_1_1_1;
  assign port_state_out_13_1_2 = port_state_in_1_1_2;
  assign port_state_out_13_1_3 = port_state_in_1_1_3;
  assign port_state_out_13_1_4 = port_state_in_1_1_4;
  assign port_state_out_13_1_5 = port_state_in_1_1_5;
  assign port_state_out_13_1_6 = port_state_in_1_1_6;
  assign port_state_out_13_1_7 = port_state_in_1_1_7;
  assign port_state_out_14_0_0 = port_state_in_6_0_0;
  assign port_state_out_14_0_1 = port_state_in_6_0_1;
  assign port_state_out_14_0_2 = port_state_in_6_0_2;
  assign port_state_out_14_0_3 = port_state_in_6_0_3;
  assign port_state_out_14_0_4 = port_state_in_6_0_4;
  assign port_state_out_14_0_5 = port_state_in_6_0_5;
  assign port_state_out_14_0_6 = port_state_in_6_0_6;
  assign port_state_out_14_0_7 = port_state_in_6_0_7;
  assign port_state_out_14_1_0 = port_state_in_6_1_0;
  assign port_state_out_14_1_1 = port_state_in_6_1_1;
  assign port_state_out_14_1_2 = port_state_in_6_1_2;
  assign port_state_out_14_1_3 = port_state_in_6_1_3;
  assign port_state_out_14_1_4 = port_state_in_6_1_4;
  assign port_state_out_14_1_5 = port_state_in_6_1_5;
  assign port_state_out_14_1_6 = port_state_in_6_1_6;
  assign port_state_out_14_1_7 = port_state_in_6_1_7;
  assign port_state_out_15_0_0 = port_state_in_11_0_0;
  assign port_state_out_15_0_1 = port_state_in_11_0_1;
  assign port_state_out_15_0_2 = port_state_in_11_0_2;
  assign port_state_out_15_0_3 = port_state_in_11_0_3;
  assign port_state_out_15_0_4 = port_state_in_11_0_4;
  assign port_state_out_15_0_5 = port_state_in_11_0_5;
  assign port_state_out_15_0_6 = port_state_in_11_0_6;
  assign port_state_out_15_0_7 = port_state_in_11_0_7;
  assign port_state_out_15_1_0 = port_state_in_11_1_0;
  assign port_state_out_15_1_1 = port_state_in_11_1_1;
  assign port_state_out_15_1_2 = port_state_in_11_1_2;
  assign port_state_out_15_1_3 = port_state_in_11_1_3;
  assign port_state_out_15_1_4 = port_state_in_11_1_4;
  assign port_state_out_15_1_5 = port_state_in_11_1_5;
  assign port_state_out_15_1_6 = port_state_in_11_1_6;
  assign port_state_out_15_1_7 = port_state_in_11_1_7;

endmodule

//Sbox_AES_Canright_CMS_2shares replaced by Sbox_AES_Canright_CMS_2shares

//Sbox_AES_Canright_CMS_2shares replaced by Sbox_AES_Canright_CMS_2shares

//Sbox_AES_Canright_CMS_2shares replaced by Sbox_AES_Canright_CMS_2shares

//Sbox_AES_Canright_CMS_2shares replaced by Sbox_AES_Canright_CMS_2shares

//Sbox_AES_Canright_CMS_2shares replaced by Sbox_AES_Canright_CMS_2shares

//Sbox_AES_Canright_CMS_2shares replaced by Sbox_AES_Canright_CMS_2shares

//Sbox_AES_Canright_CMS_2shares replaced by Sbox_AES_Canright_CMS_2shares

//Sbox_AES_Canright_CMS_2shares replaced by Sbox_AES_Canright_CMS_2shares

//Sbox_AES_Canright_CMS_2shares replaced by Sbox_AES_Canright_CMS_2shares

//Sbox_AES_Canright_CMS_2shares replaced by Sbox_AES_Canright_CMS_2shares

//Sbox_AES_Canright_CMS_2shares replaced by Sbox_AES_Canright_CMS_2shares

//Sbox_AES_Canright_CMS_2shares replaced by Sbox_AES_Canright_CMS_2shares

//Sbox_AES_Canright_CMS_2shares replaced by Sbox_AES_Canright_CMS_2shares

//Sbox_AES_Canright_CMS_2shares replaced by Sbox_AES_Canright_CMS_2shares

//Sbox_AES_Canright_CMS_2shares replaced by Sbox_AES_Canright_CMS_2shares

module Sbox_AES_Canright_CMS_2shares (
  input      [0:0]    port_i_0_0,
  input      [0:0]    port_i_0_1,
  input      [0:0]    port_i_0_2,
  input      [0:0]    port_i_0_3,
  input      [0:0]    port_i_0_4,
  input      [0:0]    port_i_0_5,
  input      [0:0]    port_i_0_6,
  input      [0:0]    port_i_0_7,
  input      [0:0]    port_i_1_0,
  input      [0:0]    port_i_1_1,
  input      [0:0]    port_i_1_2,
  input      [0:0]    port_i_1_3,
  input      [0:0]    port_i_1_4,
  input      [0:0]    port_i_1_5,
  input      [0:0]    port_i_1_6,
  input      [0:0]    port_i_1_7,
  input               port_r_0,
  input               port_r_1,
  input               port_r_2,
  input               port_r_3,
  input               port_r_4,
  input               port_r_5,
  input               port_r_6,
  input               port_r_7,
  input               port_r_8,
  input               port_r_9,
  input               port_r_10,
  input               port_r_11,
  input               port_r_12,
  input               port_r_13,
  input               port_r_14,
  input               port_r_15,
  input               port_r_16,
  input               port_r_17,
  input               port_r_18,
  input               port_r_19,
  input               port_r_20,
  input               port_r_21,
  input               port_r_22,
  input               port_r_23,
  input               port_r_24,
  input               port_r_25,
  input               port_r_26,
  input               port_r_27,
  input               port_r_28,
  input               port_r_29,
  input               port_r_30,
  input               port_r_31,
  input               port_r_32,
  input               port_r_33,
  input               port_r_34,
  input               port_r_35,
  input               port_r_36,
  input               port_r_37,
  input               port_r_38,
  input               port_r_39,
  input               port_r_40,
  input               port_r_41,
  input               port_r_42,
  input               port_r_43,
  input               port_r_44,
  input               port_r_45,
  input               port_r_46,
  input               port_r_47,
  input               port_r_48,
  input               port_r_49,
  input               port_r_50,
  input               port_r_51,
  input               port_r_52,
  input               port_r_53,
  output     [0:0]    port_o_0_0,
  output     [0:0]    port_o_0_1,
  output     [0:0]    port_o_0_2,
  output     [0:0]    port_o_0_3,
  output     [0:0]    port_o_0_4,
  output     [0:0]    port_o_0_5,
  output     [0:0]    port_o_0_6,
  output     [0:0]    port_o_0_7,
  output     [0:0]    port_o_1_0,
  output     [0:0]    port_o_1_1,
  output     [0:0]    port_o_1_2,
  output     [0:0]    port_o_1_3,
  output     [0:0]    port_o_1_4,
  output     [0:0]    port_o_1_5,
  output     [0:0]    port_o_1_6,
  output     [0:0]    port_o_1_7,
  input               clk,
  input               reset
);

  wire       [0:0]    stage6_port_i_0_0;
  wire       [0:0]    stage6_port_i_0_1;
  wire       [0:0]    stage6_port_i_0_2;
  wire       [0:0]    stage6_port_i_0_3;
  wire       [0:0]    stage6_port_i_0_4;
  wire       [0:0]    stage6_port_i_0_5;
  wire       [0:0]    stage6_port_i_0_6;
  wire       [0:0]    stage6_port_i_0_7;
  wire       [0:0]    stage6_port_i_1_0;
  wire       [0:0]    stage6_port_i_1_1;
  wire       [0:0]    stage6_port_i_1_2;
  wire       [0:0]    stage6_port_i_1_3;
  wire       [0:0]    stage6_port_i_1_4;
  wire       [0:0]    stage6_port_i_1_5;
  wire       [0:0]    stage6_port_i_1_6;
  wire       [0:0]    stage6_port_i_1_7;
  wire       [0:0]    stage1_port_o_0_0;
  wire       [0:0]    stage1_port_o_0_1;
  wire       [0:0]    stage1_port_o_0_2;
  wire       [0:0]    stage1_port_o_0_3;
  wire       [0:0]    stage1_port_o_0_4;
  wire       [0:0]    stage1_port_o_0_5;
  wire       [0:0]    stage1_port_o_0_6;
  wire       [0:0]    stage1_port_o_0_7;
  wire       [0:0]    stage1_port_o_1_0;
  wire       [0:0]    stage1_port_o_1_1;
  wire       [0:0]    stage1_port_o_1_2;
  wire       [0:0]    stage1_port_o_1_3;
  wire       [0:0]    stage1_port_o_1_4;
  wire       [0:0]    stage1_port_o_1_5;
  wire       [0:0]    stage1_port_o_1_6;
  wire       [0:0]    stage1_port_o_1_7;
  wire       [0:0]    stage2_port_y_0_0;
  wire       [0:0]    stage2_port_y_0_1;
  wire       [0:0]    stage2_port_y_0_2;
  wire       [0:0]    stage2_port_y_0_3;
  wire       [0:0]    stage2_port_y_1_0;
  wire       [0:0]    stage2_port_y_1_1;
  wire       [0:0]    stage2_port_y_1_2;
  wire       [0:0]    stage2_port_y_1_3;
  wire       [0:0]    stage2_port_y_2_0;
  wire       [0:0]    stage2_port_y_2_1;
  wire       [0:0]    stage2_port_y_2_2;
  wire       [0:0]    stage2_port_y_2_3;
  wire       [0:0]    stage2_port_y_3_0;
  wire       [0:0]    stage2_port_y_3_1;
  wire       [0:0]    stage2_port_y_3_2;
  wire       [0:0]    stage2_port_y_3_3;
  wire       [0:0]    stage3_port_y_0_0;
  wire       [0:0]    stage3_port_y_0_1;
  wire       [0:0]    stage3_port_y_1_0;
  wire       [0:0]    stage3_port_y_1_1;
  wire       [0:0]    stage3_port_y_2_0;
  wire       [0:0]    stage3_port_y_2_1;
  wire       [0:0]    stage3_port_y_3_0;
  wire       [0:0]    stage3_port_y_3_1;
  wire       [0:0]    stage4_port_y_0_0;
  wire       [0:0]    stage4_port_y_0_1;
  wire       [0:0]    stage4_port_y_0_2;
  wire       [0:0]    stage4_port_y_0_3;
  wire       [0:0]    stage4_port_y_1_0;
  wire       [0:0]    stage4_port_y_1_1;
  wire       [0:0]    stage4_port_y_1_2;
  wire       [0:0]    stage4_port_y_1_3;
  wire       [0:0]    stage4_port_y_2_0;
  wire       [0:0]    stage4_port_y_2_1;
  wire       [0:0]    stage4_port_y_2_2;
  wire       [0:0]    stage4_port_y_2_3;
  wire       [0:0]    stage4_port_y_3_0;
  wire       [0:0]    stage4_port_y_3_1;
  wire       [0:0]    stage4_port_y_3_2;
  wire       [0:0]    stage4_port_y_3_3;
  wire       [0:0]    stage5_port_y_0_0;
  wire       [0:0]    stage5_port_y_0_1;
  wire       [0:0]    stage5_port_y_0_2;
  wire       [0:0]    stage5_port_y_0_3;
  wire       [0:0]    stage5_port_y_0_4;
  wire       [0:0]    stage5_port_y_0_5;
  wire       [0:0]    stage5_port_y_0_6;
  wire       [0:0]    stage5_port_y_0_7;
  wire       [0:0]    stage5_port_y_1_0;
  wire       [0:0]    stage5_port_y_1_1;
  wire       [0:0]    stage5_port_y_1_2;
  wire       [0:0]    stage5_port_y_1_3;
  wire       [0:0]    stage5_port_y_1_4;
  wire       [0:0]    stage5_port_y_1_5;
  wire       [0:0]    stage5_port_y_1_6;
  wire       [0:0]    stage5_port_y_1_7;
  wire       [0:0]    stage5_port_y_2_0;
  wire       [0:0]    stage5_port_y_2_1;
  wire       [0:0]    stage5_port_y_2_2;
  wire       [0:0]    stage5_port_y_2_3;
  wire       [0:0]    stage5_port_y_2_4;
  wire       [0:0]    stage5_port_y_2_5;
  wire       [0:0]    stage5_port_y_2_6;
  wire       [0:0]    stage5_port_y_2_7;
  wire       [0:0]    stage5_port_y_3_0;
  wire       [0:0]    stage5_port_y_3_1;
  wire       [0:0]    stage5_port_y_3_2;
  wire       [0:0]    stage5_port_y_3_3;
  wire       [0:0]    stage5_port_y_3_4;
  wire       [0:0]    stage5_port_y_3_5;
  wire       [0:0]    stage5_port_y_3_6;
  wire       [0:0]    stage5_port_y_3_7;
  wire       [0:0]    stage6_port_o_0_0;
  wire       [0:0]    stage6_port_o_0_1;
  wire       [0:0]    stage6_port_o_0_2;
  wire       [0:0]    stage6_port_o_0_3;
  wire       [0:0]    stage6_port_o_0_4;
  wire       [0:0]    stage6_port_o_0_5;
  wire       [0:0]    stage6_port_o_0_6;
  wire       [0:0]    stage6_port_o_0_7;
  wire       [0:0]    stage6_port_o_1_0;
  wire       [0:0]    stage6_port_o_1_1;
  wire       [0:0]    stage6_port_o_1_2;
  wire       [0:0]    stage6_port_o_1_3;
  wire       [0:0]    stage6_port_o_1_4;
  wire       [0:0]    stage6_port_o_1_5;
  wire       [0:0]    stage6_port_o_1_6;
  wire       [0:0]    stage6_port_o_1_7;
  wire       [0:0]    ax_0_0;
  wire       [0:0]    ax_0_1;
  wire       [0:0]    ax_0_2;
  wire       [0:0]    ax_0_3;
  wire       [0:0]    ax_1_0;
  wire       [0:0]    ax_1_1;
  wire       [0:0]    ax_1_2;
  wire       [0:0]    ax_1_3;
  wire       [0:0]    bx_0_0;
  wire       [0:0]    bx_0_1;
  wire       [0:0]    bx_0_2;
  wire       [0:0]    bx_0_3;
  wire       [0:0]    bx_1_0;
  wire       [0:0]    bx_1_1;
  wire       [0:0]    bx_1_2;
  wire       [0:0]    bx_1_3;
  wire       [0:0]    ax1_0_0;
  wire       [0:0]    ax1_0_1;
  wire       [0:0]    ax1_1_0;
  wire       [0:0]    ax1_1_1;
  wire       [0:0]    bx1_0_0;
  wire       [0:0]    bx1_0_1;
  wire       [0:0]    bx1_1_0;
  wire       [0:0]    bx1_1_1;
  reg        [0:0]    ax4_0_0;
  reg        [0:0]    ax4_0_1;
  reg        [0:0]    ax4_1_0;
  reg        [0:0]    ax4_1_1;
  reg        [0:0]    bx4_0_0;
  reg        [0:0]    bx4_0_1;
  reg        [0:0]    bx4_1_0;
  reg        [0:0]    bx4_1_1;
  wire       [0:0]    cx4_0_0;
  wire       [0:0]    cx4_0_1;
  wire       [0:0]    cx4_1_0;
  wire       [0:0]    cx4_1_1;
  reg        [0:0]    ax_reg1_0_0;
  reg        [0:0]    ax_reg1_0_1;
  reg        [0:0]    ax_reg1_0_2;
  reg        [0:0]    ax_reg1_0_3;
  reg        [0:0]    ax_reg1_1_0;
  reg        [0:0]    ax_reg1_1_1;
  reg        [0:0]    ax_reg1_1_2;
  reg        [0:0]    ax_reg1_1_3;
  reg        [0:0]    ax_reg2_0_0;
  reg        [0:0]    ax_reg2_0_1;
  reg        [0:0]    ax_reg2_0_2;
  reg        [0:0]    ax_reg2_0_3;
  reg        [0:0]    ax_reg2_1_0;
  reg        [0:0]    ax_reg2_1_1;
  reg        [0:0]    ax_reg2_1_2;
  reg        [0:0]    ax_reg2_1_3;
  reg        [0:0]    ax_reg3_0_0;
  reg        [0:0]    ax_reg3_0_1;
  reg        [0:0]    ax_reg3_0_2;
  reg        [0:0]    ax_reg3_0_3;
  reg        [0:0]    ax_reg3_1_0;
  reg        [0:0]    ax_reg3_1_1;
  reg        [0:0]    ax_reg3_1_2;
  reg        [0:0]    ax_reg3_1_3;
  reg        [0:0]    bx_reg1_0_0;
  reg        [0:0]    bx_reg1_0_1;
  reg        [0:0]    bx_reg1_0_2;
  reg        [0:0]    bx_reg1_0_3;
  reg        [0:0]    bx_reg1_1_0;
  reg        [0:0]    bx_reg1_1_1;
  reg        [0:0]    bx_reg1_1_2;
  reg        [0:0]    bx_reg1_1_3;
  reg        [0:0]    bx_reg2_0_0;
  reg        [0:0]    bx_reg2_0_1;
  reg        [0:0]    bx_reg2_0_2;
  reg        [0:0]    bx_reg2_0_3;
  reg        [0:0]    bx_reg2_1_0;
  reg        [0:0]    bx_reg2_1_1;
  reg        [0:0]    bx_reg2_1_2;
  reg        [0:0]    bx_reg2_1_3;
  reg        [0:0]    bx_reg3_0_0;
  reg        [0:0]    bx_reg3_0_1;
  reg        [0:0]    bx_reg3_0_2;
  reg        [0:0]    bx_reg3_0_3;
  reg        [0:0]    bx_reg3_1_0;
  reg        [0:0]    bx_reg3_1_1;
  reg        [0:0]    bx_reg3_1_2;
  reg        [0:0]    bx_reg3_1_3;
  wire       [0:0]    bx5_0_0;
  wire       [0:0]    bx5_0_1;
  wire       [0:0]    bx5_0_2;
  wire       [0:0]    bx5_0_3;
  wire       [0:0]    bx5_1_0;
  wire       [0:0]    bx5_1_1;
  wire       [0:0]    bx5_1_2;
  wire       [0:0]    bx5_1_3;

  CMS_stage1 stage1 (
    .port_i_0_0 (port_i_0_0       ), //i
    .port_i_0_1 (port_i_0_1       ), //i
    .port_i_0_2 (port_i_0_2       ), //i
    .port_i_0_3 (port_i_0_3       ), //i
    .port_i_0_4 (port_i_0_4       ), //i
    .port_i_0_5 (port_i_0_5       ), //i
    .port_i_0_6 (port_i_0_6       ), //i
    .port_i_0_7 (port_i_0_7       ), //i
    .port_i_1_0 (port_i_1_0       ), //i
    .port_i_1_1 (port_i_1_1       ), //i
    .port_i_1_2 (port_i_1_2       ), //i
    .port_i_1_3 (port_i_1_3       ), //i
    .port_i_1_4 (port_i_1_4       ), //i
    .port_i_1_5 (port_i_1_5       ), //i
    .port_i_1_6 (port_i_1_6       ), //i
    .port_i_1_7 (port_i_1_7       ), //i
    .port_o_0_0 (stage1_port_o_0_0), //o
    .port_o_0_1 (stage1_port_o_0_1), //o
    .port_o_0_2 (stage1_port_o_0_2), //o
    .port_o_0_3 (stage1_port_o_0_3), //o
    .port_o_0_4 (stage1_port_o_0_4), //o
    .port_o_0_5 (stage1_port_o_0_5), //o
    .port_o_0_6 (stage1_port_o_0_6), //o
    .port_o_0_7 (stage1_port_o_0_7), //o
    .port_o_1_0 (stage1_port_o_1_0), //o
    .port_o_1_1 (stage1_port_o_1_1), //o
    .port_o_1_2 (stage1_port_o_1_2), //o
    .port_o_1_3 (stage1_port_o_1_3), //o
    .port_o_1_4 (stage1_port_o_1_4), //o
    .port_o_1_5 (stage1_port_o_1_5), //o
    .port_o_1_6 (stage1_port_o_1_6), //o
    .port_o_1_7 (stage1_port_o_1_7), //o
    .clk        (clk              ), //i
    .reset      (reset            )  //i
  );
  CMS_stage2 stage2 (
    .port_a_0_0 (ax_0_0           ), //i
    .port_a_0_1 (ax_0_1           ), //i
    .port_a_0_2 (ax_0_2           ), //i
    .port_a_0_3 (ax_0_3           ), //i
    .port_a_1_0 (ax_1_0           ), //i
    .port_a_1_1 (ax_1_1           ), //i
    .port_a_1_2 (ax_1_2           ), //i
    .port_a_1_3 (ax_1_3           ), //i
    .port_b_0_0 (bx_0_0           ), //i
    .port_b_0_1 (bx_0_1           ), //i
    .port_b_0_2 (bx_0_2           ), //i
    .port_b_0_3 (bx_0_3           ), //i
    .port_b_1_0 (bx_1_0           ), //i
    .port_b_1_1 (bx_1_1           ), //i
    .port_b_1_2 (bx_1_2           ), //i
    .port_b_1_3 (bx_1_3           ), //i
    .port_r_0_0 (port_r_0         ), //i
    .port_r_0_1 (port_r_1         ), //i
    .port_r_0_2 (port_r_2         ), //i
    .port_r_0_3 (port_r_3         ), //i
    .port_r_1_0 (port_r_4         ), //i
    .port_r_1_1 (port_r_5         ), //i
    .port_r_1_2 (port_r_6         ), //i
    .port_r_1_3 (port_r_7         ), //i
    .port_r_2_0 (port_r_8         ), //i
    .port_r_2_1 (port_r_9         ), //i
    .port_r_2_2 (port_r_10        ), //i
    .port_r_2_3 (port_r_11        ), //i
    .port_y_0_0 (stage2_port_y_0_0), //o
    .port_y_0_1 (stage2_port_y_0_1), //o
    .port_y_0_2 (stage2_port_y_0_2), //o
    .port_y_0_3 (stage2_port_y_0_3), //o
    .port_y_1_0 (stage2_port_y_1_0), //o
    .port_y_1_1 (stage2_port_y_1_1), //o
    .port_y_1_2 (stage2_port_y_1_2), //o
    .port_y_1_3 (stage2_port_y_1_3), //o
    .port_y_2_0 (stage2_port_y_2_0), //o
    .port_y_2_1 (stage2_port_y_2_1), //o
    .port_y_2_2 (stage2_port_y_2_2), //o
    .port_y_2_3 (stage2_port_y_2_3), //o
    .port_y_3_0 (stage2_port_y_3_0), //o
    .port_y_3_1 (stage2_port_y_3_1), //o
    .port_y_3_2 (stage2_port_y_3_2), //o
    .port_y_3_3 (stage2_port_y_3_3), //o
    .clk        (clk              ), //i
    .reset      (reset            )  //i
  );
  CMS_stage3 stage3 (
    .port_a_0_0 (ax1_0_0          ), //i
    .port_a_0_1 (ax1_0_1          ), //i
    .port_a_1_0 (ax1_1_0          ), //i
    .port_a_1_1 (ax1_1_1          ), //i
    .port_b_0_0 (bx1_0_0          ), //i
    .port_b_0_1 (bx1_0_1          ), //i
    .port_b_1_0 (bx1_1_0          ), //i
    .port_b_1_1 (bx1_1_1          ), //i
    .port_r_0_0 (port_r_12        ), //i
    .port_r_0_1 (port_r_13        ), //i
    .port_r_1_0 (port_r_14        ), //i
    .port_r_1_1 (port_r_15        ), //i
    .port_r_2_0 (port_r_16        ), //i
    .port_r_2_1 (port_r_17        ), //i
    .port_y_0_0 (stage3_port_y_0_0), //o
    .port_y_0_1 (stage3_port_y_0_1), //o
    .port_y_1_0 (stage3_port_y_1_0), //o
    .port_y_1_1 (stage3_port_y_1_1), //o
    .port_y_2_0 (stage3_port_y_2_0), //o
    .port_y_2_1 (stage3_port_y_2_1), //o
    .port_y_3_0 (stage3_port_y_3_0), //o
    .port_y_3_1 (stage3_port_y_3_1), //o
    .clk        (clk              ), //i
    .reset      (reset            )  //i
  );
  CMS_stage4 stage4 (
    .port_a_0_0 (ax4_0_0          ), //i
    .port_a_0_1 (ax4_0_1          ), //i
    .port_a_1_0 (ax4_1_0          ), //i
    .port_a_1_1 (ax4_1_1          ), //i
    .port_b_0_0 (cx4_0_0          ), //i
    .port_b_0_1 (cx4_0_1          ), //i
    .port_b_1_0 (cx4_1_0          ), //i
    .port_b_1_1 (cx4_1_1          ), //i
    .port_c_0_0 (bx4_0_0          ), //i
    .port_c_0_1 (bx4_0_1          ), //i
    .port_c_1_0 (bx4_1_0          ), //i
    .port_c_1_1 (bx4_1_1          ), //i
    .port_r_0_0 (port_r_18        ), //i
    .port_r_0_1 (port_r_19        ), //i
    .port_r_0_2 (port_r_20        ), //i
    .port_r_0_3 (port_r_21        ), //i
    .port_r_1_0 (port_r_22        ), //i
    .port_r_1_1 (port_r_23        ), //i
    .port_r_1_2 (port_r_24        ), //i
    .port_r_1_3 (port_r_25        ), //i
    .port_r_2_0 (port_r_26        ), //i
    .port_r_2_1 (port_r_27        ), //i
    .port_r_2_2 (port_r_28        ), //i
    .port_r_2_3 (port_r_29        ), //i
    .port_y_0_0 (stage4_port_y_0_0), //o
    .port_y_0_1 (stage4_port_y_0_1), //o
    .port_y_0_2 (stage4_port_y_0_2), //o
    .port_y_0_3 (stage4_port_y_0_3), //o
    .port_y_1_0 (stage4_port_y_1_0), //o
    .port_y_1_1 (stage4_port_y_1_1), //o
    .port_y_1_2 (stage4_port_y_1_2), //o
    .port_y_1_3 (stage4_port_y_1_3), //o
    .port_y_2_0 (stage4_port_y_2_0), //o
    .port_y_2_1 (stage4_port_y_2_1), //o
    .port_y_2_2 (stage4_port_y_2_2), //o
    .port_y_2_3 (stage4_port_y_2_3), //o
    .port_y_3_0 (stage4_port_y_3_0), //o
    .port_y_3_1 (stage4_port_y_3_1), //o
    .port_y_3_2 (stage4_port_y_3_2), //o
    .port_y_3_3 (stage4_port_y_3_3), //o
    .clk        (clk              ), //i
    .reset      (reset            )  //i
  );
  CMS_stage5 stage5 (
    .port_a_0_0 (bx_reg3_0_0      ), //i
    .port_a_0_1 (bx_reg3_0_1      ), //i
    .port_a_0_2 (bx_reg3_0_2      ), //i
    .port_a_0_3 (bx_reg3_0_3      ), //i
    .port_a_1_0 (bx_reg3_1_0      ), //i
    .port_a_1_1 (bx_reg3_1_1      ), //i
    .port_a_1_2 (bx_reg3_1_2      ), //i
    .port_a_1_3 (bx_reg3_1_3      ), //i
    .port_b_0_0 (bx5_0_0          ), //i
    .port_b_0_1 (bx5_0_1          ), //i
    .port_b_0_2 (bx5_0_2          ), //i
    .port_b_0_3 (bx5_0_3          ), //i
    .port_b_1_0 (bx5_1_0          ), //i
    .port_b_1_1 (bx5_1_1          ), //i
    .port_b_1_2 (bx5_1_2          ), //i
    .port_b_1_3 (bx5_1_3          ), //i
    .port_c_0_0 (ax_reg3_0_0      ), //i
    .port_c_0_1 (ax_reg3_0_1      ), //i
    .port_c_0_2 (ax_reg3_0_2      ), //i
    .port_c_0_3 (ax_reg3_0_3      ), //i
    .port_c_1_0 (ax_reg3_1_0      ), //i
    .port_c_1_1 (ax_reg3_1_1      ), //i
    .port_c_1_2 (ax_reg3_1_2      ), //i
    .port_c_1_3 (ax_reg3_1_3      ), //i
    .port_r_0_0 (port_r_30        ), //i
    .port_r_0_1 (port_r_31        ), //i
    .port_r_0_2 (port_r_32        ), //i
    .port_r_0_3 (port_r_33        ), //i
    .port_r_0_4 (port_r_34        ), //i
    .port_r_0_5 (port_r_35        ), //i
    .port_r_0_6 (port_r_36        ), //i
    .port_r_0_7 (port_r_37        ), //i
    .port_r_1_0 (port_r_34        ), //i
    .port_r_1_1 (port_r_35        ), //i
    .port_r_1_2 (port_r_36        ), //i
    .port_r_1_3 (port_r_37        ), //i
    .port_r_1_4 (port_r_38        ), //i
    .port_r_1_5 (port_r_39        ), //i
    .port_r_1_6 (port_r_40        ), //i
    .port_r_1_7 (port_r_41        ), //i
    .port_r_2_0 (port_r_38        ), //i
    .port_r_2_1 (port_r_39        ), //i
    .port_r_2_2 (port_r_40        ), //i
    .port_r_2_3 (port_r_41        ), //i
    .port_r_2_4 (port_r_42        ), //i
    .port_r_2_5 (port_r_43        ), //i
    .port_r_2_6 (port_r_44        ), //i
    .port_r_2_7 (port_r_45        ), //i
    .port_y_0_0 (stage5_port_y_0_0), //o
    .port_y_0_1 (stage5_port_y_0_1), //o
    .port_y_0_2 (stage5_port_y_0_2), //o
    .port_y_0_3 (stage5_port_y_0_3), //o
    .port_y_0_4 (stage5_port_y_0_4), //o
    .port_y_0_5 (stage5_port_y_0_5), //o
    .port_y_0_6 (stage5_port_y_0_6), //o
    .port_y_0_7 (stage5_port_y_0_7), //o
    .port_y_1_0 (stage5_port_y_1_0), //o
    .port_y_1_1 (stage5_port_y_1_1), //o
    .port_y_1_2 (stage5_port_y_1_2), //o
    .port_y_1_3 (stage5_port_y_1_3), //o
    .port_y_1_4 (stage5_port_y_1_4), //o
    .port_y_1_5 (stage5_port_y_1_5), //o
    .port_y_1_6 (stage5_port_y_1_6), //o
    .port_y_1_7 (stage5_port_y_1_7), //o
    .port_y_2_0 (stage5_port_y_2_0), //o
    .port_y_2_1 (stage5_port_y_2_1), //o
    .port_y_2_2 (stage5_port_y_2_2), //o
    .port_y_2_3 (stage5_port_y_2_3), //o
    .port_y_2_4 (stage5_port_y_2_4), //o
    .port_y_2_5 (stage5_port_y_2_5), //o
    .port_y_2_6 (stage5_port_y_2_6), //o
    .port_y_2_7 (stage5_port_y_2_7), //o
    .port_y_3_0 (stage5_port_y_3_0), //o
    .port_y_3_1 (stage5_port_y_3_1), //o
    .port_y_3_2 (stage5_port_y_3_2), //o
    .port_y_3_3 (stage5_port_y_3_3), //o
    .port_y_3_4 (stage5_port_y_3_4), //o
    .port_y_3_5 (stage5_port_y_3_5), //o
    .port_y_3_6 (stage5_port_y_3_6), //o
    .port_y_3_7 (stage5_port_y_3_7), //o
    .clk        (clk              ), //i
    .reset      (reset            )  //i
  );
  CMS_stage6 stage6 (
    .port_i_0_0 (stage6_port_i_0_0), //i
    .port_i_0_1 (stage6_port_i_0_1), //i
    .port_i_0_2 (stage6_port_i_0_2), //i
    .port_i_0_3 (stage6_port_i_0_3), //i
    .port_i_0_4 (stage6_port_i_0_4), //i
    .port_i_0_5 (stage6_port_i_0_5), //i
    .port_i_0_6 (stage6_port_i_0_6), //i
    .port_i_0_7 (stage6_port_i_0_7), //i
    .port_i_1_0 (stage6_port_i_1_0), //i
    .port_i_1_1 (stage6_port_i_1_1), //i
    .port_i_1_2 (stage6_port_i_1_2), //i
    .port_i_1_3 (stage6_port_i_1_3), //i
    .port_i_1_4 (stage6_port_i_1_4), //i
    .port_i_1_5 (stage6_port_i_1_5), //i
    .port_i_1_6 (stage6_port_i_1_6), //i
    .port_i_1_7 (stage6_port_i_1_7), //i
    .port_o_0_0 (stage6_port_o_0_0), //o
    .port_o_0_1 (stage6_port_o_0_1), //o
    .port_o_0_2 (stage6_port_o_0_2), //o
    .port_o_0_3 (stage6_port_o_0_3), //o
    .port_o_0_4 (stage6_port_o_0_4), //o
    .port_o_0_5 (stage6_port_o_0_5), //o
    .port_o_0_6 (stage6_port_o_0_6), //o
    .port_o_0_7 (stage6_port_o_0_7), //o
    .port_o_1_0 (stage6_port_o_1_0), //o
    .port_o_1_1 (stage6_port_o_1_1), //o
    .port_o_1_2 (stage6_port_o_1_2), //o
    .port_o_1_3 (stage6_port_o_1_3), //o
    .port_o_1_4 (stage6_port_o_1_4), //o
    .port_o_1_5 (stage6_port_o_1_5), //o
    .port_o_1_6 (stage6_port_o_1_6), //o
    .port_o_1_7 (stage6_port_o_1_7)  //o
  );
  assign ax_0_0 = stage1_port_o_0_4;
  assign bx_0_0 = stage1_port_o_0_0;
  assign ax_0_1 = stage1_port_o_0_5;
  assign bx_0_1 = stage1_port_o_0_1;
  assign ax_0_2 = stage1_port_o_0_6;
  assign bx_0_2 = stage1_port_o_0_2;
  assign ax_0_3 = stage1_port_o_0_7;
  assign bx_0_3 = stage1_port_o_0_3;
  assign ax_1_0 = stage1_port_o_1_4;
  assign bx_1_0 = stage1_port_o_1_0;
  assign ax_1_1 = stage1_port_o_1_5;
  assign bx_1_1 = stage1_port_o_1_1;
  assign ax_1_2 = stage1_port_o_1_6;
  assign bx_1_2 = stage1_port_o_1_2;
  assign ax_1_3 = stage1_port_o_1_7;
  assign bx_1_3 = stage1_port_o_1_3;
  assign ax1_0_0 = (stage2_port_y_0_2 ^ stage2_port_y_1_2);
  assign ax1_1_0 = (stage2_port_y_2_2 ^ stage2_port_y_3_2);
  assign ax1_0_1 = (stage2_port_y_0_3 ^ stage2_port_y_1_3);
  assign ax1_1_1 = (stage2_port_y_2_3 ^ stage2_port_y_3_3);
  assign bx1_0_0 = (stage2_port_y_0_0 ^ stage2_port_y_1_0);
  assign bx1_1_0 = (stage2_port_y_2_0 ^ stage2_port_y_3_0);
  assign bx1_0_1 = (stage2_port_y_0_1 ^ stage2_port_y_1_1);
  assign bx1_1_1 = (stage2_port_y_2_1 ^ stage2_port_y_3_1);
  assign cx4_0_0 = (stage3_port_y_0_0 ^ stage3_port_y_1_0);
  assign cx4_0_1 = (stage3_port_y_0_1 ^ stage3_port_y_1_1);
  assign cx4_1_0 = (stage3_port_y_2_0 ^ stage3_port_y_3_0);
  assign cx4_1_1 = (stage3_port_y_2_1 ^ stage3_port_y_3_1);
  assign bx5_0_0 = (stage4_port_y_0_0 ^ stage4_port_y_1_0);
  assign bx5_0_1 = (stage4_port_y_0_1 ^ stage4_port_y_1_1);
  assign bx5_0_2 = (stage4_port_y_0_2 ^ stage4_port_y_1_2);
  assign bx5_0_3 = (stage4_port_y_0_3 ^ stage4_port_y_1_3);
  assign bx5_1_0 = (stage4_port_y_2_0 ^ stage4_port_y_3_0);
  assign bx5_1_1 = (stage4_port_y_2_1 ^ stage4_port_y_3_1);
  assign bx5_1_2 = (stage4_port_y_2_2 ^ stage4_port_y_3_2);
  assign bx5_1_3 = (stage4_port_y_2_3 ^ stage4_port_y_3_3);
  assign stage6_port_i_0_0 = (stage5_port_y_0_0 ^ stage5_port_y_1_0);
  assign stage6_port_i_0_1 = (stage5_port_y_0_1 ^ stage5_port_y_1_1);
  assign stage6_port_i_0_2 = (stage5_port_y_0_2 ^ stage5_port_y_1_2);
  assign stage6_port_i_0_3 = (stage5_port_y_0_3 ^ stage5_port_y_1_3);
  assign stage6_port_i_0_4 = (stage5_port_y_0_4 ^ stage5_port_y_1_4);
  assign stage6_port_i_0_5 = (stage5_port_y_0_5 ^ stage5_port_y_1_5);
  assign stage6_port_i_0_6 = (stage5_port_y_0_6 ^ stage5_port_y_1_6);
  assign stage6_port_i_0_7 = (stage5_port_y_0_7 ^ stage5_port_y_1_7);
  assign stage6_port_i_1_0 = (stage5_port_y_2_0 ^ stage5_port_y_3_0);
  assign stage6_port_i_1_1 = (stage5_port_y_2_1 ^ stage5_port_y_3_1);
  assign stage6_port_i_1_2 = (stage5_port_y_2_2 ^ stage5_port_y_3_2);
  assign stage6_port_i_1_3 = (stage5_port_y_2_3 ^ stage5_port_y_3_3);
  assign stage6_port_i_1_4 = (stage5_port_y_2_4 ^ stage5_port_y_3_4);
  assign stage6_port_i_1_5 = (stage5_port_y_2_5 ^ stage5_port_y_3_5);
  assign stage6_port_i_1_6 = (stage5_port_y_2_6 ^ stage5_port_y_3_6);
  assign stage6_port_i_1_7 = (stage5_port_y_2_7 ^ stage5_port_y_3_7);
  assign port_o_0_0 = stage6_port_o_0_0;
  assign port_o_0_1 = stage6_port_o_0_1;
  assign port_o_0_2 = stage6_port_o_0_2;
  assign port_o_0_3 = stage6_port_o_0_3;
  assign port_o_0_4 = stage6_port_o_0_4;
  assign port_o_0_5 = stage6_port_o_0_5;
  assign port_o_0_6 = stage6_port_o_0_6;
  assign port_o_0_7 = stage6_port_o_0_7;
  assign port_o_1_0 = stage6_port_o_1_0;
  assign port_o_1_1 = stage6_port_o_1_1;
  assign port_o_1_2 = stage6_port_o_1_2;
  assign port_o_1_3 = stage6_port_o_1_3;
  assign port_o_1_4 = stage6_port_o_1_4;
  assign port_o_1_5 = stage6_port_o_1_5;
  assign port_o_1_6 = stage6_port_o_1_6;
  assign port_o_1_7 = stage6_port_o_1_7;
  always @(posedge clk) begin
    ax4_0_0 <= ax1_0_0;
    ax4_0_1 <= ax1_0_1;
    ax4_1_0 <= ax1_1_0;
    ax4_1_1 <= ax1_1_1;
    bx4_0_0 <= bx1_0_0;
    bx4_0_1 <= bx1_0_1;
    bx4_1_0 <= bx1_1_0;
    bx4_1_1 <= bx1_1_1;
    ax_reg1_0_0 <= ax_0_0;
    ax_reg1_0_1 <= ax_0_1;
    ax_reg1_0_2 <= ax_0_2;
    ax_reg1_0_3 <= ax_0_3;
    ax_reg1_1_0 <= ax_1_0;
    ax_reg1_1_1 <= ax_1_1;
    ax_reg1_1_2 <= ax_1_2;
    ax_reg1_1_3 <= ax_1_3;
    ax_reg2_0_0 <= ax_reg1_0_0;
    ax_reg2_0_1 <= ax_reg1_0_1;
    ax_reg2_0_2 <= ax_reg1_0_2;
    ax_reg2_0_3 <= ax_reg1_0_3;
    ax_reg2_1_0 <= ax_reg1_1_0;
    ax_reg2_1_1 <= ax_reg1_1_1;
    ax_reg2_1_2 <= ax_reg1_1_2;
    ax_reg2_1_3 <= ax_reg1_1_3;
    ax_reg3_0_0 <= ax_reg2_0_0;
    ax_reg3_0_1 <= ax_reg2_0_1;
    ax_reg3_0_2 <= ax_reg2_0_2;
    ax_reg3_0_3 <= ax_reg2_0_3;
    ax_reg3_1_0 <= ax_reg2_1_0;
    ax_reg3_1_1 <= ax_reg2_1_1;
    ax_reg3_1_2 <= ax_reg2_1_2;
    ax_reg3_1_3 <= ax_reg2_1_3;
    bx_reg1_0_0 <= bx_0_0;
    bx_reg1_0_1 <= bx_0_1;
    bx_reg1_0_2 <= bx_0_2;
    bx_reg1_0_3 <= bx_0_3;
    bx_reg1_1_0 <= bx_1_0;
    bx_reg1_1_1 <= bx_1_1;
    bx_reg1_1_2 <= bx_1_2;
    bx_reg1_1_3 <= bx_1_3;
    bx_reg2_0_0 <= bx_reg1_0_0;
    bx_reg2_0_1 <= bx_reg1_0_1;
    bx_reg2_0_2 <= bx_reg1_0_2;
    bx_reg2_0_3 <= bx_reg1_0_3;
    bx_reg2_1_0 <= bx_reg1_1_0;
    bx_reg2_1_1 <= bx_reg1_1_1;
    bx_reg2_1_2 <= bx_reg1_1_2;
    bx_reg2_1_3 <= bx_reg1_1_3;
    bx_reg3_0_0 <= bx_reg2_0_0;
    bx_reg3_0_1 <= bx_reg2_0_1;
    bx_reg3_0_2 <= bx_reg2_0_2;
    bx_reg3_0_3 <= bx_reg2_0_3;
    bx_reg3_1_0 <= bx_reg2_1_0;
    bx_reg3_1_1 <= bx_reg2_1_1;
    bx_reg3_1_2 <= bx_reg2_1_2;
    bx_reg3_1_3 <= bx_reg2_1_3;
  end


endmodule

module AES_KeyAddition (
  input      [0:0]    port_state_in_0_0_0,
  input      [0:0]    port_state_in_0_0_1,
  input      [0:0]    port_state_in_0_0_2,
  input      [0:0]    port_state_in_0_0_3,
  input      [0:0]    port_state_in_0_0_4,
  input      [0:0]    port_state_in_0_0_5,
  input      [0:0]    port_state_in_0_0_6,
  input      [0:0]    port_state_in_0_0_7,
  input      [0:0]    port_state_in_0_1_0,
  input      [0:0]    port_state_in_0_1_1,
  input      [0:0]    port_state_in_0_1_2,
  input      [0:0]    port_state_in_0_1_3,
  input      [0:0]    port_state_in_0_1_4,
  input      [0:0]    port_state_in_0_1_5,
  input      [0:0]    port_state_in_0_1_6,
  input      [0:0]    port_state_in_0_1_7,
  input      [0:0]    port_state_in_1_0_0,
  input      [0:0]    port_state_in_1_0_1,
  input      [0:0]    port_state_in_1_0_2,
  input      [0:0]    port_state_in_1_0_3,
  input      [0:0]    port_state_in_1_0_4,
  input      [0:0]    port_state_in_1_0_5,
  input      [0:0]    port_state_in_1_0_6,
  input      [0:0]    port_state_in_1_0_7,
  input      [0:0]    port_state_in_1_1_0,
  input      [0:0]    port_state_in_1_1_1,
  input      [0:0]    port_state_in_1_1_2,
  input      [0:0]    port_state_in_1_1_3,
  input      [0:0]    port_state_in_1_1_4,
  input      [0:0]    port_state_in_1_1_5,
  input      [0:0]    port_state_in_1_1_6,
  input      [0:0]    port_state_in_1_1_7,
  input      [0:0]    port_state_in_2_0_0,
  input      [0:0]    port_state_in_2_0_1,
  input      [0:0]    port_state_in_2_0_2,
  input      [0:0]    port_state_in_2_0_3,
  input      [0:0]    port_state_in_2_0_4,
  input      [0:0]    port_state_in_2_0_5,
  input      [0:0]    port_state_in_2_0_6,
  input      [0:0]    port_state_in_2_0_7,
  input      [0:0]    port_state_in_2_1_0,
  input      [0:0]    port_state_in_2_1_1,
  input      [0:0]    port_state_in_2_1_2,
  input      [0:0]    port_state_in_2_1_3,
  input      [0:0]    port_state_in_2_1_4,
  input      [0:0]    port_state_in_2_1_5,
  input      [0:0]    port_state_in_2_1_6,
  input      [0:0]    port_state_in_2_1_7,
  input      [0:0]    port_state_in_3_0_0,
  input      [0:0]    port_state_in_3_0_1,
  input      [0:0]    port_state_in_3_0_2,
  input      [0:0]    port_state_in_3_0_3,
  input      [0:0]    port_state_in_3_0_4,
  input      [0:0]    port_state_in_3_0_5,
  input      [0:0]    port_state_in_3_0_6,
  input      [0:0]    port_state_in_3_0_7,
  input      [0:0]    port_state_in_3_1_0,
  input      [0:0]    port_state_in_3_1_1,
  input      [0:0]    port_state_in_3_1_2,
  input      [0:0]    port_state_in_3_1_3,
  input      [0:0]    port_state_in_3_1_4,
  input      [0:0]    port_state_in_3_1_5,
  input      [0:0]    port_state_in_3_1_6,
  input      [0:0]    port_state_in_3_1_7,
  input      [0:0]    port_state_in_4_0_0,
  input      [0:0]    port_state_in_4_0_1,
  input      [0:0]    port_state_in_4_0_2,
  input      [0:0]    port_state_in_4_0_3,
  input      [0:0]    port_state_in_4_0_4,
  input      [0:0]    port_state_in_4_0_5,
  input      [0:0]    port_state_in_4_0_6,
  input      [0:0]    port_state_in_4_0_7,
  input      [0:0]    port_state_in_4_1_0,
  input      [0:0]    port_state_in_4_1_1,
  input      [0:0]    port_state_in_4_1_2,
  input      [0:0]    port_state_in_4_1_3,
  input      [0:0]    port_state_in_4_1_4,
  input      [0:0]    port_state_in_4_1_5,
  input      [0:0]    port_state_in_4_1_6,
  input      [0:0]    port_state_in_4_1_7,
  input      [0:0]    port_state_in_5_0_0,
  input      [0:0]    port_state_in_5_0_1,
  input      [0:0]    port_state_in_5_0_2,
  input      [0:0]    port_state_in_5_0_3,
  input      [0:0]    port_state_in_5_0_4,
  input      [0:0]    port_state_in_5_0_5,
  input      [0:0]    port_state_in_5_0_6,
  input      [0:0]    port_state_in_5_0_7,
  input      [0:0]    port_state_in_5_1_0,
  input      [0:0]    port_state_in_5_1_1,
  input      [0:0]    port_state_in_5_1_2,
  input      [0:0]    port_state_in_5_1_3,
  input      [0:0]    port_state_in_5_1_4,
  input      [0:0]    port_state_in_5_1_5,
  input      [0:0]    port_state_in_5_1_6,
  input      [0:0]    port_state_in_5_1_7,
  input      [0:0]    port_state_in_6_0_0,
  input      [0:0]    port_state_in_6_0_1,
  input      [0:0]    port_state_in_6_0_2,
  input      [0:0]    port_state_in_6_0_3,
  input      [0:0]    port_state_in_6_0_4,
  input      [0:0]    port_state_in_6_0_5,
  input      [0:0]    port_state_in_6_0_6,
  input      [0:0]    port_state_in_6_0_7,
  input      [0:0]    port_state_in_6_1_0,
  input      [0:0]    port_state_in_6_1_1,
  input      [0:0]    port_state_in_6_1_2,
  input      [0:0]    port_state_in_6_1_3,
  input      [0:0]    port_state_in_6_1_4,
  input      [0:0]    port_state_in_6_1_5,
  input      [0:0]    port_state_in_6_1_6,
  input      [0:0]    port_state_in_6_1_7,
  input      [0:0]    port_state_in_7_0_0,
  input      [0:0]    port_state_in_7_0_1,
  input      [0:0]    port_state_in_7_0_2,
  input      [0:0]    port_state_in_7_0_3,
  input      [0:0]    port_state_in_7_0_4,
  input      [0:0]    port_state_in_7_0_5,
  input      [0:0]    port_state_in_7_0_6,
  input      [0:0]    port_state_in_7_0_7,
  input      [0:0]    port_state_in_7_1_0,
  input      [0:0]    port_state_in_7_1_1,
  input      [0:0]    port_state_in_7_1_2,
  input      [0:0]    port_state_in_7_1_3,
  input      [0:0]    port_state_in_7_1_4,
  input      [0:0]    port_state_in_7_1_5,
  input      [0:0]    port_state_in_7_1_6,
  input      [0:0]    port_state_in_7_1_7,
  input      [0:0]    port_state_in_8_0_0,
  input      [0:0]    port_state_in_8_0_1,
  input      [0:0]    port_state_in_8_0_2,
  input      [0:0]    port_state_in_8_0_3,
  input      [0:0]    port_state_in_8_0_4,
  input      [0:0]    port_state_in_8_0_5,
  input      [0:0]    port_state_in_8_0_6,
  input      [0:0]    port_state_in_8_0_7,
  input      [0:0]    port_state_in_8_1_0,
  input      [0:0]    port_state_in_8_1_1,
  input      [0:0]    port_state_in_8_1_2,
  input      [0:0]    port_state_in_8_1_3,
  input      [0:0]    port_state_in_8_1_4,
  input      [0:0]    port_state_in_8_1_5,
  input      [0:0]    port_state_in_8_1_6,
  input      [0:0]    port_state_in_8_1_7,
  input      [0:0]    port_state_in_9_0_0,
  input      [0:0]    port_state_in_9_0_1,
  input      [0:0]    port_state_in_9_0_2,
  input      [0:0]    port_state_in_9_0_3,
  input      [0:0]    port_state_in_9_0_4,
  input      [0:0]    port_state_in_9_0_5,
  input      [0:0]    port_state_in_9_0_6,
  input      [0:0]    port_state_in_9_0_7,
  input      [0:0]    port_state_in_9_1_0,
  input      [0:0]    port_state_in_9_1_1,
  input      [0:0]    port_state_in_9_1_2,
  input      [0:0]    port_state_in_9_1_3,
  input      [0:0]    port_state_in_9_1_4,
  input      [0:0]    port_state_in_9_1_5,
  input      [0:0]    port_state_in_9_1_6,
  input      [0:0]    port_state_in_9_1_7,
  input      [0:0]    port_state_in_10_0_0,
  input      [0:0]    port_state_in_10_0_1,
  input      [0:0]    port_state_in_10_0_2,
  input      [0:0]    port_state_in_10_0_3,
  input      [0:0]    port_state_in_10_0_4,
  input      [0:0]    port_state_in_10_0_5,
  input      [0:0]    port_state_in_10_0_6,
  input      [0:0]    port_state_in_10_0_7,
  input      [0:0]    port_state_in_10_1_0,
  input      [0:0]    port_state_in_10_1_1,
  input      [0:0]    port_state_in_10_1_2,
  input      [0:0]    port_state_in_10_1_3,
  input      [0:0]    port_state_in_10_1_4,
  input      [0:0]    port_state_in_10_1_5,
  input      [0:0]    port_state_in_10_1_6,
  input      [0:0]    port_state_in_10_1_7,
  input      [0:0]    port_state_in_11_0_0,
  input      [0:0]    port_state_in_11_0_1,
  input      [0:0]    port_state_in_11_0_2,
  input      [0:0]    port_state_in_11_0_3,
  input      [0:0]    port_state_in_11_0_4,
  input      [0:0]    port_state_in_11_0_5,
  input      [0:0]    port_state_in_11_0_6,
  input      [0:0]    port_state_in_11_0_7,
  input      [0:0]    port_state_in_11_1_0,
  input      [0:0]    port_state_in_11_1_1,
  input      [0:0]    port_state_in_11_1_2,
  input      [0:0]    port_state_in_11_1_3,
  input      [0:0]    port_state_in_11_1_4,
  input      [0:0]    port_state_in_11_1_5,
  input      [0:0]    port_state_in_11_1_6,
  input      [0:0]    port_state_in_11_1_7,
  input      [0:0]    port_state_in_12_0_0,
  input      [0:0]    port_state_in_12_0_1,
  input      [0:0]    port_state_in_12_0_2,
  input      [0:0]    port_state_in_12_0_3,
  input      [0:0]    port_state_in_12_0_4,
  input      [0:0]    port_state_in_12_0_5,
  input      [0:0]    port_state_in_12_0_6,
  input      [0:0]    port_state_in_12_0_7,
  input      [0:0]    port_state_in_12_1_0,
  input      [0:0]    port_state_in_12_1_1,
  input      [0:0]    port_state_in_12_1_2,
  input      [0:0]    port_state_in_12_1_3,
  input      [0:0]    port_state_in_12_1_4,
  input      [0:0]    port_state_in_12_1_5,
  input      [0:0]    port_state_in_12_1_6,
  input      [0:0]    port_state_in_12_1_7,
  input      [0:0]    port_state_in_13_0_0,
  input      [0:0]    port_state_in_13_0_1,
  input      [0:0]    port_state_in_13_0_2,
  input      [0:0]    port_state_in_13_0_3,
  input      [0:0]    port_state_in_13_0_4,
  input      [0:0]    port_state_in_13_0_5,
  input      [0:0]    port_state_in_13_0_6,
  input      [0:0]    port_state_in_13_0_7,
  input      [0:0]    port_state_in_13_1_0,
  input      [0:0]    port_state_in_13_1_1,
  input      [0:0]    port_state_in_13_1_2,
  input      [0:0]    port_state_in_13_1_3,
  input      [0:0]    port_state_in_13_1_4,
  input      [0:0]    port_state_in_13_1_5,
  input      [0:0]    port_state_in_13_1_6,
  input      [0:0]    port_state_in_13_1_7,
  input      [0:0]    port_state_in_14_0_0,
  input      [0:0]    port_state_in_14_0_1,
  input      [0:0]    port_state_in_14_0_2,
  input      [0:0]    port_state_in_14_0_3,
  input      [0:0]    port_state_in_14_0_4,
  input      [0:0]    port_state_in_14_0_5,
  input      [0:0]    port_state_in_14_0_6,
  input      [0:0]    port_state_in_14_0_7,
  input      [0:0]    port_state_in_14_1_0,
  input      [0:0]    port_state_in_14_1_1,
  input      [0:0]    port_state_in_14_1_2,
  input      [0:0]    port_state_in_14_1_3,
  input      [0:0]    port_state_in_14_1_4,
  input      [0:0]    port_state_in_14_1_5,
  input      [0:0]    port_state_in_14_1_6,
  input      [0:0]    port_state_in_14_1_7,
  input      [0:0]    port_state_in_15_0_0,
  input      [0:0]    port_state_in_15_0_1,
  input      [0:0]    port_state_in_15_0_2,
  input      [0:0]    port_state_in_15_0_3,
  input      [0:0]    port_state_in_15_0_4,
  input      [0:0]    port_state_in_15_0_5,
  input      [0:0]    port_state_in_15_0_6,
  input      [0:0]    port_state_in_15_0_7,
  input      [0:0]    port_state_in_15_1_0,
  input      [0:0]    port_state_in_15_1_1,
  input      [0:0]    port_state_in_15_1_2,
  input      [0:0]    port_state_in_15_1_3,
  input      [0:0]    port_state_in_15_1_4,
  input      [0:0]    port_state_in_15_1_5,
  input      [0:0]    port_state_in_15_1_6,
  input      [0:0]    port_state_in_15_1_7,
  input      [0:0]    port_key_0_0_0,
  input      [0:0]    port_key_0_0_1,
  input      [0:0]    port_key_0_0_2,
  input      [0:0]    port_key_0_0_3,
  input      [0:0]    port_key_0_0_4,
  input      [0:0]    port_key_0_0_5,
  input      [0:0]    port_key_0_0_6,
  input      [0:0]    port_key_0_0_7,
  input      [0:0]    port_key_0_1_0,
  input      [0:0]    port_key_0_1_1,
  input      [0:0]    port_key_0_1_2,
  input      [0:0]    port_key_0_1_3,
  input      [0:0]    port_key_0_1_4,
  input      [0:0]    port_key_0_1_5,
  input      [0:0]    port_key_0_1_6,
  input      [0:0]    port_key_0_1_7,
  input      [0:0]    port_key_1_0_0,
  input      [0:0]    port_key_1_0_1,
  input      [0:0]    port_key_1_0_2,
  input      [0:0]    port_key_1_0_3,
  input      [0:0]    port_key_1_0_4,
  input      [0:0]    port_key_1_0_5,
  input      [0:0]    port_key_1_0_6,
  input      [0:0]    port_key_1_0_7,
  input      [0:0]    port_key_1_1_0,
  input      [0:0]    port_key_1_1_1,
  input      [0:0]    port_key_1_1_2,
  input      [0:0]    port_key_1_1_3,
  input      [0:0]    port_key_1_1_4,
  input      [0:0]    port_key_1_1_5,
  input      [0:0]    port_key_1_1_6,
  input      [0:0]    port_key_1_1_7,
  input      [0:0]    port_key_2_0_0,
  input      [0:0]    port_key_2_0_1,
  input      [0:0]    port_key_2_0_2,
  input      [0:0]    port_key_2_0_3,
  input      [0:0]    port_key_2_0_4,
  input      [0:0]    port_key_2_0_5,
  input      [0:0]    port_key_2_0_6,
  input      [0:0]    port_key_2_0_7,
  input      [0:0]    port_key_2_1_0,
  input      [0:0]    port_key_2_1_1,
  input      [0:0]    port_key_2_1_2,
  input      [0:0]    port_key_2_1_3,
  input      [0:0]    port_key_2_1_4,
  input      [0:0]    port_key_2_1_5,
  input      [0:0]    port_key_2_1_6,
  input      [0:0]    port_key_2_1_7,
  input      [0:0]    port_key_3_0_0,
  input      [0:0]    port_key_3_0_1,
  input      [0:0]    port_key_3_0_2,
  input      [0:0]    port_key_3_0_3,
  input      [0:0]    port_key_3_0_4,
  input      [0:0]    port_key_3_0_5,
  input      [0:0]    port_key_3_0_6,
  input      [0:0]    port_key_3_0_7,
  input      [0:0]    port_key_3_1_0,
  input      [0:0]    port_key_3_1_1,
  input      [0:0]    port_key_3_1_2,
  input      [0:0]    port_key_3_1_3,
  input      [0:0]    port_key_3_1_4,
  input      [0:0]    port_key_3_1_5,
  input      [0:0]    port_key_3_1_6,
  input      [0:0]    port_key_3_1_7,
  input      [0:0]    port_key_4_0_0,
  input      [0:0]    port_key_4_0_1,
  input      [0:0]    port_key_4_0_2,
  input      [0:0]    port_key_4_0_3,
  input      [0:0]    port_key_4_0_4,
  input      [0:0]    port_key_4_0_5,
  input      [0:0]    port_key_4_0_6,
  input      [0:0]    port_key_4_0_7,
  input      [0:0]    port_key_4_1_0,
  input      [0:0]    port_key_4_1_1,
  input      [0:0]    port_key_4_1_2,
  input      [0:0]    port_key_4_1_3,
  input      [0:0]    port_key_4_1_4,
  input      [0:0]    port_key_4_1_5,
  input      [0:0]    port_key_4_1_6,
  input      [0:0]    port_key_4_1_7,
  input      [0:0]    port_key_5_0_0,
  input      [0:0]    port_key_5_0_1,
  input      [0:0]    port_key_5_0_2,
  input      [0:0]    port_key_5_0_3,
  input      [0:0]    port_key_5_0_4,
  input      [0:0]    port_key_5_0_5,
  input      [0:0]    port_key_5_0_6,
  input      [0:0]    port_key_5_0_7,
  input      [0:0]    port_key_5_1_0,
  input      [0:0]    port_key_5_1_1,
  input      [0:0]    port_key_5_1_2,
  input      [0:0]    port_key_5_1_3,
  input      [0:0]    port_key_5_1_4,
  input      [0:0]    port_key_5_1_5,
  input      [0:0]    port_key_5_1_6,
  input      [0:0]    port_key_5_1_7,
  input      [0:0]    port_key_6_0_0,
  input      [0:0]    port_key_6_0_1,
  input      [0:0]    port_key_6_0_2,
  input      [0:0]    port_key_6_0_3,
  input      [0:0]    port_key_6_0_4,
  input      [0:0]    port_key_6_0_5,
  input      [0:0]    port_key_6_0_6,
  input      [0:0]    port_key_6_0_7,
  input      [0:0]    port_key_6_1_0,
  input      [0:0]    port_key_6_1_1,
  input      [0:0]    port_key_6_1_2,
  input      [0:0]    port_key_6_1_3,
  input      [0:0]    port_key_6_1_4,
  input      [0:0]    port_key_6_1_5,
  input      [0:0]    port_key_6_1_6,
  input      [0:0]    port_key_6_1_7,
  input      [0:0]    port_key_7_0_0,
  input      [0:0]    port_key_7_0_1,
  input      [0:0]    port_key_7_0_2,
  input      [0:0]    port_key_7_0_3,
  input      [0:0]    port_key_7_0_4,
  input      [0:0]    port_key_7_0_5,
  input      [0:0]    port_key_7_0_6,
  input      [0:0]    port_key_7_0_7,
  input      [0:0]    port_key_7_1_0,
  input      [0:0]    port_key_7_1_1,
  input      [0:0]    port_key_7_1_2,
  input      [0:0]    port_key_7_1_3,
  input      [0:0]    port_key_7_1_4,
  input      [0:0]    port_key_7_1_5,
  input      [0:0]    port_key_7_1_6,
  input      [0:0]    port_key_7_1_7,
  input      [0:0]    port_key_8_0_0,
  input      [0:0]    port_key_8_0_1,
  input      [0:0]    port_key_8_0_2,
  input      [0:0]    port_key_8_0_3,
  input      [0:0]    port_key_8_0_4,
  input      [0:0]    port_key_8_0_5,
  input      [0:0]    port_key_8_0_6,
  input      [0:0]    port_key_8_0_7,
  input      [0:0]    port_key_8_1_0,
  input      [0:0]    port_key_8_1_1,
  input      [0:0]    port_key_8_1_2,
  input      [0:0]    port_key_8_1_3,
  input      [0:0]    port_key_8_1_4,
  input      [0:0]    port_key_8_1_5,
  input      [0:0]    port_key_8_1_6,
  input      [0:0]    port_key_8_1_7,
  input      [0:0]    port_key_9_0_0,
  input      [0:0]    port_key_9_0_1,
  input      [0:0]    port_key_9_0_2,
  input      [0:0]    port_key_9_0_3,
  input      [0:0]    port_key_9_0_4,
  input      [0:0]    port_key_9_0_5,
  input      [0:0]    port_key_9_0_6,
  input      [0:0]    port_key_9_0_7,
  input      [0:0]    port_key_9_1_0,
  input      [0:0]    port_key_9_1_1,
  input      [0:0]    port_key_9_1_2,
  input      [0:0]    port_key_9_1_3,
  input      [0:0]    port_key_9_1_4,
  input      [0:0]    port_key_9_1_5,
  input      [0:0]    port_key_9_1_6,
  input      [0:0]    port_key_9_1_7,
  input      [0:0]    port_key_10_0_0,
  input      [0:0]    port_key_10_0_1,
  input      [0:0]    port_key_10_0_2,
  input      [0:0]    port_key_10_0_3,
  input      [0:0]    port_key_10_0_4,
  input      [0:0]    port_key_10_0_5,
  input      [0:0]    port_key_10_0_6,
  input      [0:0]    port_key_10_0_7,
  input      [0:0]    port_key_10_1_0,
  input      [0:0]    port_key_10_1_1,
  input      [0:0]    port_key_10_1_2,
  input      [0:0]    port_key_10_1_3,
  input      [0:0]    port_key_10_1_4,
  input      [0:0]    port_key_10_1_5,
  input      [0:0]    port_key_10_1_6,
  input      [0:0]    port_key_10_1_7,
  input      [0:0]    port_key_11_0_0,
  input      [0:0]    port_key_11_0_1,
  input      [0:0]    port_key_11_0_2,
  input      [0:0]    port_key_11_0_3,
  input      [0:0]    port_key_11_0_4,
  input      [0:0]    port_key_11_0_5,
  input      [0:0]    port_key_11_0_6,
  input      [0:0]    port_key_11_0_7,
  input      [0:0]    port_key_11_1_0,
  input      [0:0]    port_key_11_1_1,
  input      [0:0]    port_key_11_1_2,
  input      [0:0]    port_key_11_1_3,
  input      [0:0]    port_key_11_1_4,
  input      [0:0]    port_key_11_1_5,
  input      [0:0]    port_key_11_1_6,
  input      [0:0]    port_key_11_1_7,
  input      [0:0]    port_key_12_0_0,
  input      [0:0]    port_key_12_0_1,
  input      [0:0]    port_key_12_0_2,
  input      [0:0]    port_key_12_0_3,
  input      [0:0]    port_key_12_0_4,
  input      [0:0]    port_key_12_0_5,
  input      [0:0]    port_key_12_0_6,
  input      [0:0]    port_key_12_0_7,
  input      [0:0]    port_key_12_1_0,
  input      [0:0]    port_key_12_1_1,
  input      [0:0]    port_key_12_1_2,
  input      [0:0]    port_key_12_1_3,
  input      [0:0]    port_key_12_1_4,
  input      [0:0]    port_key_12_1_5,
  input      [0:0]    port_key_12_1_6,
  input      [0:0]    port_key_12_1_7,
  input      [0:0]    port_key_13_0_0,
  input      [0:0]    port_key_13_0_1,
  input      [0:0]    port_key_13_0_2,
  input      [0:0]    port_key_13_0_3,
  input      [0:0]    port_key_13_0_4,
  input      [0:0]    port_key_13_0_5,
  input      [0:0]    port_key_13_0_6,
  input      [0:0]    port_key_13_0_7,
  input      [0:0]    port_key_13_1_0,
  input      [0:0]    port_key_13_1_1,
  input      [0:0]    port_key_13_1_2,
  input      [0:0]    port_key_13_1_3,
  input      [0:0]    port_key_13_1_4,
  input      [0:0]    port_key_13_1_5,
  input      [0:0]    port_key_13_1_6,
  input      [0:0]    port_key_13_1_7,
  input      [0:0]    port_key_14_0_0,
  input      [0:0]    port_key_14_0_1,
  input      [0:0]    port_key_14_0_2,
  input      [0:0]    port_key_14_0_3,
  input      [0:0]    port_key_14_0_4,
  input      [0:0]    port_key_14_0_5,
  input      [0:0]    port_key_14_0_6,
  input      [0:0]    port_key_14_0_7,
  input      [0:0]    port_key_14_1_0,
  input      [0:0]    port_key_14_1_1,
  input      [0:0]    port_key_14_1_2,
  input      [0:0]    port_key_14_1_3,
  input      [0:0]    port_key_14_1_4,
  input      [0:0]    port_key_14_1_5,
  input      [0:0]    port_key_14_1_6,
  input      [0:0]    port_key_14_1_7,
  input      [0:0]    port_key_15_0_0,
  input      [0:0]    port_key_15_0_1,
  input      [0:0]    port_key_15_0_2,
  input      [0:0]    port_key_15_0_3,
  input      [0:0]    port_key_15_0_4,
  input      [0:0]    port_key_15_0_5,
  input      [0:0]    port_key_15_0_6,
  input      [0:0]    port_key_15_0_7,
  input      [0:0]    port_key_15_1_0,
  input      [0:0]    port_key_15_1_1,
  input      [0:0]    port_key_15_1_2,
  input      [0:0]    port_key_15_1_3,
  input      [0:0]    port_key_15_1_4,
  input      [0:0]    port_key_15_1_5,
  input      [0:0]    port_key_15_1_6,
  input      [0:0]    port_key_15_1_7,
  output     [0:0]    port_state_out_0_0_0,
  output     [0:0]    port_state_out_0_0_1,
  output     [0:0]    port_state_out_0_0_2,
  output     [0:0]    port_state_out_0_0_3,
  output     [0:0]    port_state_out_0_0_4,
  output     [0:0]    port_state_out_0_0_5,
  output     [0:0]    port_state_out_0_0_6,
  output     [0:0]    port_state_out_0_0_7,
  output     [0:0]    port_state_out_0_1_0,
  output     [0:0]    port_state_out_0_1_1,
  output     [0:0]    port_state_out_0_1_2,
  output     [0:0]    port_state_out_0_1_3,
  output     [0:0]    port_state_out_0_1_4,
  output     [0:0]    port_state_out_0_1_5,
  output     [0:0]    port_state_out_0_1_6,
  output     [0:0]    port_state_out_0_1_7,
  output     [0:0]    port_state_out_1_0_0,
  output     [0:0]    port_state_out_1_0_1,
  output     [0:0]    port_state_out_1_0_2,
  output     [0:0]    port_state_out_1_0_3,
  output     [0:0]    port_state_out_1_0_4,
  output     [0:0]    port_state_out_1_0_5,
  output     [0:0]    port_state_out_1_0_6,
  output     [0:0]    port_state_out_1_0_7,
  output     [0:0]    port_state_out_1_1_0,
  output     [0:0]    port_state_out_1_1_1,
  output     [0:0]    port_state_out_1_1_2,
  output     [0:0]    port_state_out_1_1_3,
  output     [0:0]    port_state_out_1_1_4,
  output     [0:0]    port_state_out_1_1_5,
  output     [0:0]    port_state_out_1_1_6,
  output     [0:0]    port_state_out_1_1_7,
  output     [0:0]    port_state_out_2_0_0,
  output     [0:0]    port_state_out_2_0_1,
  output     [0:0]    port_state_out_2_0_2,
  output     [0:0]    port_state_out_2_0_3,
  output     [0:0]    port_state_out_2_0_4,
  output     [0:0]    port_state_out_2_0_5,
  output     [0:0]    port_state_out_2_0_6,
  output     [0:0]    port_state_out_2_0_7,
  output     [0:0]    port_state_out_2_1_0,
  output     [0:0]    port_state_out_2_1_1,
  output     [0:0]    port_state_out_2_1_2,
  output     [0:0]    port_state_out_2_1_3,
  output     [0:0]    port_state_out_2_1_4,
  output     [0:0]    port_state_out_2_1_5,
  output     [0:0]    port_state_out_2_1_6,
  output     [0:0]    port_state_out_2_1_7,
  output     [0:0]    port_state_out_3_0_0,
  output     [0:0]    port_state_out_3_0_1,
  output     [0:0]    port_state_out_3_0_2,
  output     [0:0]    port_state_out_3_0_3,
  output     [0:0]    port_state_out_3_0_4,
  output     [0:0]    port_state_out_3_0_5,
  output     [0:0]    port_state_out_3_0_6,
  output     [0:0]    port_state_out_3_0_7,
  output     [0:0]    port_state_out_3_1_0,
  output     [0:0]    port_state_out_3_1_1,
  output     [0:0]    port_state_out_3_1_2,
  output     [0:0]    port_state_out_3_1_3,
  output     [0:0]    port_state_out_3_1_4,
  output     [0:0]    port_state_out_3_1_5,
  output     [0:0]    port_state_out_3_1_6,
  output     [0:0]    port_state_out_3_1_7,
  output     [0:0]    port_state_out_4_0_0,
  output     [0:0]    port_state_out_4_0_1,
  output     [0:0]    port_state_out_4_0_2,
  output     [0:0]    port_state_out_4_0_3,
  output     [0:0]    port_state_out_4_0_4,
  output     [0:0]    port_state_out_4_0_5,
  output     [0:0]    port_state_out_4_0_6,
  output     [0:0]    port_state_out_4_0_7,
  output     [0:0]    port_state_out_4_1_0,
  output     [0:0]    port_state_out_4_1_1,
  output     [0:0]    port_state_out_4_1_2,
  output     [0:0]    port_state_out_4_1_3,
  output     [0:0]    port_state_out_4_1_4,
  output     [0:0]    port_state_out_4_1_5,
  output     [0:0]    port_state_out_4_1_6,
  output     [0:0]    port_state_out_4_1_7,
  output     [0:0]    port_state_out_5_0_0,
  output     [0:0]    port_state_out_5_0_1,
  output     [0:0]    port_state_out_5_0_2,
  output     [0:0]    port_state_out_5_0_3,
  output     [0:0]    port_state_out_5_0_4,
  output     [0:0]    port_state_out_5_0_5,
  output     [0:0]    port_state_out_5_0_6,
  output     [0:0]    port_state_out_5_0_7,
  output     [0:0]    port_state_out_5_1_0,
  output     [0:0]    port_state_out_5_1_1,
  output     [0:0]    port_state_out_5_1_2,
  output     [0:0]    port_state_out_5_1_3,
  output     [0:0]    port_state_out_5_1_4,
  output     [0:0]    port_state_out_5_1_5,
  output     [0:0]    port_state_out_5_1_6,
  output     [0:0]    port_state_out_5_1_7,
  output     [0:0]    port_state_out_6_0_0,
  output     [0:0]    port_state_out_6_0_1,
  output     [0:0]    port_state_out_6_0_2,
  output     [0:0]    port_state_out_6_0_3,
  output     [0:0]    port_state_out_6_0_4,
  output     [0:0]    port_state_out_6_0_5,
  output     [0:0]    port_state_out_6_0_6,
  output     [0:0]    port_state_out_6_0_7,
  output     [0:0]    port_state_out_6_1_0,
  output     [0:0]    port_state_out_6_1_1,
  output     [0:0]    port_state_out_6_1_2,
  output     [0:0]    port_state_out_6_1_3,
  output     [0:0]    port_state_out_6_1_4,
  output     [0:0]    port_state_out_6_1_5,
  output     [0:0]    port_state_out_6_1_6,
  output     [0:0]    port_state_out_6_1_7,
  output     [0:0]    port_state_out_7_0_0,
  output     [0:0]    port_state_out_7_0_1,
  output     [0:0]    port_state_out_7_0_2,
  output     [0:0]    port_state_out_7_0_3,
  output     [0:0]    port_state_out_7_0_4,
  output     [0:0]    port_state_out_7_0_5,
  output     [0:0]    port_state_out_7_0_6,
  output     [0:0]    port_state_out_7_0_7,
  output     [0:0]    port_state_out_7_1_0,
  output     [0:0]    port_state_out_7_1_1,
  output     [0:0]    port_state_out_7_1_2,
  output     [0:0]    port_state_out_7_1_3,
  output     [0:0]    port_state_out_7_1_4,
  output     [0:0]    port_state_out_7_1_5,
  output     [0:0]    port_state_out_7_1_6,
  output     [0:0]    port_state_out_7_1_7,
  output     [0:0]    port_state_out_8_0_0,
  output     [0:0]    port_state_out_8_0_1,
  output     [0:0]    port_state_out_8_0_2,
  output     [0:0]    port_state_out_8_0_3,
  output     [0:0]    port_state_out_8_0_4,
  output     [0:0]    port_state_out_8_0_5,
  output     [0:0]    port_state_out_8_0_6,
  output     [0:0]    port_state_out_8_0_7,
  output     [0:0]    port_state_out_8_1_0,
  output     [0:0]    port_state_out_8_1_1,
  output     [0:0]    port_state_out_8_1_2,
  output     [0:0]    port_state_out_8_1_3,
  output     [0:0]    port_state_out_8_1_4,
  output     [0:0]    port_state_out_8_1_5,
  output     [0:0]    port_state_out_8_1_6,
  output     [0:0]    port_state_out_8_1_7,
  output     [0:0]    port_state_out_9_0_0,
  output     [0:0]    port_state_out_9_0_1,
  output     [0:0]    port_state_out_9_0_2,
  output     [0:0]    port_state_out_9_0_3,
  output     [0:0]    port_state_out_9_0_4,
  output     [0:0]    port_state_out_9_0_5,
  output     [0:0]    port_state_out_9_0_6,
  output     [0:0]    port_state_out_9_0_7,
  output     [0:0]    port_state_out_9_1_0,
  output     [0:0]    port_state_out_9_1_1,
  output     [0:0]    port_state_out_9_1_2,
  output     [0:0]    port_state_out_9_1_3,
  output     [0:0]    port_state_out_9_1_4,
  output     [0:0]    port_state_out_9_1_5,
  output     [0:0]    port_state_out_9_1_6,
  output     [0:0]    port_state_out_9_1_7,
  output     [0:0]    port_state_out_10_0_0,
  output     [0:0]    port_state_out_10_0_1,
  output     [0:0]    port_state_out_10_0_2,
  output     [0:0]    port_state_out_10_0_3,
  output     [0:0]    port_state_out_10_0_4,
  output     [0:0]    port_state_out_10_0_5,
  output     [0:0]    port_state_out_10_0_6,
  output     [0:0]    port_state_out_10_0_7,
  output     [0:0]    port_state_out_10_1_0,
  output     [0:0]    port_state_out_10_1_1,
  output     [0:0]    port_state_out_10_1_2,
  output     [0:0]    port_state_out_10_1_3,
  output     [0:0]    port_state_out_10_1_4,
  output     [0:0]    port_state_out_10_1_5,
  output     [0:0]    port_state_out_10_1_6,
  output     [0:0]    port_state_out_10_1_7,
  output     [0:0]    port_state_out_11_0_0,
  output     [0:0]    port_state_out_11_0_1,
  output     [0:0]    port_state_out_11_0_2,
  output     [0:0]    port_state_out_11_0_3,
  output     [0:0]    port_state_out_11_0_4,
  output     [0:0]    port_state_out_11_0_5,
  output     [0:0]    port_state_out_11_0_6,
  output     [0:0]    port_state_out_11_0_7,
  output     [0:0]    port_state_out_11_1_0,
  output     [0:0]    port_state_out_11_1_1,
  output     [0:0]    port_state_out_11_1_2,
  output     [0:0]    port_state_out_11_1_3,
  output     [0:0]    port_state_out_11_1_4,
  output     [0:0]    port_state_out_11_1_5,
  output     [0:0]    port_state_out_11_1_6,
  output     [0:0]    port_state_out_11_1_7,
  output     [0:0]    port_state_out_12_0_0,
  output     [0:0]    port_state_out_12_0_1,
  output     [0:0]    port_state_out_12_0_2,
  output     [0:0]    port_state_out_12_0_3,
  output     [0:0]    port_state_out_12_0_4,
  output     [0:0]    port_state_out_12_0_5,
  output     [0:0]    port_state_out_12_0_6,
  output     [0:0]    port_state_out_12_0_7,
  output     [0:0]    port_state_out_12_1_0,
  output     [0:0]    port_state_out_12_1_1,
  output     [0:0]    port_state_out_12_1_2,
  output     [0:0]    port_state_out_12_1_3,
  output     [0:0]    port_state_out_12_1_4,
  output     [0:0]    port_state_out_12_1_5,
  output     [0:0]    port_state_out_12_1_6,
  output     [0:0]    port_state_out_12_1_7,
  output     [0:0]    port_state_out_13_0_0,
  output     [0:0]    port_state_out_13_0_1,
  output     [0:0]    port_state_out_13_0_2,
  output     [0:0]    port_state_out_13_0_3,
  output     [0:0]    port_state_out_13_0_4,
  output     [0:0]    port_state_out_13_0_5,
  output     [0:0]    port_state_out_13_0_6,
  output     [0:0]    port_state_out_13_0_7,
  output     [0:0]    port_state_out_13_1_0,
  output     [0:0]    port_state_out_13_1_1,
  output     [0:0]    port_state_out_13_1_2,
  output     [0:0]    port_state_out_13_1_3,
  output     [0:0]    port_state_out_13_1_4,
  output     [0:0]    port_state_out_13_1_5,
  output     [0:0]    port_state_out_13_1_6,
  output     [0:0]    port_state_out_13_1_7,
  output     [0:0]    port_state_out_14_0_0,
  output     [0:0]    port_state_out_14_0_1,
  output     [0:0]    port_state_out_14_0_2,
  output     [0:0]    port_state_out_14_0_3,
  output     [0:0]    port_state_out_14_0_4,
  output     [0:0]    port_state_out_14_0_5,
  output     [0:0]    port_state_out_14_0_6,
  output     [0:0]    port_state_out_14_0_7,
  output     [0:0]    port_state_out_14_1_0,
  output     [0:0]    port_state_out_14_1_1,
  output     [0:0]    port_state_out_14_1_2,
  output     [0:0]    port_state_out_14_1_3,
  output     [0:0]    port_state_out_14_1_4,
  output     [0:0]    port_state_out_14_1_5,
  output     [0:0]    port_state_out_14_1_6,
  output     [0:0]    port_state_out_14_1_7,
  output     [0:0]    port_state_out_15_0_0,
  output     [0:0]    port_state_out_15_0_1,
  output     [0:0]    port_state_out_15_0_2,
  output     [0:0]    port_state_out_15_0_3,
  output     [0:0]    port_state_out_15_0_4,
  output     [0:0]    port_state_out_15_0_5,
  output     [0:0]    port_state_out_15_0_6,
  output     [0:0]    port_state_out_15_0_7,
  output     [0:0]    port_state_out_15_1_0,
  output     [0:0]    port_state_out_15_1_1,
  output     [0:0]    port_state_out_15_1_2,
  output     [0:0]    port_state_out_15_1_3,
  output     [0:0]    port_state_out_15_1_4,
  output     [0:0]    port_state_out_15_1_5,
  output     [0:0]    port_state_out_15_1_6,
  output     [0:0]    port_state_out_15_1_7
);


  assign port_state_out_0_0_0 = (port_state_in_0_0_0 ^ port_key_0_0_0);
  assign port_state_out_0_0_1 = (port_state_in_0_0_1 ^ port_key_0_0_1);
  assign port_state_out_0_0_2 = (port_state_in_0_0_2 ^ port_key_0_0_2);
  assign port_state_out_0_0_3 = (port_state_in_0_0_3 ^ port_key_0_0_3);
  assign port_state_out_0_0_4 = (port_state_in_0_0_4 ^ port_key_0_0_4);
  assign port_state_out_0_0_5 = (port_state_in_0_0_5 ^ port_key_0_0_5);
  assign port_state_out_0_0_6 = (port_state_in_0_0_6 ^ port_key_0_0_6);
  assign port_state_out_0_0_7 = (port_state_in_0_0_7 ^ port_key_0_0_7);
  assign port_state_out_0_1_0 = (port_state_in_0_1_0 ^ port_key_0_1_0);
  assign port_state_out_0_1_1 = (port_state_in_0_1_1 ^ port_key_0_1_1);
  assign port_state_out_0_1_2 = (port_state_in_0_1_2 ^ port_key_0_1_2);
  assign port_state_out_0_1_3 = (port_state_in_0_1_3 ^ port_key_0_1_3);
  assign port_state_out_0_1_4 = (port_state_in_0_1_4 ^ port_key_0_1_4);
  assign port_state_out_0_1_5 = (port_state_in_0_1_5 ^ port_key_0_1_5);
  assign port_state_out_0_1_6 = (port_state_in_0_1_6 ^ port_key_0_1_6);
  assign port_state_out_0_1_7 = (port_state_in_0_1_7 ^ port_key_0_1_7);
  assign port_state_out_1_0_0 = (port_state_in_1_0_0 ^ port_key_1_0_0);
  assign port_state_out_1_0_1 = (port_state_in_1_0_1 ^ port_key_1_0_1);
  assign port_state_out_1_0_2 = (port_state_in_1_0_2 ^ port_key_1_0_2);
  assign port_state_out_1_0_3 = (port_state_in_1_0_3 ^ port_key_1_0_3);
  assign port_state_out_1_0_4 = (port_state_in_1_0_4 ^ port_key_1_0_4);
  assign port_state_out_1_0_5 = (port_state_in_1_0_5 ^ port_key_1_0_5);
  assign port_state_out_1_0_6 = (port_state_in_1_0_6 ^ port_key_1_0_6);
  assign port_state_out_1_0_7 = (port_state_in_1_0_7 ^ port_key_1_0_7);
  assign port_state_out_1_1_0 = (port_state_in_1_1_0 ^ port_key_1_1_0);
  assign port_state_out_1_1_1 = (port_state_in_1_1_1 ^ port_key_1_1_1);
  assign port_state_out_1_1_2 = (port_state_in_1_1_2 ^ port_key_1_1_2);
  assign port_state_out_1_1_3 = (port_state_in_1_1_3 ^ port_key_1_1_3);
  assign port_state_out_1_1_4 = (port_state_in_1_1_4 ^ port_key_1_1_4);
  assign port_state_out_1_1_5 = (port_state_in_1_1_5 ^ port_key_1_1_5);
  assign port_state_out_1_1_6 = (port_state_in_1_1_6 ^ port_key_1_1_6);
  assign port_state_out_1_1_7 = (port_state_in_1_1_7 ^ port_key_1_1_7);
  assign port_state_out_2_0_0 = (port_state_in_2_0_0 ^ port_key_2_0_0);
  assign port_state_out_2_0_1 = (port_state_in_2_0_1 ^ port_key_2_0_1);
  assign port_state_out_2_0_2 = (port_state_in_2_0_2 ^ port_key_2_0_2);
  assign port_state_out_2_0_3 = (port_state_in_2_0_3 ^ port_key_2_0_3);
  assign port_state_out_2_0_4 = (port_state_in_2_0_4 ^ port_key_2_0_4);
  assign port_state_out_2_0_5 = (port_state_in_2_0_5 ^ port_key_2_0_5);
  assign port_state_out_2_0_6 = (port_state_in_2_0_6 ^ port_key_2_0_6);
  assign port_state_out_2_0_7 = (port_state_in_2_0_7 ^ port_key_2_0_7);
  assign port_state_out_2_1_0 = (port_state_in_2_1_0 ^ port_key_2_1_0);
  assign port_state_out_2_1_1 = (port_state_in_2_1_1 ^ port_key_2_1_1);
  assign port_state_out_2_1_2 = (port_state_in_2_1_2 ^ port_key_2_1_2);
  assign port_state_out_2_1_3 = (port_state_in_2_1_3 ^ port_key_2_1_3);
  assign port_state_out_2_1_4 = (port_state_in_2_1_4 ^ port_key_2_1_4);
  assign port_state_out_2_1_5 = (port_state_in_2_1_5 ^ port_key_2_1_5);
  assign port_state_out_2_1_6 = (port_state_in_2_1_6 ^ port_key_2_1_6);
  assign port_state_out_2_1_7 = (port_state_in_2_1_7 ^ port_key_2_1_7);
  assign port_state_out_3_0_0 = (port_state_in_3_0_0 ^ port_key_3_0_0);
  assign port_state_out_3_0_1 = (port_state_in_3_0_1 ^ port_key_3_0_1);
  assign port_state_out_3_0_2 = (port_state_in_3_0_2 ^ port_key_3_0_2);
  assign port_state_out_3_0_3 = (port_state_in_3_0_3 ^ port_key_3_0_3);
  assign port_state_out_3_0_4 = (port_state_in_3_0_4 ^ port_key_3_0_4);
  assign port_state_out_3_0_5 = (port_state_in_3_0_5 ^ port_key_3_0_5);
  assign port_state_out_3_0_6 = (port_state_in_3_0_6 ^ port_key_3_0_6);
  assign port_state_out_3_0_7 = (port_state_in_3_0_7 ^ port_key_3_0_7);
  assign port_state_out_3_1_0 = (port_state_in_3_1_0 ^ port_key_3_1_0);
  assign port_state_out_3_1_1 = (port_state_in_3_1_1 ^ port_key_3_1_1);
  assign port_state_out_3_1_2 = (port_state_in_3_1_2 ^ port_key_3_1_2);
  assign port_state_out_3_1_3 = (port_state_in_3_1_3 ^ port_key_3_1_3);
  assign port_state_out_3_1_4 = (port_state_in_3_1_4 ^ port_key_3_1_4);
  assign port_state_out_3_1_5 = (port_state_in_3_1_5 ^ port_key_3_1_5);
  assign port_state_out_3_1_6 = (port_state_in_3_1_6 ^ port_key_3_1_6);
  assign port_state_out_3_1_7 = (port_state_in_3_1_7 ^ port_key_3_1_7);
  assign port_state_out_4_0_0 = (port_state_in_4_0_0 ^ port_key_4_0_0);
  assign port_state_out_4_0_1 = (port_state_in_4_0_1 ^ port_key_4_0_1);
  assign port_state_out_4_0_2 = (port_state_in_4_0_2 ^ port_key_4_0_2);
  assign port_state_out_4_0_3 = (port_state_in_4_0_3 ^ port_key_4_0_3);
  assign port_state_out_4_0_4 = (port_state_in_4_0_4 ^ port_key_4_0_4);
  assign port_state_out_4_0_5 = (port_state_in_4_0_5 ^ port_key_4_0_5);
  assign port_state_out_4_0_6 = (port_state_in_4_0_6 ^ port_key_4_0_6);
  assign port_state_out_4_0_7 = (port_state_in_4_0_7 ^ port_key_4_0_7);
  assign port_state_out_4_1_0 = (port_state_in_4_1_0 ^ port_key_4_1_0);
  assign port_state_out_4_1_1 = (port_state_in_4_1_1 ^ port_key_4_1_1);
  assign port_state_out_4_1_2 = (port_state_in_4_1_2 ^ port_key_4_1_2);
  assign port_state_out_4_1_3 = (port_state_in_4_1_3 ^ port_key_4_1_3);
  assign port_state_out_4_1_4 = (port_state_in_4_1_4 ^ port_key_4_1_4);
  assign port_state_out_4_1_5 = (port_state_in_4_1_5 ^ port_key_4_1_5);
  assign port_state_out_4_1_6 = (port_state_in_4_1_6 ^ port_key_4_1_6);
  assign port_state_out_4_1_7 = (port_state_in_4_1_7 ^ port_key_4_1_7);
  assign port_state_out_5_0_0 = (port_state_in_5_0_0 ^ port_key_5_0_0);
  assign port_state_out_5_0_1 = (port_state_in_5_0_1 ^ port_key_5_0_1);
  assign port_state_out_5_0_2 = (port_state_in_5_0_2 ^ port_key_5_0_2);
  assign port_state_out_5_0_3 = (port_state_in_5_0_3 ^ port_key_5_0_3);
  assign port_state_out_5_0_4 = (port_state_in_5_0_4 ^ port_key_5_0_4);
  assign port_state_out_5_0_5 = (port_state_in_5_0_5 ^ port_key_5_0_5);
  assign port_state_out_5_0_6 = (port_state_in_5_0_6 ^ port_key_5_0_6);
  assign port_state_out_5_0_7 = (port_state_in_5_0_7 ^ port_key_5_0_7);
  assign port_state_out_5_1_0 = (port_state_in_5_1_0 ^ port_key_5_1_0);
  assign port_state_out_5_1_1 = (port_state_in_5_1_1 ^ port_key_5_1_1);
  assign port_state_out_5_1_2 = (port_state_in_5_1_2 ^ port_key_5_1_2);
  assign port_state_out_5_1_3 = (port_state_in_5_1_3 ^ port_key_5_1_3);
  assign port_state_out_5_1_4 = (port_state_in_5_1_4 ^ port_key_5_1_4);
  assign port_state_out_5_1_5 = (port_state_in_5_1_5 ^ port_key_5_1_5);
  assign port_state_out_5_1_6 = (port_state_in_5_1_6 ^ port_key_5_1_6);
  assign port_state_out_5_1_7 = (port_state_in_5_1_7 ^ port_key_5_1_7);
  assign port_state_out_6_0_0 = (port_state_in_6_0_0 ^ port_key_6_0_0);
  assign port_state_out_6_0_1 = (port_state_in_6_0_1 ^ port_key_6_0_1);
  assign port_state_out_6_0_2 = (port_state_in_6_0_2 ^ port_key_6_0_2);
  assign port_state_out_6_0_3 = (port_state_in_6_0_3 ^ port_key_6_0_3);
  assign port_state_out_6_0_4 = (port_state_in_6_0_4 ^ port_key_6_0_4);
  assign port_state_out_6_0_5 = (port_state_in_6_0_5 ^ port_key_6_0_5);
  assign port_state_out_6_0_6 = (port_state_in_6_0_6 ^ port_key_6_0_6);
  assign port_state_out_6_0_7 = (port_state_in_6_0_7 ^ port_key_6_0_7);
  assign port_state_out_6_1_0 = (port_state_in_6_1_0 ^ port_key_6_1_0);
  assign port_state_out_6_1_1 = (port_state_in_6_1_1 ^ port_key_6_1_1);
  assign port_state_out_6_1_2 = (port_state_in_6_1_2 ^ port_key_6_1_2);
  assign port_state_out_6_1_3 = (port_state_in_6_1_3 ^ port_key_6_1_3);
  assign port_state_out_6_1_4 = (port_state_in_6_1_4 ^ port_key_6_1_4);
  assign port_state_out_6_1_5 = (port_state_in_6_1_5 ^ port_key_6_1_5);
  assign port_state_out_6_1_6 = (port_state_in_6_1_6 ^ port_key_6_1_6);
  assign port_state_out_6_1_7 = (port_state_in_6_1_7 ^ port_key_6_1_7);
  assign port_state_out_7_0_0 = (port_state_in_7_0_0 ^ port_key_7_0_0);
  assign port_state_out_7_0_1 = (port_state_in_7_0_1 ^ port_key_7_0_1);
  assign port_state_out_7_0_2 = (port_state_in_7_0_2 ^ port_key_7_0_2);
  assign port_state_out_7_0_3 = (port_state_in_7_0_3 ^ port_key_7_0_3);
  assign port_state_out_7_0_4 = (port_state_in_7_0_4 ^ port_key_7_0_4);
  assign port_state_out_7_0_5 = (port_state_in_7_0_5 ^ port_key_7_0_5);
  assign port_state_out_7_0_6 = (port_state_in_7_0_6 ^ port_key_7_0_6);
  assign port_state_out_7_0_7 = (port_state_in_7_0_7 ^ port_key_7_0_7);
  assign port_state_out_7_1_0 = (port_state_in_7_1_0 ^ port_key_7_1_0);
  assign port_state_out_7_1_1 = (port_state_in_7_1_1 ^ port_key_7_1_1);
  assign port_state_out_7_1_2 = (port_state_in_7_1_2 ^ port_key_7_1_2);
  assign port_state_out_7_1_3 = (port_state_in_7_1_3 ^ port_key_7_1_3);
  assign port_state_out_7_1_4 = (port_state_in_7_1_4 ^ port_key_7_1_4);
  assign port_state_out_7_1_5 = (port_state_in_7_1_5 ^ port_key_7_1_5);
  assign port_state_out_7_1_6 = (port_state_in_7_1_6 ^ port_key_7_1_6);
  assign port_state_out_7_1_7 = (port_state_in_7_1_7 ^ port_key_7_1_7);
  assign port_state_out_8_0_0 = (port_state_in_8_0_0 ^ port_key_8_0_0);
  assign port_state_out_8_0_1 = (port_state_in_8_0_1 ^ port_key_8_0_1);
  assign port_state_out_8_0_2 = (port_state_in_8_0_2 ^ port_key_8_0_2);
  assign port_state_out_8_0_3 = (port_state_in_8_0_3 ^ port_key_8_0_3);
  assign port_state_out_8_0_4 = (port_state_in_8_0_4 ^ port_key_8_0_4);
  assign port_state_out_8_0_5 = (port_state_in_8_0_5 ^ port_key_8_0_5);
  assign port_state_out_8_0_6 = (port_state_in_8_0_6 ^ port_key_8_0_6);
  assign port_state_out_8_0_7 = (port_state_in_8_0_7 ^ port_key_8_0_7);
  assign port_state_out_8_1_0 = (port_state_in_8_1_0 ^ port_key_8_1_0);
  assign port_state_out_8_1_1 = (port_state_in_8_1_1 ^ port_key_8_1_1);
  assign port_state_out_8_1_2 = (port_state_in_8_1_2 ^ port_key_8_1_2);
  assign port_state_out_8_1_3 = (port_state_in_8_1_3 ^ port_key_8_1_3);
  assign port_state_out_8_1_4 = (port_state_in_8_1_4 ^ port_key_8_1_4);
  assign port_state_out_8_1_5 = (port_state_in_8_1_5 ^ port_key_8_1_5);
  assign port_state_out_8_1_6 = (port_state_in_8_1_6 ^ port_key_8_1_6);
  assign port_state_out_8_1_7 = (port_state_in_8_1_7 ^ port_key_8_1_7);
  assign port_state_out_9_0_0 = (port_state_in_9_0_0 ^ port_key_9_0_0);
  assign port_state_out_9_0_1 = (port_state_in_9_0_1 ^ port_key_9_0_1);
  assign port_state_out_9_0_2 = (port_state_in_9_0_2 ^ port_key_9_0_2);
  assign port_state_out_9_0_3 = (port_state_in_9_0_3 ^ port_key_9_0_3);
  assign port_state_out_9_0_4 = (port_state_in_9_0_4 ^ port_key_9_0_4);
  assign port_state_out_9_0_5 = (port_state_in_9_0_5 ^ port_key_9_0_5);
  assign port_state_out_9_0_6 = (port_state_in_9_0_6 ^ port_key_9_0_6);
  assign port_state_out_9_0_7 = (port_state_in_9_0_7 ^ port_key_9_0_7);
  assign port_state_out_9_1_0 = (port_state_in_9_1_0 ^ port_key_9_1_0);
  assign port_state_out_9_1_1 = (port_state_in_9_1_1 ^ port_key_9_1_1);
  assign port_state_out_9_1_2 = (port_state_in_9_1_2 ^ port_key_9_1_2);
  assign port_state_out_9_1_3 = (port_state_in_9_1_3 ^ port_key_9_1_3);
  assign port_state_out_9_1_4 = (port_state_in_9_1_4 ^ port_key_9_1_4);
  assign port_state_out_9_1_5 = (port_state_in_9_1_5 ^ port_key_9_1_5);
  assign port_state_out_9_1_6 = (port_state_in_9_1_6 ^ port_key_9_1_6);
  assign port_state_out_9_1_7 = (port_state_in_9_1_7 ^ port_key_9_1_7);
  assign port_state_out_10_0_0 = (port_state_in_10_0_0 ^ port_key_10_0_0);
  assign port_state_out_10_0_1 = (port_state_in_10_0_1 ^ port_key_10_0_1);
  assign port_state_out_10_0_2 = (port_state_in_10_0_2 ^ port_key_10_0_2);
  assign port_state_out_10_0_3 = (port_state_in_10_0_3 ^ port_key_10_0_3);
  assign port_state_out_10_0_4 = (port_state_in_10_0_4 ^ port_key_10_0_4);
  assign port_state_out_10_0_5 = (port_state_in_10_0_5 ^ port_key_10_0_5);
  assign port_state_out_10_0_6 = (port_state_in_10_0_6 ^ port_key_10_0_6);
  assign port_state_out_10_0_7 = (port_state_in_10_0_7 ^ port_key_10_0_7);
  assign port_state_out_10_1_0 = (port_state_in_10_1_0 ^ port_key_10_1_0);
  assign port_state_out_10_1_1 = (port_state_in_10_1_1 ^ port_key_10_1_1);
  assign port_state_out_10_1_2 = (port_state_in_10_1_2 ^ port_key_10_1_2);
  assign port_state_out_10_1_3 = (port_state_in_10_1_3 ^ port_key_10_1_3);
  assign port_state_out_10_1_4 = (port_state_in_10_1_4 ^ port_key_10_1_4);
  assign port_state_out_10_1_5 = (port_state_in_10_1_5 ^ port_key_10_1_5);
  assign port_state_out_10_1_6 = (port_state_in_10_1_6 ^ port_key_10_1_6);
  assign port_state_out_10_1_7 = (port_state_in_10_1_7 ^ port_key_10_1_7);
  assign port_state_out_11_0_0 = (port_state_in_11_0_0 ^ port_key_11_0_0);
  assign port_state_out_11_0_1 = (port_state_in_11_0_1 ^ port_key_11_0_1);
  assign port_state_out_11_0_2 = (port_state_in_11_0_2 ^ port_key_11_0_2);
  assign port_state_out_11_0_3 = (port_state_in_11_0_3 ^ port_key_11_0_3);
  assign port_state_out_11_0_4 = (port_state_in_11_0_4 ^ port_key_11_0_4);
  assign port_state_out_11_0_5 = (port_state_in_11_0_5 ^ port_key_11_0_5);
  assign port_state_out_11_0_6 = (port_state_in_11_0_6 ^ port_key_11_0_6);
  assign port_state_out_11_0_7 = (port_state_in_11_0_7 ^ port_key_11_0_7);
  assign port_state_out_11_1_0 = (port_state_in_11_1_0 ^ port_key_11_1_0);
  assign port_state_out_11_1_1 = (port_state_in_11_1_1 ^ port_key_11_1_1);
  assign port_state_out_11_1_2 = (port_state_in_11_1_2 ^ port_key_11_1_2);
  assign port_state_out_11_1_3 = (port_state_in_11_1_3 ^ port_key_11_1_3);
  assign port_state_out_11_1_4 = (port_state_in_11_1_4 ^ port_key_11_1_4);
  assign port_state_out_11_1_5 = (port_state_in_11_1_5 ^ port_key_11_1_5);
  assign port_state_out_11_1_6 = (port_state_in_11_1_6 ^ port_key_11_1_6);
  assign port_state_out_11_1_7 = (port_state_in_11_1_7 ^ port_key_11_1_7);
  assign port_state_out_12_0_0 = (port_state_in_12_0_0 ^ port_key_12_0_0);
  assign port_state_out_12_0_1 = (port_state_in_12_0_1 ^ port_key_12_0_1);
  assign port_state_out_12_0_2 = (port_state_in_12_0_2 ^ port_key_12_0_2);
  assign port_state_out_12_0_3 = (port_state_in_12_0_3 ^ port_key_12_0_3);
  assign port_state_out_12_0_4 = (port_state_in_12_0_4 ^ port_key_12_0_4);
  assign port_state_out_12_0_5 = (port_state_in_12_0_5 ^ port_key_12_0_5);
  assign port_state_out_12_0_6 = (port_state_in_12_0_6 ^ port_key_12_0_6);
  assign port_state_out_12_0_7 = (port_state_in_12_0_7 ^ port_key_12_0_7);
  assign port_state_out_12_1_0 = (port_state_in_12_1_0 ^ port_key_12_1_0);
  assign port_state_out_12_1_1 = (port_state_in_12_1_1 ^ port_key_12_1_1);
  assign port_state_out_12_1_2 = (port_state_in_12_1_2 ^ port_key_12_1_2);
  assign port_state_out_12_1_3 = (port_state_in_12_1_3 ^ port_key_12_1_3);
  assign port_state_out_12_1_4 = (port_state_in_12_1_4 ^ port_key_12_1_4);
  assign port_state_out_12_1_5 = (port_state_in_12_1_5 ^ port_key_12_1_5);
  assign port_state_out_12_1_6 = (port_state_in_12_1_6 ^ port_key_12_1_6);
  assign port_state_out_12_1_7 = (port_state_in_12_1_7 ^ port_key_12_1_7);
  assign port_state_out_13_0_0 = (port_state_in_13_0_0 ^ port_key_13_0_0);
  assign port_state_out_13_0_1 = (port_state_in_13_0_1 ^ port_key_13_0_1);
  assign port_state_out_13_0_2 = (port_state_in_13_0_2 ^ port_key_13_0_2);
  assign port_state_out_13_0_3 = (port_state_in_13_0_3 ^ port_key_13_0_3);
  assign port_state_out_13_0_4 = (port_state_in_13_0_4 ^ port_key_13_0_4);
  assign port_state_out_13_0_5 = (port_state_in_13_0_5 ^ port_key_13_0_5);
  assign port_state_out_13_0_6 = (port_state_in_13_0_6 ^ port_key_13_0_6);
  assign port_state_out_13_0_7 = (port_state_in_13_0_7 ^ port_key_13_0_7);
  assign port_state_out_13_1_0 = (port_state_in_13_1_0 ^ port_key_13_1_0);
  assign port_state_out_13_1_1 = (port_state_in_13_1_1 ^ port_key_13_1_1);
  assign port_state_out_13_1_2 = (port_state_in_13_1_2 ^ port_key_13_1_2);
  assign port_state_out_13_1_3 = (port_state_in_13_1_3 ^ port_key_13_1_3);
  assign port_state_out_13_1_4 = (port_state_in_13_1_4 ^ port_key_13_1_4);
  assign port_state_out_13_1_5 = (port_state_in_13_1_5 ^ port_key_13_1_5);
  assign port_state_out_13_1_6 = (port_state_in_13_1_6 ^ port_key_13_1_6);
  assign port_state_out_13_1_7 = (port_state_in_13_1_7 ^ port_key_13_1_7);
  assign port_state_out_14_0_0 = (port_state_in_14_0_0 ^ port_key_14_0_0);
  assign port_state_out_14_0_1 = (port_state_in_14_0_1 ^ port_key_14_0_1);
  assign port_state_out_14_0_2 = (port_state_in_14_0_2 ^ port_key_14_0_2);
  assign port_state_out_14_0_3 = (port_state_in_14_0_3 ^ port_key_14_0_3);
  assign port_state_out_14_0_4 = (port_state_in_14_0_4 ^ port_key_14_0_4);
  assign port_state_out_14_0_5 = (port_state_in_14_0_5 ^ port_key_14_0_5);
  assign port_state_out_14_0_6 = (port_state_in_14_0_6 ^ port_key_14_0_6);
  assign port_state_out_14_0_7 = (port_state_in_14_0_7 ^ port_key_14_0_7);
  assign port_state_out_14_1_0 = (port_state_in_14_1_0 ^ port_key_14_1_0);
  assign port_state_out_14_1_1 = (port_state_in_14_1_1 ^ port_key_14_1_1);
  assign port_state_out_14_1_2 = (port_state_in_14_1_2 ^ port_key_14_1_2);
  assign port_state_out_14_1_3 = (port_state_in_14_1_3 ^ port_key_14_1_3);
  assign port_state_out_14_1_4 = (port_state_in_14_1_4 ^ port_key_14_1_4);
  assign port_state_out_14_1_5 = (port_state_in_14_1_5 ^ port_key_14_1_5);
  assign port_state_out_14_1_6 = (port_state_in_14_1_6 ^ port_key_14_1_6);
  assign port_state_out_14_1_7 = (port_state_in_14_1_7 ^ port_key_14_1_7);
  assign port_state_out_15_0_0 = (port_state_in_15_0_0 ^ port_key_15_0_0);
  assign port_state_out_15_0_1 = (port_state_in_15_0_1 ^ port_key_15_0_1);
  assign port_state_out_15_0_2 = (port_state_in_15_0_2 ^ port_key_15_0_2);
  assign port_state_out_15_0_3 = (port_state_in_15_0_3 ^ port_key_15_0_3);
  assign port_state_out_15_0_4 = (port_state_in_15_0_4 ^ port_key_15_0_4);
  assign port_state_out_15_0_5 = (port_state_in_15_0_5 ^ port_key_15_0_5);
  assign port_state_out_15_0_6 = (port_state_in_15_0_6 ^ port_key_15_0_6);
  assign port_state_out_15_0_7 = (port_state_in_15_0_7 ^ port_key_15_0_7);
  assign port_state_out_15_1_0 = (port_state_in_15_1_0 ^ port_key_15_1_0);
  assign port_state_out_15_1_1 = (port_state_in_15_1_1 ^ port_key_15_1_1);
  assign port_state_out_15_1_2 = (port_state_in_15_1_2 ^ port_key_15_1_2);
  assign port_state_out_15_1_3 = (port_state_in_15_1_3 ^ port_key_15_1_3);
  assign port_state_out_15_1_4 = (port_state_in_15_1_4 ^ port_key_15_1_4);
  assign port_state_out_15_1_5 = (port_state_in_15_1_5 ^ port_key_15_1_5);
  assign port_state_out_15_1_6 = (port_state_in_15_1_6 ^ port_key_15_1_6);
  assign port_state_out_15_1_7 = (port_state_in_15_1_7 ^ port_key_15_1_7);

endmodule

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

module Mul3 (
  input      [0:0]    port_byte_in_0,
  input      [0:0]    port_byte_in_1,
  input      [0:0]    port_byte_in_2,
  input      [0:0]    port_byte_in_3,
  input      [0:0]    port_byte_in_4,
  input      [0:0]    port_byte_in_5,
  input      [0:0]    port_byte_in_6,
  input      [0:0]    port_byte_in_7,
  output     [0:0]    port_byte_out_0,
  output     [0:0]    port_byte_out_1,
  output     [0:0]    port_byte_out_2,
  output     [0:0]    port_byte_out_3,
  output     [0:0]    port_byte_out_4,
  output     [0:0]    port_byte_out_5,
  output     [0:0]    port_byte_out_6,
  output     [0:0]    port_byte_out_7
);


  assign port_byte_out_7 = (port_byte_in_7 ^ port_byte_in_6);
  assign port_byte_out_6 = (port_byte_in_6 ^ port_byte_in_5);
  assign port_byte_out_5 = (port_byte_in_5 ^ port_byte_in_4);
  assign port_byte_out_4 = ((port_byte_in_7 ^ port_byte_in_4) ^ port_byte_in_3);
  assign port_byte_out_3 = ((port_byte_in_7 ^ port_byte_in_3) ^ port_byte_in_2);
  assign port_byte_out_2 = (port_byte_in_2 ^ port_byte_in_1);
  assign port_byte_out_1 = ((port_byte_in_7 ^ port_byte_in_1) ^ port_byte_in_0);
  assign port_byte_out_0 = (port_byte_in_7 ^ port_byte_in_0);

endmodule

module Mul2 (
  input      [0:0]    port_byte_in_0,
  input      [0:0]    port_byte_in_1,
  input      [0:0]    port_byte_in_2,
  input      [0:0]    port_byte_in_3,
  input      [0:0]    port_byte_in_4,
  input      [0:0]    port_byte_in_5,
  input      [0:0]    port_byte_in_6,
  input      [0:0]    port_byte_in_7,
  output     [0:0]    port_byte_out_0,
  output     [0:0]    port_byte_out_1,
  output     [0:0]    port_byte_out_2,
  output     [0:0]    port_byte_out_3,
  output     [0:0]    port_byte_out_4,
  output     [0:0]    port_byte_out_5,
  output     [0:0]    port_byte_out_6,
  output     [0:0]    port_byte_out_7
);


  assign port_byte_out_7 = port_byte_in_6;
  assign port_byte_out_6 = port_byte_in_5;
  assign port_byte_out_5 = port_byte_in_4;
  assign port_byte_out_4 = (port_byte_in_7 ^ port_byte_in_3);
  assign port_byte_out_3 = (port_byte_in_7 ^ port_byte_in_2);
  assign port_byte_out_2 = port_byte_in_1;
  assign port_byte_out_1 = (port_byte_in_7 ^ port_byte_in_0);
  assign port_byte_out_0 = port_byte_in_7;

endmodule

//CMS_stage6 replaced by CMS_stage6

//CMS_stage5 replaced by CMS_stage5

//CMS_stage4 replaced by CMS_stage4

//CMS_stage3 replaced by CMS_stage3

//CMS_stage2 replaced by CMS_stage2

//CMS_stage1 replaced by CMS_stage1

//CMS_stage6 replaced by CMS_stage6

//CMS_stage5 replaced by CMS_stage5

//CMS_stage4 replaced by CMS_stage4

//CMS_stage3 replaced by CMS_stage3

//CMS_stage2 replaced by CMS_stage2

//CMS_stage1 replaced by CMS_stage1

//CMS_stage6 replaced by CMS_stage6

//CMS_stage5 replaced by CMS_stage5

//CMS_stage4 replaced by CMS_stage4

//CMS_stage3 replaced by CMS_stage3

//CMS_stage2 replaced by CMS_stage2

//CMS_stage1 replaced by CMS_stage1

//CMS_stage6 replaced by CMS_stage6

//CMS_stage5 replaced by CMS_stage5

//CMS_stage4 replaced by CMS_stage4

//CMS_stage3 replaced by CMS_stage3

//CMS_stage2 replaced by CMS_stage2

//CMS_stage1 replaced by CMS_stage1

//CMS_stage6 replaced by CMS_stage6

//CMS_stage5 replaced by CMS_stage5

//CMS_stage4 replaced by CMS_stage4

//CMS_stage3 replaced by CMS_stage3

//CMS_stage2 replaced by CMS_stage2

//CMS_stage1 replaced by CMS_stage1

//CMS_stage6 replaced by CMS_stage6

//CMS_stage5 replaced by CMS_stage5

//CMS_stage4 replaced by CMS_stage4

//CMS_stage3 replaced by CMS_stage3

//CMS_stage2 replaced by CMS_stage2

//CMS_stage1 replaced by CMS_stage1

//CMS_stage6 replaced by CMS_stage6

//CMS_stage5 replaced by CMS_stage5

//CMS_stage4 replaced by CMS_stage4

//CMS_stage3 replaced by CMS_stage3

//CMS_stage2 replaced by CMS_stage2

//CMS_stage1 replaced by CMS_stage1

//CMS_stage6 replaced by CMS_stage6

//CMS_stage5 replaced by CMS_stage5

//CMS_stage4 replaced by CMS_stage4

//CMS_stage3 replaced by CMS_stage3

//CMS_stage2 replaced by CMS_stage2

//CMS_stage1 replaced by CMS_stage1

//CMS_stage6 replaced by CMS_stage6

//CMS_stage5 replaced by CMS_stage5

//CMS_stage4 replaced by CMS_stage4

//CMS_stage3 replaced by CMS_stage3

//CMS_stage2 replaced by CMS_stage2

//CMS_stage1 replaced by CMS_stage1

//CMS_stage6 replaced by CMS_stage6

//CMS_stage5 replaced by CMS_stage5

//CMS_stage4 replaced by CMS_stage4

//CMS_stage3 replaced by CMS_stage3

//CMS_stage2 replaced by CMS_stage2

//CMS_stage1 replaced by CMS_stage1

//CMS_stage6 replaced by CMS_stage6

//CMS_stage5 replaced by CMS_stage5

//CMS_stage4 replaced by CMS_stage4

//CMS_stage3 replaced by CMS_stage3

//CMS_stage2 replaced by CMS_stage2

//CMS_stage1 replaced by CMS_stage1

//CMS_stage6 replaced by CMS_stage6

//CMS_stage5 replaced by CMS_stage5

//CMS_stage4 replaced by CMS_stage4

//CMS_stage3 replaced by CMS_stage3

//CMS_stage2 replaced by CMS_stage2

//CMS_stage1 replaced by CMS_stage1

//CMS_stage6 replaced by CMS_stage6

//CMS_stage5 replaced by CMS_stage5

//CMS_stage4 replaced by CMS_stage4

//CMS_stage3 replaced by CMS_stage3

//CMS_stage2 replaced by CMS_stage2

//CMS_stage1 replaced by CMS_stage1

//CMS_stage6 replaced by CMS_stage6

//CMS_stage5 replaced by CMS_stage5

//CMS_stage4 replaced by CMS_stage4

//CMS_stage3 replaced by CMS_stage3

//CMS_stage2 replaced by CMS_stage2

//CMS_stage1 replaced by CMS_stage1

//CMS_stage6 replaced by CMS_stage6

//CMS_stage5 replaced by CMS_stage5

//CMS_stage4 replaced by CMS_stage4

//CMS_stage3 replaced by CMS_stage3

//CMS_stage2 replaced by CMS_stage2

//CMS_stage1 replaced by CMS_stage1

module CMS_stage6 (
  input      [0:0]    port_i_0_0,
  input      [0:0]    port_i_0_1,
  input      [0:0]    port_i_0_2,
  input      [0:0]    port_i_0_3,
  input      [0:0]    port_i_0_4,
  input      [0:0]    port_i_0_5,
  input      [0:0]    port_i_0_6,
  input      [0:0]    port_i_0_7,
  input      [0:0]    port_i_1_0,
  input      [0:0]    port_i_1_1,
  input      [0:0]    port_i_1_2,
  input      [0:0]    port_i_1_3,
  input      [0:0]    port_i_1_4,
  input      [0:0]    port_i_1_5,
  input      [0:0]    port_i_1_6,
  input      [0:0]    port_i_1_7,
  output     [0:0]    port_o_0_0,
  output     [0:0]    port_o_0_1,
  output     [0:0]    port_o_0_2,
  output     [0:0]    port_o_0_3,
  output     [0:0]    port_o_0_4,
  output     [0:0]    port_o_0_5,
  output     [0:0]    port_o_0_6,
  output     [0:0]    port_o_0_7,
  output     [0:0]    port_o_1_0,
  output     [0:0]    port_o_1_1,
  output     [0:0]    port_o_1_2,
  output     [0:0]    port_o_1_3,
  output     [0:0]    port_o_1_4,
  output     [0:0]    port_o_1_5,
  output     [0:0]    port_o_1_6,
  output     [0:0]    port_o_1_7
);

  wire       [0:0]    tx1_0;
  wire       [0:0]    tx2_0;
  wire       [0:0]    tx3_0;
  wire       [0:0]    tx4_0;
  wire       [0:0]    tx5_0;
  wire       [0:0]    tx6_0;
  wire       [0:0]    tx7_0;
  wire       [0:0]    tx8_0;
  wire       [0:0]    tx9_0;
  wire       [0:0]    tx10_0;
  wire       [0:0]    tx1_1;
  wire       [0:0]    tx2_1;
  wire       [0:0]    tx3_1;
  wire       [0:0]    tx4_1;
  wire       [0:0]    tx5_1;
  wire       [0:0]    tx6_1;
  wire       [0:0]    tx7_1;
  wire       [0:0]    tx8_1;
  wire       [0:0]    tx9_1;
  wire       [0:0]    tx10_1;

  assign tx1_0 = (port_i_0_7 ^ port_i_0_3);
  assign tx2_0 = (port_i_0_6 ^ port_i_0_4);
  assign tx3_0 = (port_i_0_6 ^ port_i_0_0);
  assign tx4_0 = (~ (port_i_0_5 ^ port_i_0_3));
  assign tx5_0 = (~ (port_i_0_5 ^ tx1_0));
  assign tx6_0 = (~ (port_i_0_5 ^ port_i_0_1));
  assign tx7_0 = (~ (port_i_0_4 ^ tx6_0));
  assign tx8_0 = (port_i_0_2 ^ tx4_0);
  assign tx9_0 = (port_i_0_1 ^ tx2_0);
  assign tx10_0 = (tx3_0 ^ tx5_0);
  assign port_o_0_7 = (~ tx4_0);
  assign port_o_0_6 = (~ tx1_0);
  assign port_o_0_5 = (~ tx3_0);
  assign port_o_0_4 = (~ tx5_0);
  assign port_o_0_3 = (~ (tx2_0 ^ tx5_0));
  assign port_o_0_2 = (~ (tx3_0 ^ tx8_0));
  assign port_o_0_1 = (~ tx7_0);
  assign port_o_0_0 = (~ tx9_0);
  assign tx1_1 = (port_i_1_7 ^ port_i_1_3);
  assign tx2_1 = (port_i_1_6 ^ port_i_1_4);
  assign tx3_1 = (port_i_1_6 ^ port_i_1_0);
  assign tx4_1 = (port_i_1_5 ^ port_i_1_3);
  assign tx5_1 = (port_i_1_5 ^ tx1_1);
  assign tx6_1 = (port_i_1_5 ^ port_i_1_1);
  assign tx7_1 = (port_i_1_4 ^ tx6_1);
  assign tx8_1 = (port_i_1_2 ^ tx4_1);
  assign tx9_1 = (port_i_1_1 ^ tx2_1);
  assign tx10_1 = (tx3_1 ^ tx5_1);
  assign port_o_1_7 = tx4_1;
  assign port_o_1_6 = tx1_1;
  assign port_o_1_5 = tx3_1;
  assign port_o_1_4 = tx5_1;
  assign port_o_1_3 = (tx2_1 ^ tx5_1);
  assign port_o_1_2 = (tx3_1 ^ tx8_1);
  assign port_o_1_1 = tx7_1;
  assign port_o_1_0 = tx9_1;

endmodule

module CMS_stage5 (
  input      [0:0]    port_a_0_0,
  input      [0:0]    port_a_0_1,
  input      [0:0]    port_a_0_2,
  input      [0:0]    port_a_0_3,
  input      [0:0]    port_a_1_0,
  input      [0:0]    port_a_1_1,
  input      [0:0]    port_a_1_2,
  input      [0:0]    port_a_1_3,
  input      [0:0]    port_b_0_0,
  input      [0:0]    port_b_0_1,
  input      [0:0]    port_b_0_2,
  input      [0:0]    port_b_0_3,
  input      [0:0]    port_b_1_0,
  input      [0:0]    port_b_1_1,
  input      [0:0]    port_b_1_2,
  input      [0:0]    port_b_1_3,
  input      [0:0]    port_c_0_0,
  input      [0:0]    port_c_0_1,
  input      [0:0]    port_c_0_2,
  input      [0:0]    port_c_0_3,
  input      [0:0]    port_c_1_0,
  input      [0:0]    port_c_1_1,
  input      [0:0]    port_c_1_2,
  input      [0:0]    port_c_1_3,
  input               port_r_0_0,
  input               port_r_0_1,
  input               port_r_0_2,
  input               port_r_0_3,
  input               port_r_0_4,
  input               port_r_0_5,
  input               port_r_0_6,
  input               port_r_0_7,
  input               port_r_1_0,
  input               port_r_1_1,
  input               port_r_1_2,
  input               port_r_1_3,
  input               port_r_1_4,
  input               port_r_1_5,
  input               port_r_1_6,
  input               port_r_1_7,
  input               port_r_2_0,
  input               port_r_2_1,
  input               port_r_2_2,
  input               port_r_2_3,
  input               port_r_2_4,
  input               port_r_2_5,
  input               port_r_2_6,
  input               port_r_2_7,
  output     [0:0]    port_y_0_0,
  output     [0:0]    port_y_0_1,
  output     [0:0]    port_y_0_2,
  output     [0:0]    port_y_0_3,
  output     [0:0]    port_y_0_4,
  output     [0:0]    port_y_0_5,
  output     [0:0]    port_y_0_6,
  output     [0:0]    port_y_0_7,
  output     [0:0]    port_y_1_0,
  output     [0:0]    port_y_1_1,
  output     [0:0]    port_y_1_2,
  output     [0:0]    port_y_1_3,
  output     [0:0]    port_y_1_4,
  output     [0:0]    port_y_1_5,
  output     [0:0]    port_y_1_6,
  output     [0:0]    port_y_1_7,
  output     [0:0]    port_y_2_0,
  output     [0:0]    port_y_2_1,
  output     [0:0]    port_y_2_2,
  output     [0:0]    port_y_2_3,
  output     [0:0]    port_y_2_4,
  output     [0:0]    port_y_2_5,
  output     [0:0]    port_y_2_6,
  output     [0:0]    port_y_2_7,
  output     [0:0]    port_y_3_0,
  output     [0:0]    port_y_3_1,
  output     [0:0]    port_y_3_2,
  output     [0:0]    port_y_3_3,
  output     [0:0]    port_y_3_4,
  output     [0:0]    port_y_3_5,
  output     [0:0]    port_y_3_6,
  output     [0:0]    port_y_3_7,
  input               clk,
  input               reset
);

  wire       [0:0]    gF_MULS_4_192_port_o_0;
  wire       [0:0]    gF_MULS_4_192_port_o_1;
  wire       [0:0]    gF_MULS_4_192_port_o_2;
  wire       [0:0]    gF_MULS_4_192_port_o_3;
  wire       [0:0]    gF_MULS_4_193_port_o_0;
  wire       [0:0]    gF_MULS_4_193_port_o_1;
  wire       [0:0]    gF_MULS_4_193_port_o_2;
  wire       [0:0]    gF_MULS_4_193_port_o_3;
  wire       [0:0]    gF_MULS_4_194_port_o_0;
  wire       [0:0]    gF_MULS_4_194_port_o_1;
  wire       [0:0]    gF_MULS_4_194_port_o_2;
  wire       [0:0]    gF_MULS_4_194_port_o_3;
  wire       [0:0]    gF_MULS_4_195_port_o_0;
  wire       [0:0]    gF_MULS_4_195_port_o_1;
  wire       [0:0]    gF_MULS_4_195_port_o_2;
  wire       [0:0]    gF_MULS_4_195_port_o_3;
  wire       [0:0]    gF_MULS_4_196_port_o_0;
  wire       [0:0]    gF_MULS_4_196_port_o_1;
  wire       [0:0]    gF_MULS_4_196_port_o_2;
  wire       [0:0]    gF_MULS_4_196_port_o_3;
  wire       [0:0]    gF_MULS_4_197_port_o_0;
  wire       [0:0]    gF_MULS_4_197_port_o_1;
  wire       [0:0]    gF_MULS_4_197_port_o_2;
  wire       [0:0]    gF_MULS_4_197_port_o_3;
  wire       [0:0]    gF_MULS_4_198_port_o_0;
  wire       [0:0]    gF_MULS_4_198_port_o_1;
  wire       [0:0]    gF_MULS_4_198_port_o_2;
  wire       [0:0]    gF_MULS_4_198_port_o_3;
  wire       [0:0]    gF_MULS_4_199_port_o_0;
  wire       [0:0]    gF_MULS_4_199_port_o_1;
  wire       [0:0]    gF_MULS_4_199_port_o_2;
  wire       [0:0]    gF_MULS_4_199_port_o_3;
  reg        [0:0]    outReg_0_0;
  reg        [0:0]    outReg_0_1;
  reg        [0:0]    outReg_0_2;
  reg        [0:0]    outReg_0_3;
  reg        [0:0]    outReg_0_4;
  reg        [0:0]    outReg_0_5;
  reg        [0:0]    outReg_0_6;
  reg        [0:0]    outReg_0_7;
  reg        [0:0]    outReg_1_0;
  reg        [0:0]    outReg_1_1;
  reg        [0:0]    outReg_1_2;
  reg        [0:0]    outReg_1_3;
  reg        [0:0]    outReg_1_4;
  reg        [0:0]    outReg_1_5;
  reg        [0:0]    outReg_1_6;
  reg        [0:0]    outReg_1_7;
  reg        [0:0]    outReg_2_0;
  reg        [0:0]    outReg_2_1;
  reg        [0:0]    outReg_2_2;
  reg        [0:0]    outReg_2_3;
  reg        [0:0]    outReg_2_4;
  reg        [0:0]    outReg_2_5;
  reg        [0:0]    outReg_2_6;
  reg        [0:0]    outReg_2_7;
  reg        [0:0]    outReg_3_0;
  reg        [0:0]    outReg_3_1;
  reg        [0:0]    outReg_3_2;
  reg        [0:0]    outReg_3_3;
  reg        [0:0]    outReg_3_4;
  reg        [0:0]    outReg_3_5;
  reg        [0:0]    outReg_3_6;
  reg        [0:0]    outReg_3_7;
  wire       [0:0]    outVal_0_0;
  wire       [0:0]    outVal_0_1;
  wire       [0:0]    outVal_0_2;
  wire       [0:0]    outVal_0_3;
  wire       [0:0]    outVal_0_4;
  wire       [0:0]    outVal_0_5;
  wire       [0:0]    outVal_0_6;
  wire       [0:0]    outVal_0_7;
  wire       [0:0]    outVal_1_0;
  wire       [0:0]    outVal_1_1;
  wire       [0:0]    outVal_1_2;
  wire       [0:0]    outVal_1_3;
  wire       [0:0]    outVal_1_4;
  wire       [0:0]    outVal_1_5;
  wire       [0:0]    outVal_1_6;
  wire       [0:0]    outVal_1_7;
  wire       [0:0]    outVal_2_0;
  wire       [0:0]    outVal_2_1;
  wire       [0:0]    outVal_2_2;
  wire       [0:0]    outVal_2_3;
  wire       [0:0]    outVal_2_4;
  wire       [0:0]    outVal_2_5;
  wire       [0:0]    outVal_2_6;
  wire       [0:0]    outVal_2_7;
  wire       [0:0]    outVal_3_0;
  wire       [0:0]    outVal_3_1;
  wire       [0:0]    outVal_3_2;
  wire       [0:0]    outVal_3_3;
  wire       [0:0]    outVal_3_4;
  wire       [0:0]    outVal_3_5;
  wire       [0:0]    outVal_3_6;
  wire       [0:0]    outVal_3_7;
  wire       [0:0]    refVal_0_0;
  wire       [0:0]    refVal_0_1;
  wire       [0:0]    refVal_0_2;
  wire       [0:0]    refVal_0_3;
  wire       [0:0]    refVal_0_4;
  wire       [0:0]    refVal_0_5;
  wire       [0:0]    refVal_0_6;
  wire       [0:0]    refVal_0_7;
  wire       [0:0]    refVal_1_0;
  wire       [0:0]    refVal_1_1;
  wire       [0:0]    refVal_1_2;
  wire       [0:0]    refVal_1_3;
  wire       [0:0]    refVal_1_4;
  wire       [0:0]    refVal_1_5;
  wire       [0:0]    refVal_1_6;
  wire       [0:0]    refVal_1_7;
  wire       [0:0]    refVal_2_0;
  wire       [0:0]    refVal_2_1;
  wire       [0:0]    refVal_2_2;
  wire       [0:0]    refVal_2_3;
  wire       [0:0]    refVal_2_4;
  wire       [0:0]    refVal_2_5;
  wire       [0:0]    refVal_2_6;
  wire       [0:0]    refVal_2_7;
  wire       [0:0]    refVal_3_0;
  wire       [0:0]    refVal_3_1;
  wire       [0:0]    refVal_3_2;
  wire       [0:0]    refVal_3_3;
  wire       [0:0]    refVal_3_4;
  wire       [0:0]    refVal_3_5;
  wire       [0:0]    refVal_3_6;
  wire       [0:0]    refVal_3_7;
  wire       [0:0]    sax_0_0;
  wire       [0:0]    sax_0_1;
  wire       [0:0]    sax_1_0;
  wire       [0:0]    sax_1_1;
  wire       [0:0]    sbx_0_0;
  wire       [0:0]    sbx_0_1;
  wire       [0:0]    sbx_1_0;
  wire       [0:0]    sbx_1_1;
  wire       [0:0]    scx_0_0;
  wire       [0:0]    scx_0_1;
  wire       [0:0]    scx_1_0;
  wire       [0:0]    scx_1_1;
  wire       [0:0]    al_0;
  wire       [0:0]    al_1;
  wire       [0:0]    ah_0;
  wire       [0:0]    ah_1;
  wire       [0:0]    aa_0;
  wire       [0:0]    aa_1;
  wire       [0:0]    bl_0;
  wire       [0:0]    bl_1;
  wire       [0:0]    bh_0;
  wire       [0:0]    bh_1;
  wire       [0:0]    bb_0;
  wire       [0:0]    bb_1;
  wire       [0:0]    cl_0;
  wire       [0:0]    cl_1;
  wire       [0:0]    ch_0;
  wire       [0:0]    ch_1;
  wire       [0:0]    cc_0;
  wire       [0:0]    cc_1;

  GF_MULS_4 gF_MULS_4_192 (
    .port_A_0   (port_b_0_0            ), //i
    .port_A_1   (port_b_0_1            ), //i
    .port_A_2   (port_b_0_2            ), //i
    .port_A_3   (port_b_0_3            ), //i
    .port_a_0_1 (sbx_0_0               ), //i
    .port_a_1_1 (sbx_0_1               ), //i
    .port_Al    (bl_0                  ), //i
    .port_Ah    (bh_0                  ), //i
    .port_aa    (bb_0                  ), //i
    .port_B_0   (port_a_0_0            ), //i
    .port_B_1   (port_a_0_1            ), //i
    .port_B_2   (port_a_0_2            ), //i
    .port_B_3   (port_a_0_3            ), //i
    .port_b_0_1 (sax_0_0               ), //i
    .port_b_1_1 (sax_0_1               ), //i
    .port_Bl    (al_0                  ), //i
    .port_Bh    (ah_0                  ), //i
    .port_bb    (aa_0                  ), //i
    .port_o_0   (gF_MULS_4_192_port_o_0), //o
    .port_o_1   (gF_MULS_4_192_port_o_1), //o
    .port_o_2   (gF_MULS_4_192_port_o_2), //o
    .port_o_3   (gF_MULS_4_192_port_o_3)  //o
  );
  GF_MULS_4 gF_MULS_4_193 (
    .port_A_0   (port_b_0_0            ), //i
    .port_A_1   (port_b_0_1            ), //i
    .port_A_2   (port_b_0_2            ), //i
    .port_A_3   (port_b_0_3            ), //i
    .port_a_0_1 (sbx_0_0               ), //i
    .port_a_1_1 (sbx_0_1               ), //i
    .port_Al    (bl_0                  ), //i
    .port_Ah    (bh_0                  ), //i
    .port_aa    (bb_0                  ), //i
    .port_B_0   (port_c_0_0            ), //i
    .port_B_1   (port_c_0_1            ), //i
    .port_B_2   (port_c_0_2            ), //i
    .port_B_3   (port_c_0_3            ), //i
    .port_b_0_1 (scx_0_0               ), //i
    .port_b_1_1 (scx_0_1               ), //i
    .port_Bl    (cl_0                  ), //i
    .port_Bh    (ch_0                  ), //i
    .port_bb    (cc_0                  ), //i
    .port_o_0   (gF_MULS_4_193_port_o_0), //o
    .port_o_1   (gF_MULS_4_193_port_o_1), //o
    .port_o_2   (gF_MULS_4_193_port_o_2), //o
    .port_o_3   (gF_MULS_4_193_port_o_3)  //o
  );
  GF_MULS_4 gF_MULS_4_194 (
    .port_A_0   (port_b_0_0            ), //i
    .port_A_1   (port_b_0_1            ), //i
    .port_A_2   (port_b_0_2            ), //i
    .port_A_3   (port_b_0_3            ), //i
    .port_a_0_1 (sbx_0_0               ), //i
    .port_a_1_1 (sbx_0_1               ), //i
    .port_Al    (bl_0                  ), //i
    .port_Ah    (bh_0                  ), //i
    .port_aa    (bb_0                  ), //i
    .port_B_0   (port_a_1_0            ), //i
    .port_B_1   (port_a_1_1            ), //i
    .port_B_2   (port_a_1_2            ), //i
    .port_B_3   (port_a_1_3            ), //i
    .port_b_0_1 (sax_1_0               ), //i
    .port_b_1_1 (sax_1_1               ), //i
    .port_Bl    (al_1                  ), //i
    .port_Bh    (ah_1                  ), //i
    .port_bb    (aa_1                  ), //i
    .port_o_0   (gF_MULS_4_194_port_o_0), //o
    .port_o_1   (gF_MULS_4_194_port_o_1), //o
    .port_o_2   (gF_MULS_4_194_port_o_2), //o
    .port_o_3   (gF_MULS_4_194_port_o_3)  //o
  );
  GF_MULS_4 gF_MULS_4_195 (
    .port_A_0   (port_b_0_0            ), //i
    .port_A_1   (port_b_0_1            ), //i
    .port_A_2   (port_b_0_2            ), //i
    .port_A_3   (port_b_0_3            ), //i
    .port_a_0_1 (sbx_0_0               ), //i
    .port_a_1_1 (sbx_0_1               ), //i
    .port_Al    (bl_0                  ), //i
    .port_Ah    (bh_0                  ), //i
    .port_aa    (bb_0                  ), //i
    .port_B_0   (port_c_1_0            ), //i
    .port_B_1   (port_c_1_1            ), //i
    .port_B_2   (port_c_1_2            ), //i
    .port_B_3   (port_c_1_3            ), //i
    .port_b_0_1 (scx_1_0               ), //i
    .port_b_1_1 (scx_1_1               ), //i
    .port_Bl    (cl_1                  ), //i
    .port_Bh    (ch_1                  ), //i
    .port_bb    (cc_1                  ), //i
    .port_o_0   (gF_MULS_4_195_port_o_0), //o
    .port_o_1   (gF_MULS_4_195_port_o_1), //o
    .port_o_2   (gF_MULS_4_195_port_o_2), //o
    .port_o_3   (gF_MULS_4_195_port_o_3)  //o
  );
  GF_MULS_4 gF_MULS_4_196 (
    .port_A_0   (port_b_1_0            ), //i
    .port_A_1   (port_b_1_1            ), //i
    .port_A_2   (port_b_1_2            ), //i
    .port_A_3   (port_b_1_3            ), //i
    .port_a_0_1 (sbx_1_0               ), //i
    .port_a_1_1 (sbx_1_1               ), //i
    .port_Al    (bl_1                  ), //i
    .port_Ah    (bh_1                  ), //i
    .port_aa    (bb_1                  ), //i
    .port_B_0   (port_a_0_0            ), //i
    .port_B_1   (port_a_0_1            ), //i
    .port_B_2   (port_a_0_2            ), //i
    .port_B_3   (port_a_0_3            ), //i
    .port_b_0_1 (sax_0_0               ), //i
    .port_b_1_1 (sax_0_1               ), //i
    .port_Bl    (al_0                  ), //i
    .port_Bh    (ah_0                  ), //i
    .port_bb    (aa_0                  ), //i
    .port_o_0   (gF_MULS_4_196_port_o_0), //o
    .port_o_1   (gF_MULS_4_196_port_o_1), //o
    .port_o_2   (gF_MULS_4_196_port_o_2), //o
    .port_o_3   (gF_MULS_4_196_port_o_3)  //o
  );
  GF_MULS_4 gF_MULS_4_197 (
    .port_A_0   (port_b_1_0            ), //i
    .port_A_1   (port_b_1_1            ), //i
    .port_A_2   (port_b_1_2            ), //i
    .port_A_3   (port_b_1_3            ), //i
    .port_a_0_1 (sbx_1_0               ), //i
    .port_a_1_1 (sbx_1_1               ), //i
    .port_Al    (bl_1                  ), //i
    .port_Ah    (bh_1                  ), //i
    .port_aa    (bb_1                  ), //i
    .port_B_0   (port_c_0_0            ), //i
    .port_B_1   (port_c_0_1            ), //i
    .port_B_2   (port_c_0_2            ), //i
    .port_B_3   (port_c_0_3            ), //i
    .port_b_0_1 (scx_0_0               ), //i
    .port_b_1_1 (scx_0_1               ), //i
    .port_Bl    (cl_0                  ), //i
    .port_Bh    (ch_0                  ), //i
    .port_bb    (cc_0                  ), //i
    .port_o_0   (gF_MULS_4_197_port_o_0), //o
    .port_o_1   (gF_MULS_4_197_port_o_1), //o
    .port_o_2   (gF_MULS_4_197_port_o_2), //o
    .port_o_3   (gF_MULS_4_197_port_o_3)  //o
  );
  GF_MULS_4 gF_MULS_4_198 (
    .port_A_0   (port_b_1_0            ), //i
    .port_A_1   (port_b_1_1            ), //i
    .port_A_2   (port_b_1_2            ), //i
    .port_A_3   (port_b_1_3            ), //i
    .port_a_0_1 (sbx_1_0               ), //i
    .port_a_1_1 (sbx_1_1               ), //i
    .port_Al    (bl_1                  ), //i
    .port_Ah    (bh_1                  ), //i
    .port_aa    (bb_1                  ), //i
    .port_B_0   (port_a_1_0            ), //i
    .port_B_1   (port_a_1_1            ), //i
    .port_B_2   (port_a_1_2            ), //i
    .port_B_3   (port_a_1_3            ), //i
    .port_b_0_1 (sax_1_0               ), //i
    .port_b_1_1 (sax_1_1               ), //i
    .port_Bl    (al_1                  ), //i
    .port_Bh    (ah_1                  ), //i
    .port_bb    (aa_1                  ), //i
    .port_o_0   (gF_MULS_4_198_port_o_0), //o
    .port_o_1   (gF_MULS_4_198_port_o_1), //o
    .port_o_2   (gF_MULS_4_198_port_o_2), //o
    .port_o_3   (gF_MULS_4_198_port_o_3)  //o
  );
  GF_MULS_4 gF_MULS_4_199 (
    .port_A_0   (port_b_1_0            ), //i
    .port_A_1   (port_b_1_1            ), //i
    .port_A_2   (port_b_1_2            ), //i
    .port_A_3   (port_b_1_3            ), //i
    .port_a_0_1 (sbx_1_0               ), //i
    .port_a_1_1 (sbx_1_1               ), //i
    .port_Al    (bl_1                  ), //i
    .port_Ah    (bh_1                  ), //i
    .port_aa    (bb_1                  ), //i
    .port_B_0   (port_c_1_0            ), //i
    .port_B_1   (port_c_1_1            ), //i
    .port_B_2   (port_c_1_2            ), //i
    .port_B_3   (port_c_1_3            ), //i
    .port_b_0_1 (scx_1_0               ), //i
    .port_b_1_1 (scx_1_1               ), //i
    .port_Bl    (cl_1                  ), //i
    .port_Bh    (ch_1                  ), //i
    .port_bb    (cc_1                  ), //i
    .port_o_0   (gF_MULS_4_199_port_o_0), //o
    .port_o_1   (gF_MULS_4_199_port_o_1), //o
    .port_o_2   (gF_MULS_4_199_port_o_2), //o
    .port_o_3   (gF_MULS_4_199_port_o_3)  //o
  );
  assign sax_0_0 = (port_a_0_2 ^ port_a_0_0);
  assign sax_0_1 = (port_a_0_3 ^ port_a_0_1);
  assign al_0 = (port_a_0_1 ^ port_a_0_0);
  assign ah_0 = (port_a_0_3 ^ port_a_0_2);
  assign aa_0 = (sax_0_1 ^ sax_0_0);
  assign sbx_0_0 = (port_b_0_2 ^ port_b_0_0);
  assign sbx_0_1 = (port_b_0_3 ^ port_b_0_1);
  assign bl_0 = (port_b_0_1 ^ port_b_0_0);
  assign bh_0 = (port_b_0_3 ^ port_b_0_2);
  assign bb_0 = (sbx_0_1 ^ sbx_0_0);
  assign scx_0_0 = (port_c_0_2 ^ port_c_0_0);
  assign scx_0_1 = (port_c_0_3 ^ port_c_0_1);
  assign cl_0 = (port_c_0_1 ^ port_c_0_0);
  assign ch_0 = (port_c_0_3 ^ port_c_0_2);
  assign cc_0 = (scx_0_1 ^ scx_0_0);
  assign sax_1_0 = (port_a_1_2 ^ port_a_1_0);
  assign sax_1_1 = (port_a_1_3 ^ port_a_1_1);
  assign al_1 = (port_a_1_1 ^ port_a_1_0);
  assign ah_1 = (port_a_1_3 ^ port_a_1_2);
  assign aa_1 = (sax_1_1 ^ sax_1_0);
  assign sbx_1_0 = (port_b_1_2 ^ port_b_1_0);
  assign sbx_1_1 = (port_b_1_3 ^ port_b_1_1);
  assign bl_1 = (port_b_1_1 ^ port_b_1_0);
  assign bh_1 = (port_b_1_3 ^ port_b_1_2);
  assign bb_1 = (sbx_1_1 ^ sbx_1_0);
  assign scx_1_0 = (port_c_1_2 ^ port_c_1_0);
  assign scx_1_1 = (port_c_1_3 ^ port_c_1_1);
  assign cl_1 = (port_c_1_1 ^ port_c_1_0);
  assign ch_1 = (port_c_1_3 ^ port_c_1_2);
  assign cc_1 = (scx_1_1 ^ scx_1_0);
  assign outVal_0_0 = gF_MULS_4_193_port_o_0;
  assign outVal_0_1 = gF_MULS_4_193_port_o_1;
  assign outVal_0_2 = gF_MULS_4_193_port_o_2;
  assign outVal_0_3 = gF_MULS_4_193_port_o_3;
  assign outVal_0_4 = gF_MULS_4_192_port_o_0;
  assign outVal_0_5 = gF_MULS_4_192_port_o_1;
  assign outVal_0_6 = gF_MULS_4_192_port_o_2;
  assign outVal_0_7 = gF_MULS_4_192_port_o_3;
  assign outVal_2_0 = gF_MULS_4_195_port_o_0;
  assign outVal_2_1 = gF_MULS_4_195_port_o_1;
  assign outVal_2_2 = gF_MULS_4_195_port_o_2;
  assign outVal_2_3 = gF_MULS_4_195_port_o_3;
  assign outVal_2_4 = gF_MULS_4_194_port_o_0;
  assign outVal_2_5 = gF_MULS_4_194_port_o_1;
  assign outVal_2_6 = gF_MULS_4_194_port_o_2;
  assign outVal_2_7 = gF_MULS_4_194_port_o_3;
  assign outVal_1_0 = gF_MULS_4_197_port_o_0;
  assign outVal_1_1 = gF_MULS_4_197_port_o_1;
  assign outVal_1_2 = gF_MULS_4_197_port_o_2;
  assign outVal_1_3 = gF_MULS_4_197_port_o_3;
  assign outVal_1_4 = gF_MULS_4_196_port_o_0;
  assign outVal_1_5 = gF_MULS_4_196_port_o_1;
  assign outVal_1_6 = gF_MULS_4_196_port_o_2;
  assign outVal_1_7 = gF_MULS_4_196_port_o_3;
  assign outVal_3_0 = gF_MULS_4_199_port_o_0;
  assign outVal_3_1 = gF_MULS_4_199_port_o_1;
  assign outVal_3_2 = gF_MULS_4_199_port_o_2;
  assign outVal_3_3 = gF_MULS_4_199_port_o_3;
  assign outVal_3_4 = gF_MULS_4_198_port_o_0;
  assign outVal_3_5 = gF_MULS_4_198_port_o_1;
  assign outVal_3_6 = gF_MULS_4_198_port_o_2;
  assign outVal_3_7 = gF_MULS_4_198_port_o_3;
  assign refVal_0_0[0] = (outVal_0_0[0] ^ port_r_0_0);
  assign refVal_0_1[0] = (outVal_0_1[0] ^ port_r_0_1);
  assign refVal_0_2[0] = (outVal_0_2[0] ^ port_r_0_2);
  assign refVal_0_3[0] = (outVal_0_3[0] ^ port_r_0_3);
  assign refVal_0_4[0] = (outVal_0_4[0] ^ port_r_0_4);
  assign refVal_0_5[0] = (outVal_0_5[0] ^ port_r_0_5);
  assign refVal_0_6[0] = (outVal_0_6[0] ^ port_r_0_6);
  assign refVal_0_7[0] = (outVal_0_7[0] ^ port_r_0_7);
  assign refVal_1_0[0] = (outVal_1_0[0] ^ port_r_1_0);
  assign refVal_1_1[0] = (outVal_1_1[0] ^ port_r_1_1);
  assign refVal_1_2[0] = (outVal_1_2[0] ^ port_r_1_2);
  assign refVal_1_3[0] = (outVal_1_3[0] ^ port_r_1_3);
  assign refVal_1_4[0] = (outVal_1_4[0] ^ port_r_1_4);
  assign refVal_1_5[0] = (outVal_1_5[0] ^ port_r_1_5);
  assign refVal_1_6[0] = (outVal_1_6[0] ^ port_r_1_6);
  assign refVal_1_7[0] = (outVal_1_7[0] ^ port_r_1_7);
  assign refVal_2_0[0] = (outVal_2_0[0] ^ port_r_2_0);
  assign refVal_2_1[0] = (outVal_2_1[0] ^ port_r_2_1);
  assign refVal_2_2[0] = (outVal_2_2[0] ^ port_r_2_2);
  assign refVal_2_3[0] = (outVal_2_3[0] ^ port_r_2_3);
  assign refVal_2_4[0] = (outVal_2_4[0] ^ port_r_2_4);
  assign refVal_2_5[0] = (outVal_2_5[0] ^ port_r_2_5);
  assign refVal_2_6[0] = (outVal_2_6[0] ^ port_r_2_6);
  assign refVal_2_7[0] = (outVal_2_7[0] ^ port_r_2_7);
  assign refVal_3_0[0] = (outVal_3_0[0] ^ ((port_r_0_0 ^ port_r_1_0) ^ port_r_2_0));
  assign refVal_3_1[0] = (outVal_3_1[0] ^ ((port_r_0_1 ^ port_r_1_1) ^ port_r_2_1));
  assign refVal_3_2[0] = (outVal_3_2[0] ^ ((port_r_0_2 ^ port_r_1_2) ^ port_r_2_2));
  assign refVal_3_3[0] = (outVal_3_3[0] ^ ((port_r_0_3 ^ port_r_1_3) ^ port_r_2_3));
  assign refVal_3_4[0] = (outVal_3_4[0] ^ ((port_r_0_4 ^ port_r_1_4) ^ port_r_2_4));
  assign refVal_3_5[0] = (outVal_3_5[0] ^ ((port_r_0_5 ^ port_r_1_5) ^ port_r_2_5));
  assign refVal_3_6[0] = (outVal_3_6[0] ^ ((port_r_0_6 ^ port_r_1_6) ^ port_r_2_6));
  assign refVal_3_7[0] = (outVal_3_7[0] ^ ((port_r_0_7 ^ port_r_1_7) ^ port_r_2_7));
  assign port_y_0_0 = outReg_0_0;
  assign port_y_0_1 = outReg_0_1;
  assign port_y_0_2 = outReg_0_2;
  assign port_y_0_3 = outReg_0_3;
  assign port_y_0_4 = outReg_0_4;
  assign port_y_0_5 = outReg_0_5;
  assign port_y_0_6 = outReg_0_6;
  assign port_y_0_7 = outReg_0_7;
  assign port_y_1_0 = outReg_1_0;
  assign port_y_1_1 = outReg_1_1;
  assign port_y_1_2 = outReg_1_2;
  assign port_y_1_3 = outReg_1_3;
  assign port_y_1_4 = outReg_1_4;
  assign port_y_1_5 = outReg_1_5;
  assign port_y_1_6 = outReg_1_6;
  assign port_y_1_7 = outReg_1_7;
  assign port_y_2_0 = outReg_2_0;
  assign port_y_2_1 = outReg_2_1;
  assign port_y_2_2 = outReg_2_2;
  assign port_y_2_3 = outReg_2_3;
  assign port_y_2_4 = outReg_2_4;
  assign port_y_2_5 = outReg_2_5;
  assign port_y_2_6 = outReg_2_6;
  assign port_y_2_7 = outReg_2_7;
  assign port_y_3_0 = outReg_3_0;
  assign port_y_3_1 = outReg_3_1;
  assign port_y_3_2 = outReg_3_2;
  assign port_y_3_3 = outReg_3_3;
  assign port_y_3_4 = outReg_3_4;
  assign port_y_3_5 = outReg_3_5;
  assign port_y_3_6 = outReg_3_6;
  assign port_y_3_7 = outReg_3_7;
  always @(posedge clk) begin
    outReg_0_0 <= refVal_0_0;
    outReg_0_1 <= refVal_0_1;
    outReg_0_2 <= refVal_0_2;
    outReg_0_3 <= refVal_0_3;
    outReg_0_4 <= refVal_0_4;
    outReg_0_5 <= refVal_0_5;
    outReg_0_6 <= refVal_0_6;
    outReg_0_7 <= refVal_0_7;
    outReg_1_0 <= refVal_1_0;
    outReg_1_1 <= refVal_1_1;
    outReg_1_2 <= refVal_1_2;
    outReg_1_3 <= refVal_1_3;
    outReg_1_4 <= refVal_1_4;
    outReg_1_5 <= refVal_1_5;
    outReg_1_6 <= refVal_1_6;
    outReg_1_7 <= refVal_1_7;
    outReg_2_0 <= refVal_2_0;
    outReg_2_1 <= refVal_2_1;
    outReg_2_2 <= refVal_2_2;
    outReg_2_3 <= refVal_2_3;
    outReg_2_4 <= refVal_2_4;
    outReg_2_5 <= refVal_2_5;
    outReg_2_6 <= refVal_2_6;
    outReg_2_7 <= refVal_2_7;
    outReg_3_0 <= refVal_3_0;
    outReg_3_1 <= refVal_3_1;
    outReg_3_2 <= refVal_3_2;
    outReg_3_3 <= refVal_3_3;
    outReg_3_4 <= refVal_3_4;
    outReg_3_5 <= refVal_3_5;
    outReg_3_6 <= refVal_3_6;
    outReg_3_7 <= refVal_3_7;
  end


endmodule

module CMS_stage4 (
  input      [0:0]    port_a_0_0,
  input      [0:0]    port_a_0_1,
  input      [0:0]    port_a_1_0,
  input      [0:0]    port_a_1_1,
  input      [0:0]    port_b_0_0,
  input      [0:0]    port_b_0_1,
  input      [0:0]    port_b_1_0,
  input      [0:0]    port_b_1_1,
  input      [0:0]    port_c_0_0,
  input      [0:0]    port_c_0_1,
  input      [0:0]    port_c_1_0,
  input      [0:0]    port_c_1_1,
  input               port_r_0_0,
  input               port_r_0_1,
  input               port_r_0_2,
  input               port_r_0_3,
  input               port_r_1_0,
  input               port_r_1_1,
  input               port_r_1_2,
  input               port_r_1_3,
  input               port_r_2_0,
  input               port_r_2_1,
  input               port_r_2_2,
  input               port_r_2_3,
  output     [0:0]    port_y_0_0,
  output     [0:0]    port_y_0_1,
  output     [0:0]    port_y_0_2,
  output     [0:0]    port_y_0_3,
  output     [0:0]    port_y_1_0,
  output     [0:0]    port_y_1_1,
  output     [0:0]    port_y_1_2,
  output     [0:0]    port_y_1_3,
  output     [0:0]    port_y_2_0,
  output     [0:0]    port_y_2_1,
  output     [0:0]    port_y_2_2,
  output     [0:0]    port_y_2_3,
  output     [0:0]    port_y_3_0,
  output     [0:0]    port_y_3_1,
  output     [0:0]    port_y_3_2,
  output     [0:0]    port_y_3_3,
  input               clk,
  input               reset
);

  wire       [0:0]    sq_0_port_o_0;
  wire       [0:0]    sq_0_port_o_1;
  wire       [0:0]    sq_1_port_o_0;
  wire       [0:0]    sq_1_port_o_1;
  wire       [0:0]    gF_MULS_2_576_port_o_0;
  wire       [0:0]    gF_MULS_2_576_port_o_1;
  wire       [0:0]    gF_MULS_2_577_port_o_0;
  wire       [0:0]    gF_MULS_2_577_port_o_1;
  wire       [0:0]    gF_MULS_2_578_port_o_0;
  wire       [0:0]    gF_MULS_2_578_port_o_1;
  wire       [0:0]    gF_MULS_2_579_port_o_0;
  wire       [0:0]    gF_MULS_2_579_port_o_1;
  wire       [0:0]    gF_MULS_2_580_port_o_0;
  wire       [0:0]    gF_MULS_2_580_port_o_1;
  wire       [0:0]    gF_MULS_2_581_port_o_0;
  wire       [0:0]    gF_MULS_2_581_port_o_1;
  wire       [0:0]    gF_MULS_2_582_port_o_0;
  wire       [0:0]    gF_MULS_2_582_port_o_1;
  wire       [0:0]    gF_MULS_2_583_port_o_0;
  wire       [0:0]    gF_MULS_2_583_port_o_1;
  reg        [0:0]    outReg_0_0;
  reg        [0:0]    outReg_0_1;
  reg        [0:0]    outReg_0_2;
  reg        [0:0]    outReg_0_3;
  reg        [0:0]    outReg_1_0;
  reg        [0:0]    outReg_1_1;
  reg        [0:0]    outReg_1_2;
  reg        [0:0]    outReg_1_3;
  reg        [0:0]    outReg_2_0;
  reg        [0:0]    outReg_2_1;
  reg        [0:0]    outReg_2_2;
  reg        [0:0]    outReg_2_3;
  reg        [0:0]    outReg_3_0;
  reg        [0:0]    outReg_3_1;
  reg        [0:0]    outReg_3_2;
  reg        [0:0]    outReg_3_3;
  wire       [0:0]    outVal_0_0;
  wire       [0:0]    outVal_0_1;
  wire       [0:0]    outVal_0_2;
  wire       [0:0]    outVal_0_3;
  wire       [0:0]    outVal_1_0;
  wire       [0:0]    outVal_1_1;
  wire       [0:0]    outVal_1_2;
  wire       [0:0]    outVal_1_3;
  wire       [0:0]    outVal_2_0;
  wire       [0:0]    outVal_2_1;
  wire       [0:0]    outVal_2_2;
  wire       [0:0]    outVal_2_3;
  wire       [0:0]    outVal_3_0;
  wire       [0:0]    outVal_3_1;
  wire       [0:0]    outVal_3_2;
  wire       [0:0]    outVal_3_3;
  wire       [0:0]    refVal_0_0;
  wire       [0:0]    refVal_0_1;
  wire       [0:0]    refVal_0_2;
  wire       [0:0]    refVal_0_3;
  wire       [0:0]    refVal_1_0;
  wire       [0:0]    refVal_1_1;
  wire       [0:0]    refVal_1_2;
  wire       [0:0]    refVal_1_3;
  wire       [0:0]    refVal_2_0;
  wire       [0:0]    refVal_2_1;
  wire       [0:0]    refVal_2_2;
  wire       [0:0]    refVal_2_3;
  wire       [0:0]    refVal_3_0;
  wire       [0:0]    refVal_3_1;
  wire       [0:0]    refVal_3_2;
  wire       [0:0]    refVal_3_3;
  wire       [0:0]    sq_0_0;
  wire       [0:0]    sq_0_1;
  wire       [0:0]    sq_1_0;
  wire       [0:0]    sq_1_1;
  wire       [0:0]    sax_0;
  wire       [0:0]    sax_1;
  wire       [0:0]    sqx_0;
  wire       [0:0]    sqx_1;
  wire       [0:0]    scx_0;
  wire       [0:0]    scx_1;

  GF_SQ_2 sq_0 (
    .port_i_0 (port_b_0_0   ), //i
    .port_i_1 (port_b_0_1   ), //i
    .port_o_0 (sq_0_port_o_0), //o
    .port_o_1 (sq_0_port_o_1)  //o
  );
  GF_SQ_2 sq_1 (
    .port_i_0 (port_b_1_0   ), //i
    .port_i_1 (port_b_1_1   ), //i
    .port_o_0 (sq_1_port_o_0), //o
    .port_o_1 (sq_1_port_o_1)  //o
  );
  GF_MULS_2 gF_MULS_2_576 (
    .port_a_0 (port_a_0_0            ), //i
    .port_a_1 (port_a_0_1            ), //i
    .port_ab  (sax_0                 ), //i
    .port_b_0 (sq_0_0                ), //i
    .port_b_1 (sq_0_1                ), //i
    .port_cd  (sqx_0                 ), //i
    .port_o_0 (gF_MULS_2_576_port_o_0), //o
    .port_o_1 (gF_MULS_2_576_port_o_1)  //o
  );
  GF_MULS_2 gF_MULS_2_577 (
    .port_a_0 (port_c_0_0            ), //i
    .port_a_1 (port_c_0_1            ), //i
    .port_ab  (scx_0                 ), //i
    .port_b_0 (sq_0_0                ), //i
    .port_b_1 (sq_0_1                ), //i
    .port_cd  (sqx_0                 ), //i
    .port_o_0 (gF_MULS_2_577_port_o_0), //o
    .port_o_1 (gF_MULS_2_577_port_o_1)  //o
  );
  GF_MULS_2 gF_MULS_2_578 (
    .port_a_0 (port_a_0_0            ), //i
    .port_a_1 (port_a_0_1            ), //i
    .port_ab  (sax_0                 ), //i
    .port_b_0 (sq_1_0                ), //i
    .port_b_1 (sq_1_1                ), //i
    .port_cd  (sqx_1                 ), //i
    .port_o_0 (gF_MULS_2_578_port_o_0), //o
    .port_o_1 (gF_MULS_2_578_port_o_1)  //o
  );
  GF_MULS_2 gF_MULS_2_579 (
    .port_a_0 (port_c_0_0            ), //i
    .port_a_1 (port_c_0_1            ), //i
    .port_ab  (scx_0                 ), //i
    .port_b_0 (sq_1_0                ), //i
    .port_b_1 (sq_1_1                ), //i
    .port_cd  (sqx_1                 ), //i
    .port_o_0 (gF_MULS_2_579_port_o_0), //o
    .port_o_1 (gF_MULS_2_579_port_o_1)  //o
  );
  GF_MULS_2 gF_MULS_2_580 (
    .port_a_0 (port_a_1_0            ), //i
    .port_a_1 (port_a_1_1            ), //i
    .port_ab  (sax_1                 ), //i
    .port_b_0 (sq_0_0                ), //i
    .port_b_1 (sq_0_1                ), //i
    .port_cd  (sqx_0                 ), //i
    .port_o_0 (gF_MULS_2_580_port_o_0), //o
    .port_o_1 (gF_MULS_2_580_port_o_1)  //o
  );
  GF_MULS_2 gF_MULS_2_581 (
    .port_a_0 (port_c_1_0            ), //i
    .port_a_1 (port_c_1_1            ), //i
    .port_ab  (scx_1                 ), //i
    .port_b_0 (sq_0_0                ), //i
    .port_b_1 (sq_0_1                ), //i
    .port_cd  (sqx_0                 ), //i
    .port_o_0 (gF_MULS_2_581_port_o_0), //o
    .port_o_1 (gF_MULS_2_581_port_o_1)  //o
  );
  GF_MULS_2 gF_MULS_2_582 (
    .port_a_0 (port_a_1_0            ), //i
    .port_a_1 (port_a_1_1            ), //i
    .port_ab  (sax_1                 ), //i
    .port_b_0 (sq_1_0                ), //i
    .port_b_1 (sq_1_1                ), //i
    .port_cd  (sqx_1                 ), //i
    .port_o_0 (gF_MULS_2_582_port_o_0), //o
    .port_o_1 (gF_MULS_2_582_port_o_1)  //o
  );
  GF_MULS_2 gF_MULS_2_583 (
    .port_a_0 (port_c_1_0            ), //i
    .port_a_1 (port_c_1_1            ), //i
    .port_ab  (scx_1                 ), //i
    .port_b_0 (sq_1_0                ), //i
    .port_b_1 (sq_1_1                ), //i
    .port_cd  (sqx_1                 ), //i
    .port_o_0 (gF_MULS_2_583_port_o_0), //o
    .port_o_1 (gF_MULS_2_583_port_o_1)  //o
  );
  assign sq_0_0 = sq_0_port_o_0;
  assign sq_0_1 = sq_0_port_o_1;
  assign sq_1_0 = sq_1_port_o_0;
  assign sq_1_1 = sq_1_port_o_1;
  assign sax_0 = (port_a_0_0 ^ port_a_0_1);
  assign sqx_0 = (sq_0_0 ^ sq_0_1);
  assign scx_0 = (port_c_0_0 ^ port_c_0_1);
  assign sax_1 = (port_a_1_0 ^ port_a_1_1);
  assign sqx_1 = (sq_1_0 ^ sq_1_1);
  assign scx_1 = (port_c_1_0 ^ port_c_1_1);
  assign outVal_0_0 = gF_MULS_2_576_port_o_0;
  assign outVal_0_1 = gF_MULS_2_576_port_o_1;
  assign outVal_0_2 = gF_MULS_2_577_port_o_0;
  assign outVal_0_3 = gF_MULS_2_577_port_o_1;
  assign outVal_2_0 = gF_MULS_2_578_port_o_0;
  assign outVal_2_1 = gF_MULS_2_578_port_o_1;
  assign outVal_2_2 = gF_MULS_2_579_port_o_0;
  assign outVal_2_3 = gF_MULS_2_579_port_o_1;
  assign outVal_1_0 = gF_MULS_2_580_port_o_0;
  assign outVal_1_1 = gF_MULS_2_580_port_o_1;
  assign outVal_1_2 = gF_MULS_2_581_port_o_0;
  assign outVal_1_3 = gF_MULS_2_581_port_o_1;
  assign outVal_3_0 = gF_MULS_2_582_port_o_0;
  assign outVal_3_1 = gF_MULS_2_582_port_o_1;
  assign outVal_3_2 = gF_MULS_2_583_port_o_0;
  assign outVal_3_3 = gF_MULS_2_583_port_o_1;
  assign refVal_0_0[0] = (outVal_0_0[0] ^ port_r_0_0);
  assign refVal_0_1[0] = (outVal_0_1[0] ^ port_r_0_1);
  assign refVal_0_2[0] = (outVal_0_2[0] ^ port_r_0_2);
  assign refVal_0_3[0] = (outVal_0_3[0] ^ port_r_0_3);
  assign refVal_1_0[0] = (outVal_1_0[0] ^ port_r_1_0);
  assign refVal_1_1[0] = (outVal_1_1[0] ^ port_r_1_1);
  assign refVal_1_2[0] = (outVal_1_2[0] ^ port_r_1_2);
  assign refVal_1_3[0] = (outVal_1_3[0] ^ port_r_1_3);
  assign refVal_2_0[0] = (outVal_2_0[0] ^ port_r_2_0);
  assign refVal_2_1[0] = (outVal_2_1[0] ^ port_r_2_1);
  assign refVal_2_2[0] = (outVal_2_2[0] ^ port_r_2_2);
  assign refVal_2_3[0] = (outVal_2_3[0] ^ port_r_2_3);
  assign refVal_3_0[0] = (outVal_3_0[0] ^ ((port_r_0_0 ^ port_r_1_0) ^ port_r_2_0));
  assign refVal_3_1[0] = (outVal_3_1[0] ^ ((port_r_0_1 ^ port_r_1_1) ^ port_r_2_1));
  assign refVal_3_2[0] = (outVal_3_2[0] ^ ((port_r_0_2 ^ port_r_1_2) ^ port_r_2_2));
  assign refVal_3_3[0] = (outVal_3_3[0] ^ ((port_r_0_3 ^ port_r_1_3) ^ port_r_2_3));
  assign port_y_0_0 = outReg_0_0;
  assign port_y_0_1 = outReg_0_1;
  assign port_y_0_2 = outReg_0_2;
  assign port_y_0_3 = outReg_0_3;
  assign port_y_1_0 = outReg_1_0;
  assign port_y_1_1 = outReg_1_1;
  assign port_y_1_2 = outReg_1_2;
  assign port_y_1_3 = outReg_1_3;
  assign port_y_2_0 = outReg_2_0;
  assign port_y_2_1 = outReg_2_1;
  assign port_y_2_2 = outReg_2_2;
  assign port_y_2_3 = outReg_2_3;
  assign port_y_3_0 = outReg_3_0;
  assign port_y_3_1 = outReg_3_1;
  assign port_y_3_2 = outReg_3_2;
  assign port_y_3_3 = outReg_3_3;
  always @(posedge clk) begin
    outReg_0_0 <= refVal_0_0;
    outReg_0_1 <= refVal_0_1;
    outReg_0_2 <= refVal_0_2;
    outReg_0_3 <= refVal_0_3;
    outReg_1_0 <= refVal_1_0;
    outReg_1_1 <= refVal_1_1;
    outReg_1_2 <= refVal_1_2;
    outReg_1_3 <= refVal_1_3;
    outReg_2_0 <= refVal_2_0;
    outReg_2_1 <= refVal_2_1;
    outReg_2_2 <= refVal_2_2;
    outReg_2_3 <= refVal_2_3;
    outReg_3_0 <= refVal_3_0;
    outReg_3_1 <= refVal_3_1;
    outReg_3_2 <= refVal_3_2;
    outReg_3_3 <= refVal_3_3;
  end


endmodule

module CMS_stage3 (
  input      [0:0]    port_a_0_0,
  input      [0:0]    port_a_0_1,
  input      [0:0]    port_a_1_0,
  input      [0:0]    port_a_1_1,
  input      [0:0]    port_b_0_0,
  input      [0:0]    port_b_0_1,
  input      [0:0]    port_b_1_0,
  input      [0:0]    port_b_1_1,
  input               port_r_0_0,
  input               port_r_0_1,
  input               port_r_1_0,
  input               port_r_1_1,
  input               port_r_2_0,
  input               port_r_2_1,
  output     [0:0]    port_y_0_0,
  output     [0:0]    port_y_0_1,
  output     [0:0]    port_y_1_0,
  output     [0:0]    port_y_1_1,
  output     [0:0]    port_y_2_0,
  output     [0:0]    port_y_2_1,
  output     [0:0]    port_y_3_0,
  output     [0:0]    port_y_3_1,
  input               clk,
  input               reset
);

  wire       [0:0]    gF_SQ_2_128_port_i_0;
  wire       [0:0]    gF_SQ_2_128_port_i_1;
  wire       [0:0]    gF_SQ_2_129_port_i_0;
  wire       [0:0]    gF_SQ_2_129_port_i_1;
  wire       [0:0]    gF_SQ_2_128_port_o_0;
  wire       [0:0]    gF_SQ_2_128_port_o_1;
  wire       [0:0]    gF_SCLW2_2_32_port_o_0;
  wire       [0:0]    gF_SCLW2_2_32_port_o_1;
  wire       [0:0]    gF_SQ_2_129_port_o_0;
  wire       [0:0]    gF_SQ_2_129_port_o_1;
  wire       [0:0]    gF_SCLW2_2_33_port_o_0;
  wire       [0:0]    gF_SCLW2_2_33_port_o_1;
  wire       [0:0]    gF_MULS_2_576_port_o_0;
  wire       [0:0]    gF_MULS_2_576_port_o_1;
  wire       [0:0]    gF_MULS_2_577_port_o_0;
  wire       [0:0]    gF_MULS_2_577_port_o_1;
  wire       [0:0]    gF_MULS_2_578_port_o_0;
  wire       [0:0]    gF_MULS_2_578_port_o_1;
  wire       [0:0]    gF_MULS_2_579_port_o_0;
  wire       [0:0]    gF_MULS_2_579_port_o_1;
  reg        [0:0]    outReg_0_0;
  reg        [0:0]    outReg_0_1;
  reg        [0:0]    outReg_1_0;
  reg        [0:0]    outReg_1_1;
  reg        [0:0]    outReg_2_0;
  reg        [0:0]    outReg_2_1;
  reg        [0:0]    outReg_3_0;
  reg        [0:0]    outReg_3_1;
  wire       [0:0]    outVal_0_0;
  wire       [0:0]    outVal_0_1;
  wire       [0:0]    outVal_1_0;
  wire       [0:0]    outVal_1_1;
  wire       [0:0]    outVal_2_0;
  wire       [0:0]    outVal_2_1;
  wire       [0:0]    outVal_3_0;
  wire       [0:0]    outVal_3_1;
  wire       [0:0]    refVal_0_0;
  wire       [0:0]    refVal_0_1;
  wire       [0:0]    refVal_1_0;
  wire       [0:0]    refVal_1_1;
  wire       [0:0]    refVal_2_0;
  wire       [0:0]    refVal_2_1;
  wire       [0:0]    refVal_3_0;
  wire       [0:0]    refVal_3_1;
  wire       [0:0]    sax_0;
  wire       [0:0]    sax_1;
  wire       [0:0]    sbx_0;
  wire       [0:0]    sbx_1;
  wire       [0:0]    sq_0_0;
  wire       [0:0]    sq_0_1;
  wire       [0:0]    sq_1_0;
  wire       [0:0]    sq_1_1;

  GF_SQ_2 gF_SQ_2_128 (
    .port_i_0 (gF_SQ_2_128_port_i_0), //i
    .port_i_1 (gF_SQ_2_128_port_i_1), //i
    .port_o_0 (gF_SQ_2_128_port_o_0), //o
    .port_o_1 (gF_SQ_2_128_port_o_1)  //o
  );
  GF_SCLW2_2 gF_SCLW2_2_32 (
    .port_i_0 (gF_SQ_2_128_port_o_0  ), //i
    .port_i_1 (gF_SQ_2_128_port_o_1  ), //i
    .port_o_0 (gF_SCLW2_2_32_port_o_0), //o
    .port_o_1 (gF_SCLW2_2_32_port_o_1)  //o
  );
  GF_SQ_2 gF_SQ_2_129 (
    .port_i_0 (gF_SQ_2_129_port_i_0), //i
    .port_i_1 (gF_SQ_2_129_port_i_1), //i
    .port_o_0 (gF_SQ_2_129_port_o_0), //o
    .port_o_1 (gF_SQ_2_129_port_o_1)  //o
  );
  GF_SCLW2_2 gF_SCLW2_2_33 (
    .port_i_0 (gF_SQ_2_129_port_o_0  ), //i
    .port_i_1 (gF_SQ_2_129_port_o_1  ), //i
    .port_o_0 (gF_SCLW2_2_33_port_o_0), //o
    .port_o_1 (gF_SCLW2_2_33_port_o_1)  //o
  );
  GF_MULS_2 gF_MULS_2_576 (
    .port_a_0 (port_a_0_0            ), //i
    .port_a_1 (port_a_0_1            ), //i
    .port_ab  (sax_0                 ), //i
    .port_b_0 (port_b_0_0            ), //i
    .port_b_1 (port_b_0_1            ), //i
    .port_cd  (sbx_0                 ), //i
    .port_o_0 (gF_MULS_2_576_port_o_0), //o
    .port_o_1 (gF_MULS_2_576_port_o_1)  //o
  );
  GF_MULS_2 gF_MULS_2_577 (
    .port_a_0 (port_a_0_0            ), //i
    .port_a_1 (port_a_0_1            ), //i
    .port_ab  (sax_0                 ), //i
    .port_b_0 (port_b_1_0            ), //i
    .port_b_1 (port_b_1_1            ), //i
    .port_cd  (sbx_1                 ), //i
    .port_o_0 (gF_MULS_2_577_port_o_0), //o
    .port_o_1 (gF_MULS_2_577_port_o_1)  //o
  );
  GF_MULS_2 gF_MULS_2_578 (
    .port_a_0 (port_a_1_0            ), //i
    .port_a_1 (port_a_1_1            ), //i
    .port_ab  (sax_1                 ), //i
    .port_b_0 (port_b_0_0            ), //i
    .port_b_1 (port_b_0_1            ), //i
    .port_cd  (sbx_0                 ), //i
    .port_o_0 (gF_MULS_2_578_port_o_0), //o
    .port_o_1 (gF_MULS_2_578_port_o_1)  //o
  );
  GF_MULS_2 gF_MULS_2_579 (
    .port_a_0 (port_a_1_0            ), //i
    .port_a_1 (port_a_1_1            ), //i
    .port_ab  (sax_1                 ), //i
    .port_b_0 (port_b_1_0            ), //i
    .port_b_1 (port_b_1_1            ), //i
    .port_cd  (sbx_1                 ), //i
    .port_o_0 (gF_MULS_2_579_port_o_0), //o
    .port_o_1 (gF_MULS_2_579_port_o_1)  //o
  );
  assign sax_0 = (port_a_0_0 ^ port_a_0_1);
  assign sbx_0 = (port_b_0_0 ^ port_b_0_1);
  assign sax_1 = (port_a_1_0 ^ port_a_1_1);
  assign sbx_1 = (port_b_1_0 ^ port_b_1_1);
  assign gF_SQ_2_128_port_i_0 = (port_a_0_0 ^ port_b_0_0);
  assign gF_SQ_2_128_port_i_1 = (port_a_0_1 ^ port_b_0_1);
  assign sq_0_0 = gF_SCLW2_2_32_port_o_0;
  assign sq_0_1 = gF_SCLW2_2_32_port_o_1;
  assign gF_SQ_2_129_port_i_0 = (port_a_1_0 ^ port_b_1_0);
  assign gF_SQ_2_129_port_i_1 = (port_a_1_1 ^ port_b_1_1);
  assign sq_1_0 = gF_SCLW2_2_33_port_o_0;
  assign sq_1_1 = gF_SCLW2_2_33_port_o_1;
  assign outVal_0_0 = (gF_MULS_2_576_port_o_0 ^ sq_0_0);
  assign outVal_0_1 = (gF_MULS_2_576_port_o_1 ^ sq_0_1);
  assign outVal_2_0 = gF_MULS_2_577_port_o_0;
  assign outVal_2_1 = gF_MULS_2_577_port_o_1;
  assign outVal_1_0 = gF_MULS_2_578_port_o_0;
  assign outVal_1_1 = gF_MULS_2_578_port_o_1;
  assign outVal_3_0 = (gF_MULS_2_579_port_o_0 ^ sq_1_0);
  assign outVal_3_1 = (gF_MULS_2_579_port_o_1 ^ sq_1_1);
  assign refVal_0_0[0] = (outVal_0_0[0] ^ port_r_0_0);
  assign refVal_0_1[0] = (outVal_0_1[0] ^ port_r_0_1);
  assign refVal_1_0[0] = (outVal_1_0[0] ^ port_r_1_0);
  assign refVal_1_1[0] = (outVal_1_1[0] ^ port_r_1_1);
  assign refVal_2_0[0] = (outVal_2_0[0] ^ port_r_2_0);
  assign refVal_2_1[0] = (outVal_2_1[0] ^ port_r_2_1);
  assign refVal_3_0[0] = (outVal_3_0[0] ^ ((port_r_0_0 ^ port_r_1_0) ^ port_r_2_0));
  assign refVal_3_1[0] = (outVal_3_1[0] ^ ((port_r_0_1 ^ port_r_1_1) ^ port_r_2_1));
  assign port_y_0_0 = outReg_0_0;
  assign port_y_0_1 = outReg_0_1;
  assign port_y_1_0 = outReg_1_0;
  assign port_y_1_1 = outReg_1_1;
  assign port_y_2_0 = outReg_2_0;
  assign port_y_2_1 = outReg_2_1;
  assign port_y_3_0 = outReg_3_0;
  assign port_y_3_1 = outReg_3_1;
  always @(posedge clk) begin
    outReg_0_0 <= refVal_0_0;
    outReg_0_1 <= refVal_0_1;
    outReg_1_0 <= refVal_1_0;
    outReg_1_1 <= refVal_1_1;
    outReg_2_0 <= refVal_2_0;
    outReg_2_1 <= refVal_2_1;
    outReg_3_0 <= refVal_3_0;
    outReg_3_1 <= refVal_3_1;
  end


endmodule

module CMS_stage2 (
  input      [0:0]    port_a_0_0,
  input      [0:0]    port_a_0_1,
  input      [0:0]    port_a_0_2,
  input      [0:0]    port_a_0_3,
  input      [0:0]    port_a_1_0,
  input      [0:0]    port_a_1_1,
  input      [0:0]    port_a_1_2,
  input      [0:0]    port_a_1_3,
  input      [0:0]    port_b_0_0,
  input      [0:0]    port_b_0_1,
  input      [0:0]    port_b_0_2,
  input      [0:0]    port_b_0_3,
  input      [0:0]    port_b_1_0,
  input      [0:0]    port_b_1_1,
  input      [0:0]    port_b_1_2,
  input      [0:0]    port_b_1_3,
  input               port_r_0_0,
  input               port_r_0_1,
  input               port_r_0_2,
  input               port_r_0_3,
  input               port_r_1_0,
  input               port_r_1_1,
  input               port_r_1_2,
  input               port_r_1_3,
  input               port_r_2_0,
  input               port_r_2_1,
  input               port_r_2_2,
  input               port_r_2_3,
  output     [0:0]    port_y_0_0,
  output     [0:0]    port_y_0_1,
  output     [0:0]    port_y_0_2,
  output     [0:0]    port_y_0_3,
  output     [0:0]    port_y_1_0,
  output     [0:0]    port_y_1_1,
  output     [0:0]    port_y_1_2,
  output     [0:0]    port_y_1_3,
  output     [0:0]    port_y_2_0,
  output     [0:0]    port_y_2_1,
  output     [0:0]    port_y_2_2,
  output     [0:0]    port_y_2_3,
  output     [0:0]    port_y_3_0,
  output     [0:0]    port_y_3_1,
  output     [0:0]    port_y_3_2,
  output     [0:0]    port_y_3_3,
  input               clk,
  input               reset
);

  wire       [0:0]    sq_0_port_i_0;
  wire       [0:0]    sq_0_port_i_1;
  wire       [0:0]    sq_0_port_i_2;
  wire       [0:0]    sq_0_port_i_3;
  wire       [0:0]    sq_1_port_i_0;
  wire       [0:0]    sq_1_port_i_1;
  wire       [0:0]    sq_1_port_i_2;
  wire       [0:0]    sq_1_port_i_3;
  wire       [0:0]    sq_0_port_o_0;
  wire       [0:0]    sq_0_port_o_1;
  wire       [0:0]    sq_0_port_o_2;
  wire       [0:0]    sq_0_port_o_3;
  wire       [0:0]    sq_1_port_o_0;
  wire       [0:0]    sq_1_port_o_1;
  wire       [0:0]    sq_1_port_o_2;
  wire       [0:0]    sq_1_port_o_3;
  wire       [0:0]    gF_MULS_4_192_port_o_0;
  wire       [0:0]    gF_MULS_4_192_port_o_1;
  wire       [0:0]    gF_MULS_4_192_port_o_2;
  wire       [0:0]    gF_MULS_4_192_port_o_3;
  wire       [0:0]    gF_MULS_4_193_port_o_0;
  wire       [0:0]    gF_MULS_4_193_port_o_1;
  wire       [0:0]    gF_MULS_4_193_port_o_2;
  wire       [0:0]    gF_MULS_4_193_port_o_3;
  wire       [0:0]    gF_MULS_4_194_port_o_0;
  wire       [0:0]    gF_MULS_4_194_port_o_1;
  wire       [0:0]    gF_MULS_4_194_port_o_2;
  wire       [0:0]    gF_MULS_4_194_port_o_3;
  wire       [0:0]    gF_MULS_4_195_port_o_0;
  wire       [0:0]    gF_MULS_4_195_port_o_1;
  wire       [0:0]    gF_MULS_4_195_port_o_2;
  wire       [0:0]    gF_MULS_4_195_port_o_3;
  reg        [0:0]    outReg_0_0;
  reg        [0:0]    outReg_0_1;
  reg        [0:0]    outReg_0_2;
  reg        [0:0]    outReg_0_3;
  reg        [0:0]    outReg_1_0;
  reg        [0:0]    outReg_1_1;
  reg        [0:0]    outReg_1_2;
  reg        [0:0]    outReg_1_3;
  reg        [0:0]    outReg_2_0;
  reg        [0:0]    outReg_2_1;
  reg        [0:0]    outReg_2_2;
  reg        [0:0]    outReg_2_3;
  reg        [0:0]    outReg_3_0;
  reg        [0:0]    outReg_3_1;
  reg        [0:0]    outReg_3_2;
  reg        [0:0]    outReg_3_3;
  wire       [0:0]    outVal_0_0;
  wire       [0:0]    outVal_0_1;
  wire       [0:0]    outVal_0_2;
  wire       [0:0]    outVal_0_3;
  wire       [0:0]    outVal_1_0;
  wire       [0:0]    outVal_1_1;
  wire       [0:0]    outVal_1_2;
  wire       [0:0]    outVal_1_3;
  wire       [0:0]    outVal_2_0;
  wire       [0:0]    outVal_2_1;
  wire       [0:0]    outVal_2_2;
  wire       [0:0]    outVal_2_3;
  wire       [0:0]    outVal_3_0;
  wire       [0:0]    outVal_3_1;
  wire       [0:0]    outVal_3_2;
  wire       [0:0]    outVal_3_3;
  wire       [0:0]    refVal_0_0;
  wire       [0:0]    refVal_0_1;
  wire       [0:0]    refVal_0_2;
  wire       [0:0]    refVal_0_3;
  wire       [0:0]    refVal_1_0;
  wire       [0:0]    refVal_1_1;
  wire       [0:0]    refVal_1_2;
  wire       [0:0]    refVal_1_3;
  wire       [0:0]    refVal_2_0;
  wire       [0:0]    refVal_2_1;
  wire       [0:0]    refVal_2_2;
  wire       [0:0]    refVal_2_3;
  wire       [0:0]    refVal_3_0;
  wire       [0:0]    refVal_3_1;
  wire       [0:0]    refVal_3_2;
  wire       [0:0]    refVal_3_3;
  wire       [0:0]    sq_0_0;
  wire       [0:0]    sq_0_1;
  wire       [0:0]    sq_0_2;
  wire       [0:0]    sq_0_3;
  wire       [0:0]    sq_1_0;
  wire       [0:0]    sq_1_1;
  wire       [0:0]    sq_1_2;
  wire       [0:0]    sq_1_3;
  wire       [0:0]    sax_0_0;
  wire       [0:0]    sax_0_1;
  wire       [0:0]    sax_1_0;
  wire       [0:0]    sax_1_1;
  wire       [0:0]    sbx_0_0;
  wire       [0:0]    sbx_0_1;
  wire       [0:0]    sbx_1_0;
  wire       [0:0]    sbx_1_1;
  wire       [0:0]    al_0;
  wire       [0:0]    al_1;
  wire       [0:0]    ah_0;
  wire       [0:0]    ah_1;
  wire       [0:0]    aa_0;
  wire       [0:0]    aa_1;
  wire       [0:0]    bl_0;
  wire       [0:0]    bl_1;
  wire       [0:0]    bh_0;
  wire       [0:0]    bh_1;
  wire       [0:0]    bb_0;
  wire       [0:0]    bb_1;

  GF_SQ_SCL_4 sq_0 (
    .port_i_0 (sq_0_port_i_0), //i
    .port_i_1 (sq_0_port_i_1), //i
    .port_i_2 (sq_0_port_i_2), //i
    .port_i_3 (sq_0_port_i_3), //i
    .port_o_0 (sq_0_port_o_0), //o
    .port_o_1 (sq_0_port_o_1), //o
    .port_o_2 (sq_0_port_o_2), //o
    .port_o_3 (sq_0_port_o_3)  //o
  );
  GF_SQ_SCL_4 sq_1 (
    .port_i_0 (sq_1_port_i_0), //i
    .port_i_1 (sq_1_port_i_1), //i
    .port_i_2 (sq_1_port_i_2), //i
    .port_i_3 (sq_1_port_i_3), //i
    .port_o_0 (sq_1_port_o_0), //o
    .port_o_1 (sq_1_port_o_1), //o
    .port_o_2 (sq_1_port_o_2), //o
    .port_o_3 (sq_1_port_o_3)  //o
  );
  GF_MULS_4 gF_MULS_4_192 (
    .port_A_0   (port_a_0_0            ), //i
    .port_A_1   (port_a_0_1            ), //i
    .port_A_2   (port_a_0_2            ), //i
    .port_A_3   (port_a_0_3            ), //i
    .port_a_0_1 (sax_0_0               ), //i
    .port_a_1_1 (sax_0_1               ), //i
    .port_Al    (al_0                  ), //i
    .port_Ah    (ah_0                  ), //i
    .port_aa    (aa_0                  ), //i
    .port_B_0   (port_b_0_0            ), //i
    .port_B_1   (port_b_0_1            ), //i
    .port_B_2   (port_b_0_2            ), //i
    .port_B_3   (port_b_0_3            ), //i
    .port_b_0_1 (sbx_0_0               ), //i
    .port_b_1_1 (sbx_0_1               ), //i
    .port_Bl    (bl_0                  ), //i
    .port_Bh    (bh_0                  ), //i
    .port_bb    (bb_0                  ), //i
    .port_o_0   (gF_MULS_4_192_port_o_0), //o
    .port_o_1   (gF_MULS_4_192_port_o_1), //o
    .port_o_2   (gF_MULS_4_192_port_o_2), //o
    .port_o_3   (gF_MULS_4_192_port_o_3)  //o
  );
  GF_MULS_4 gF_MULS_4_193 (
    .port_A_0   (port_a_0_0            ), //i
    .port_A_1   (port_a_0_1            ), //i
    .port_A_2   (port_a_0_2            ), //i
    .port_A_3   (port_a_0_3            ), //i
    .port_a_0_1 (sax_0_0               ), //i
    .port_a_1_1 (sax_0_1               ), //i
    .port_Al    (al_0                  ), //i
    .port_Ah    (ah_0                  ), //i
    .port_aa    (aa_0                  ), //i
    .port_B_0   (port_b_1_0            ), //i
    .port_B_1   (port_b_1_1            ), //i
    .port_B_2   (port_b_1_2            ), //i
    .port_B_3   (port_b_1_3            ), //i
    .port_b_0_1 (sbx_1_0               ), //i
    .port_b_1_1 (sbx_1_1               ), //i
    .port_Bl    (bl_1                  ), //i
    .port_Bh    (bh_1                  ), //i
    .port_bb    (bb_1                  ), //i
    .port_o_0   (gF_MULS_4_193_port_o_0), //o
    .port_o_1   (gF_MULS_4_193_port_o_1), //o
    .port_o_2   (gF_MULS_4_193_port_o_2), //o
    .port_o_3   (gF_MULS_4_193_port_o_3)  //o
  );
  GF_MULS_4 gF_MULS_4_194 (
    .port_A_0   (port_a_1_0            ), //i
    .port_A_1   (port_a_1_1            ), //i
    .port_A_2   (port_a_1_2            ), //i
    .port_A_3   (port_a_1_3            ), //i
    .port_a_0_1 (sax_1_0               ), //i
    .port_a_1_1 (sax_1_1               ), //i
    .port_Al    (al_1                  ), //i
    .port_Ah    (ah_1                  ), //i
    .port_aa    (aa_1                  ), //i
    .port_B_0   (port_b_0_0            ), //i
    .port_B_1   (port_b_0_1            ), //i
    .port_B_2   (port_b_0_2            ), //i
    .port_B_3   (port_b_0_3            ), //i
    .port_b_0_1 (sbx_0_0               ), //i
    .port_b_1_1 (sbx_0_1               ), //i
    .port_Bl    (bl_0                  ), //i
    .port_Bh    (bh_0                  ), //i
    .port_bb    (bb_0                  ), //i
    .port_o_0   (gF_MULS_4_194_port_o_0), //o
    .port_o_1   (gF_MULS_4_194_port_o_1), //o
    .port_o_2   (gF_MULS_4_194_port_o_2), //o
    .port_o_3   (gF_MULS_4_194_port_o_3)  //o
  );
  GF_MULS_4 gF_MULS_4_195 (
    .port_A_0   (port_a_1_0            ), //i
    .port_A_1   (port_a_1_1            ), //i
    .port_A_2   (port_a_1_2            ), //i
    .port_A_3   (port_a_1_3            ), //i
    .port_a_0_1 (sax_1_0               ), //i
    .port_a_1_1 (sax_1_1               ), //i
    .port_Al    (al_1                  ), //i
    .port_Ah    (ah_1                  ), //i
    .port_aa    (aa_1                  ), //i
    .port_B_0   (port_b_1_0            ), //i
    .port_B_1   (port_b_1_1            ), //i
    .port_B_2   (port_b_1_2            ), //i
    .port_B_3   (port_b_1_3            ), //i
    .port_b_0_1 (sbx_1_0               ), //i
    .port_b_1_1 (sbx_1_1               ), //i
    .port_Bl    (bl_1                  ), //i
    .port_Bh    (bh_1                  ), //i
    .port_bb    (bb_1                  ), //i
    .port_o_0   (gF_MULS_4_195_port_o_0), //o
    .port_o_1   (gF_MULS_4_195_port_o_1), //o
    .port_o_2   (gF_MULS_4_195_port_o_2), //o
    .port_o_3   (gF_MULS_4_195_port_o_3)  //o
  );
  assign sq_0_port_i_0 = (port_a_0_0 ^ port_b_0_0);
  assign sq_0_port_i_1 = (port_a_0_1 ^ port_b_0_1);
  assign sq_0_port_i_2 = (port_a_0_2 ^ port_b_0_2);
  assign sq_0_port_i_3 = (port_a_0_3 ^ port_b_0_3);
  assign sq_0_0 = sq_0_port_o_0;
  assign sq_0_1 = sq_0_port_o_1;
  assign sq_0_2 = sq_0_port_o_2;
  assign sq_0_3 = sq_0_port_o_3;
  assign sq_1_port_i_0 = (port_a_1_0 ^ port_b_1_0);
  assign sq_1_port_i_1 = (port_a_1_1 ^ port_b_1_1);
  assign sq_1_port_i_2 = (port_a_1_2 ^ port_b_1_2);
  assign sq_1_port_i_3 = (port_a_1_3 ^ port_b_1_3);
  assign sq_1_0 = sq_1_port_o_0;
  assign sq_1_1 = sq_1_port_o_1;
  assign sq_1_2 = sq_1_port_o_2;
  assign sq_1_3 = sq_1_port_o_3;
  assign sax_0_0 = (port_a_0_2 ^ port_a_0_0);
  assign sax_0_1 = (port_a_0_3 ^ port_a_0_1);
  assign sbx_0_0 = (port_b_0_2 ^ port_b_0_0);
  assign sbx_0_1 = (port_b_0_3 ^ port_b_0_1);
  assign al_0 = (port_a_0_1 ^ port_a_0_0);
  assign ah_0 = (port_a_0_3 ^ port_a_0_2);
  assign aa_0 = (sax_0_1 ^ sax_0_0);
  assign bl_0 = (port_b_0_1 ^ port_b_0_0);
  assign bh_0 = (port_b_0_3 ^ port_b_0_2);
  assign bb_0 = (sbx_0_1 ^ sbx_0_0);
  assign sax_1_0 = (port_a_1_2 ^ port_a_1_0);
  assign sax_1_1 = (port_a_1_3 ^ port_a_1_1);
  assign sbx_1_0 = (port_b_1_2 ^ port_b_1_0);
  assign sbx_1_1 = (port_b_1_3 ^ port_b_1_1);
  assign al_1 = (port_a_1_1 ^ port_a_1_0);
  assign ah_1 = (port_a_1_3 ^ port_a_1_2);
  assign aa_1 = (sax_1_1 ^ sax_1_0);
  assign bl_1 = (port_b_1_1 ^ port_b_1_0);
  assign bh_1 = (port_b_1_3 ^ port_b_1_2);
  assign bb_1 = (sbx_1_1 ^ sbx_1_0);
  assign outVal_0_0 = (gF_MULS_4_192_port_o_0 ^ sq_0_0);
  assign outVal_0_1 = (gF_MULS_4_192_port_o_1 ^ sq_0_1);
  assign outVal_0_2 = (gF_MULS_4_192_port_o_2 ^ sq_0_2);
  assign outVal_0_3 = (gF_MULS_4_192_port_o_3 ^ sq_0_3);
  assign outVal_2_0 = gF_MULS_4_193_port_o_0;
  assign outVal_2_1 = gF_MULS_4_193_port_o_1;
  assign outVal_2_2 = gF_MULS_4_193_port_o_2;
  assign outVal_2_3 = gF_MULS_4_193_port_o_3;
  assign outVal_1_0 = gF_MULS_4_194_port_o_0;
  assign outVal_1_1 = gF_MULS_4_194_port_o_1;
  assign outVal_1_2 = gF_MULS_4_194_port_o_2;
  assign outVal_1_3 = gF_MULS_4_194_port_o_3;
  assign outVal_3_0 = (gF_MULS_4_195_port_o_0 ^ sq_1_0);
  assign outVal_3_1 = (gF_MULS_4_195_port_o_1 ^ sq_1_1);
  assign outVal_3_2 = (gF_MULS_4_195_port_o_2 ^ sq_1_2);
  assign outVal_3_3 = (gF_MULS_4_195_port_o_3 ^ sq_1_3);
  assign refVal_0_0[0] = (outVal_0_0[0] ^ port_r_0_0);
  assign refVal_0_1[0] = (outVal_0_1[0] ^ port_r_0_1);
  assign refVal_0_2[0] = (outVal_0_2[0] ^ port_r_0_2);
  assign refVal_0_3[0] = (outVal_0_3[0] ^ port_r_0_3);
  assign refVal_1_0[0] = (outVal_1_0[0] ^ port_r_1_0);
  assign refVal_1_1[0] = (outVal_1_1[0] ^ port_r_1_1);
  assign refVal_1_2[0] = (outVal_1_2[0] ^ port_r_1_2);
  assign refVal_1_3[0] = (outVal_1_3[0] ^ port_r_1_3);
  assign refVal_2_0[0] = (outVal_2_0[0] ^ port_r_2_0);
  assign refVal_2_1[0] = (outVal_2_1[0] ^ port_r_2_1);
  assign refVal_2_2[0] = (outVal_2_2[0] ^ port_r_2_2);
  assign refVal_2_3[0] = (outVal_2_3[0] ^ port_r_2_3);
  assign refVal_3_0[0] = (outVal_3_0[0] ^ ((port_r_0_0 ^ port_r_1_0) ^ port_r_2_0));
  assign refVal_3_1[0] = (outVal_3_1[0] ^ ((port_r_0_1 ^ port_r_1_1) ^ port_r_2_1));
  assign refVal_3_2[0] = (outVal_3_2[0] ^ ((port_r_0_2 ^ port_r_1_2) ^ port_r_2_2));
  assign refVal_3_3[0] = (outVal_3_3[0] ^ ((port_r_0_3 ^ port_r_1_3) ^ port_r_2_3));
  assign port_y_0_0 = outReg_0_0;
  assign port_y_0_1 = outReg_0_1;
  assign port_y_0_2 = outReg_0_2;
  assign port_y_0_3 = outReg_0_3;
  assign port_y_1_0 = outReg_1_0;
  assign port_y_1_1 = outReg_1_1;
  assign port_y_1_2 = outReg_1_2;
  assign port_y_1_3 = outReg_1_3;
  assign port_y_2_0 = outReg_2_0;
  assign port_y_2_1 = outReg_2_1;
  assign port_y_2_2 = outReg_2_2;
  assign port_y_2_3 = outReg_2_3;
  assign port_y_3_0 = outReg_3_0;
  assign port_y_3_1 = outReg_3_1;
  assign port_y_3_2 = outReg_3_2;
  assign port_y_3_3 = outReg_3_3;
  always @(posedge clk) begin
    outReg_0_0 <= refVal_0_0;
    outReg_0_1 <= refVal_0_1;
    outReg_0_2 <= refVal_0_2;
    outReg_0_3 <= refVal_0_3;
    outReg_1_0 <= refVal_1_0;
    outReg_1_1 <= refVal_1_1;
    outReg_1_2 <= refVal_1_2;
    outReg_1_3 <= refVal_1_3;
    outReg_2_0 <= refVal_2_0;
    outReg_2_1 <= refVal_2_1;
    outReg_2_2 <= refVal_2_2;
    outReg_2_3 <= refVal_2_3;
    outReg_3_0 <= refVal_3_0;
    outReg_3_1 <= refVal_3_1;
    outReg_3_2 <= refVal_3_2;
    outReg_3_3 <= refVal_3_3;
  end


endmodule

module CMS_stage1 (
  input      [0:0]    port_i_0_0,
  input      [0:0]    port_i_0_1,
  input      [0:0]    port_i_0_2,
  input      [0:0]    port_i_0_3,
  input      [0:0]    port_i_0_4,
  input      [0:0]    port_i_0_5,
  input      [0:0]    port_i_0_6,
  input      [0:0]    port_i_0_7,
  input      [0:0]    port_i_1_0,
  input      [0:0]    port_i_1_1,
  input      [0:0]    port_i_1_2,
  input      [0:0]    port_i_1_3,
  input      [0:0]    port_i_1_4,
  input      [0:0]    port_i_1_5,
  input      [0:0]    port_i_1_6,
  input      [0:0]    port_i_1_7,
  output     [0:0]    port_o_0_0,
  output     [0:0]    port_o_0_1,
  output     [0:0]    port_o_0_2,
  output     [0:0]    port_o_0_3,
  output     [0:0]    port_o_0_4,
  output     [0:0]    port_o_0_5,
  output     [0:0]    port_o_0_6,
  output     [0:0]    port_o_0_7,
  output     [0:0]    port_o_1_0,
  output     [0:0]    port_o_1_1,
  output     [0:0]    port_o_1_2,
  output     [0:0]    port_o_1_3,
  output     [0:0]    port_o_1_4,
  output     [0:0]    port_o_1_5,
  output     [0:0]    port_o_1_6,
  output     [0:0]    port_o_1_7,
  input               clk,
  input               reset
);

  reg        [0:0]    outReg_0_0;
  reg        [0:0]    outReg_0_1;
  reg        [0:0]    outReg_0_2;
  reg        [0:0]    outReg_0_3;
  reg        [0:0]    outReg_0_4;
  reg        [0:0]    outReg_0_5;
  reg        [0:0]    outReg_0_6;
  reg        [0:0]    outReg_0_7;
  reg        [0:0]    outReg_1_0;
  reg        [0:0]    outReg_1_1;
  reg        [0:0]    outReg_1_2;
  reg        [0:0]    outReg_1_3;
  reg        [0:0]    outReg_1_4;
  reg        [0:0]    outReg_1_5;
  reg        [0:0]    outReg_1_6;
  reg        [0:0]    outReg_1_7;
  wire       [0:0]    outVal_0_0;
  wire       [0:0]    outVal_0_1;
  wire       [0:0]    outVal_0_2;
  wire       [0:0]    outVal_0_3;
  wire       [0:0]    outVal_0_4;
  wire       [0:0]    outVal_0_5;
  wire       [0:0]    outVal_0_6;
  wire       [0:0]    outVal_0_7;
  wire       [0:0]    outVal_1_0;
  wire       [0:0]    outVal_1_1;
  wire       [0:0]    outVal_1_2;
  wire       [0:0]    outVal_1_3;
  wire       [0:0]    outVal_1_4;
  wire       [0:0]    outVal_1_5;
  wire       [0:0]    outVal_1_6;
  wire       [0:0]    outVal_1_7;
  wire       [0:0]    rx1_0;
  wire       [0:0]    rx2_0;
  wire       [0:0]    rx3_0;
  wire       [0:0]    rx4_0;
  wire       [0:0]    rx5_0;
  wire       [0:0]    rx6_0;
  wire       [0:0]    rx7_0;
  wire       [0:0]    rx8_0;
  wire       [0:0]    rx9_0;
  wire       [0:0]    rx1_1;
  wire       [0:0]    rx2_1;
  wire       [0:0]    rx3_1;
  wire       [0:0]    rx4_1;
  wire       [0:0]    rx5_1;
  wire       [0:0]    rx6_1;
  wire       [0:0]    rx7_1;
  wire       [0:0]    rx8_1;
  wire       [0:0]    rx9_1;

  assign rx1_0 = (port_i_0_7 ^ port_i_0_5);
  assign rx2_0 = (~ (port_i_0_7 ^ port_i_0_4));
  assign rx3_0 = (port_i_0_6 ^ port_i_0_0);
  assign rx4_0 = (~ (port_i_0_5 ^ rx3_0));
  assign rx5_0 = (port_i_0_4 ^ rx4_0);
  assign rx6_0 = (port_i_0_3 ^ port_i_0_0);
  assign rx7_0 = (port_i_0_2 ^ rx1_0);
  assign rx8_0 = (port_i_0_1 ^ rx3_0);
  assign rx9_0 = (port_i_0_3 ^ rx8_0);
  assign outVal_0_7 = (rx7_0 ^ rx8_0);
  assign outVal_0_6 = (~ rx5_0);
  assign outVal_0_5 = (~ (port_i_0_1 ^ rx4_0));
  assign outVal_0_4 = (rx1_0 ^ rx3_0);
  assign outVal_0_3 = (~ ((port_i_0_1 ^ rx2_0) ^ rx6_0));
  assign outVal_0_2 = port_i_0_0;
  assign outVal_0_1 = (~ rx4_0);
  assign outVal_0_0 = (port_i_0_2 ^ rx9_0);
  assign rx1_1 = (port_i_1_7 ^ port_i_1_5);
  assign rx2_1 = (port_i_1_7 ^ port_i_1_4);
  assign rx3_1 = (port_i_1_6 ^ port_i_1_0);
  assign rx4_1 = (port_i_1_5 ^ rx3_1);
  assign rx5_1 = (port_i_1_4 ^ rx4_1);
  assign rx6_1 = (port_i_1_3 ^ port_i_1_0);
  assign rx7_1 = (port_i_1_2 ^ rx1_1);
  assign rx8_1 = (port_i_1_1 ^ rx3_1);
  assign rx9_1 = (port_i_1_3 ^ rx8_1);
  assign outVal_1_7 = (rx7_1 ^ rx8_1);
  assign outVal_1_6 = rx5_1;
  assign outVal_1_5 = (port_i_1_1 ^ rx4_1);
  assign outVal_1_4 = (rx1_1 ^ rx3_1);
  assign outVal_1_3 = ((port_i_1_1 ^ rx2_1) ^ rx6_1);
  assign outVal_1_2 = port_i_1_0;
  assign outVal_1_1 = rx4_1;
  assign outVal_1_0 = (port_i_1_2 ^ rx9_1);
  assign port_o_0_0 = outReg_0_0;
  assign port_o_0_1 = outReg_0_1;
  assign port_o_0_2 = outReg_0_2;
  assign port_o_0_3 = outReg_0_3;
  assign port_o_0_4 = outReg_0_4;
  assign port_o_0_5 = outReg_0_5;
  assign port_o_0_6 = outReg_0_6;
  assign port_o_0_7 = outReg_0_7;
  assign port_o_1_0 = outReg_1_0;
  assign port_o_1_1 = outReg_1_1;
  assign port_o_1_2 = outReg_1_2;
  assign port_o_1_3 = outReg_1_3;
  assign port_o_1_4 = outReg_1_4;
  assign port_o_1_5 = outReg_1_5;
  assign port_o_1_6 = outReg_1_6;
  assign port_o_1_7 = outReg_1_7;
  always @(posedge clk) begin
    outReg_0_0 <= outVal_0_0;
    outReg_0_1 <= outVal_0_1;
    outReg_0_2 <= outVal_0_2;
    outReg_0_3 <= outVal_0_3;
    outReg_0_4 <= outVal_0_4;
    outReg_0_5 <= outVal_0_5;
    outReg_0_6 <= outVal_0_6;
    outReg_0_7 <= outVal_0_7;
    outReg_1_0 <= outVal_1_0;
    outReg_1_1 <= outVal_1_1;
    outReg_1_2 <= outVal_1_2;
    outReg_1_3 <= outVal_1_3;
    outReg_1_4 <= outVal_1_4;
    outReg_1_5 <= outVal_1_5;
    outReg_1_6 <= outVal_1_6;
    outReg_1_7 <= outVal_1_7;
  end


endmodule

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_SCLW2_2 replaced by GF_SCLW2_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_SCLW2_2 replaced by GF_SCLW2_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_SQ_SCL_4 replaced by GF_SQ_SCL_4

//GF_SQ_SCL_4 replaced by GF_SQ_SCL_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_SCLW2_2 replaced by GF_SCLW2_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_SCLW2_2 replaced by GF_SCLW2_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_SQ_SCL_4 replaced by GF_SQ_SCL_4

//GF_SQ_SCL_4 replaced by GF_SQ_SCL_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_SCLW2_2 replaced by GF_SCLW2_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_SCLW2_2 replaced by GF_SCLW2_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_SQ_SCL_4 replaced by GF_SQ_SCL_4

//GF_SQ_SCL_4 replaced by GF_SQ_SCL_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_SCLW2_2 replaced by GF_SCLW2_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_SCLW2_2 replaced by GF_SCLW2_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_SQ_SCL_4 replaced by GF_SQ_SCL_4

//GF_SQ_SCL_4 replaced by GF_SQ_SCL_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_SCLW2_2 replaced by GF_SCLW2_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_SCLW2_2 replaced by GF_SCLW2_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_SQ_SCL_4 replaced by GF_SQ_SCL_4

//GF_SQ_SCL_4 replaced by GF_SQ_SCL_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_SCLW2_2 replaced by GF_SCLW2_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_SCLW2_2 replaced by GF_SCLW2_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_SQ_SCL_4 replaced by GF_SQ_SCL_4

//GF_SQ_SCL_4 replaced by GF_SQ_SCL_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_SCLW2_2 replaced by GF_SCLW2_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_SCLW2_2 replaced by GF_SCLW2_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_SQ_SCL_4 replaced by GF_SQ_SCL_4

//GF_SQ_SCL_4 replaced by GF_SQ_SCL_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_SCLW2_2 replaced by GF_SCLW2_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_SCLW2_2 replaced by GF_SCLW2_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_SQ_SCL_4 replaced by GF_SQ_SCL_4

//GF_SQ_SCL_4 replaced by GF_SQ_SCL_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_SCLW2_2 replaced by GF_SCLW2_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_SCLW2_2 replaced by GF_SCLW2_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_SQ_SCL_4 replaced by GF_SQ_SCL_4

//GF_SQ_SCL_4 replaced by GF_SQ_SCL_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_SCLW2_2 replaced by GF_SCLW2_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_SCLW2_2 replaced by GF_SCLW2_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_SQ_SCL_4 replaced by GF_SQ_SCL_4

//GF_SQ_SCL_4 replaced by GF_SQ_SCL_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_SCLW2_2 replaced by GF_SCLW2_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_SCLW2_2 replaced by GF_SCLW2_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_SQ_SCL_4 replaced by GF_SQ_SCL_4

//GF_SQ_SCL_4 replaced by GF_SQ_SCL_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_SCLW2_2 replaced by GF_SCLW2_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_SCLW2_2 replaced by GF_SCLW2_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_SQ_SCL_4 replaced by GF_SQ_SCL_4

//GF_SQ_SCL_4 replaced by GF_SQ_SCL_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_SCLW2_2 replaced by GF_SCLW2_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_SCLW2_2 replaced by GF_SCLW2_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_SQ_SCL_4 replaced by GF_SQ_SCL_4

//GF_SQ_SCL_4 replaced by GF_SQ_SCL_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_SCLW2_2 replaced by GF_SCLW2_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_SCLW2_2 replaced by GF_SCLW2_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_SQ_SCL_4 replaced by GF_SQ_SCL_4

//GF_SQ_SCL_4 replaced by GF_SQ_SCL_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_SCLW2_2 replaced by GF_SCLW2_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_SCLW2_2 replaced by GF_SCLW2_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_SQ_SCL_4 replaced by GF_SQ_SCL_4

//GF_SQ_SCL_4 replaced by GF_SQ_SCL_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_SCLW2_2 replaced by GF_SCLW2_2

//GF_SQ_2 replaced by GF_SQ_2

module GF_SCLW2_2 (
  input      [0:0]    port_i_0,
  input      [0:0]    port_i_1,
  output     [0:0]    port_o_0,
  output     [0:0]    port_o_1
);


  assign port_o_0 = (port_i_1 ^ port_i_0);
  assign port_o_1 = port_i_0;

endmodule

//GF_SQ_2 replaced by GF_SQ_2

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

//GF_MULS_4 replaced by GF_MULS_4

module GF_MULS_4 (
  input      [0:0]    port_A_0,
  input      [0:0]    port_A_1,
  input      [0:0]    port_A_2,
  input      [0:0]    port_A_3,
  input      [0:0]    port_a_0_1,
  input      [0:0]    port_a_1_1,
  input      [0:0]    port_Al,
  input      [0:0]    port_Ah,
  input      [0:0]    port_aa,
  input      [0:0]    port_B_0,
  input      [0:0]    port_B_1,
  input      [0:0]    port_B_2,
  input      [0:0]    port_B_3,
  input      [0:0]    port_b_0_1,
  input      [0:0]    port_b_1_1,
  input      [0:0]    port_Bl,
  input      [0:0]    port_Bh,
  input      [0:0]    port_bb,
  output     [0:0]    port_o_0,
  output     [0:0]    port_o_1,
  output     [0:0]    port_o_2,
  output     [0:0]    port_o_3
);

  wire       [0:0]    hi_mul_port_o_0;
  wire       [0:0]    hi_mul_port_o_1;
  wire       [0:0]    lo_mul_port_o_0;
  wire       [0:0]    lo_mul_port_o_1;
  wire       [0:0]    sum_mul_port_o_0;
  wire       [0:0]    sum_mul_port_o_1;
  wire       [0:0]    ph_0;
  wire       [0:0]    ph_1;
  wire       [0:0]    pl_0;
  wire       [0:0]    pl_1;
  wire       [0:0]    p_0;
  wire       [0:0]    p_1;

  GF_MULS_2 hi_mul (
    .port_a_0 (port_A_2       ), //i
    .port_a_1 (port_A_3       ), //i
    .port_ab  (port_Ah        ), //i
    .port_b_0 (port_B_2       ), //i
    .port_b_1 (port_B_3       ), //i
    .port_cd  (port_Bh        ), //i
    .port_o_0 (hi_mul_port_o_0), //o
    .port_o_1 (hi_mul_port_o_1)  //o
  );
  GF_MULS_2 lo_mul (
    .port_a_0 (port_A_0       ), //i
    .port_a_1 (port_A_1       ), //i
    .port_ab  (port_Al        ), //i
    .port_b_0 (port_B_0       ), //i
    .port_b_1 (port_B_1       ), //i
    .port_cd  (port_Bl        ), //i
    .port_o_0 (lo_mul_port_o_0), //o
    .port_o_1 (lo_mul_port_o_1)  //o
  );
  GF_MULS_SCL_2 sum_mul (
    .port_a_0 (port_a_0_1      ), //i
    .port_a_1 (port_a_1_1      ), //i
    .port_ab  (port_aa         ), //i
    .port_b_0 (port_b_0_1      ), //i
    .port_b_1 (port_b_1_1      ), //i
    .port_cd  (port_bb         ), //i
    .port_o_0 (sum_mul_port_o_0), //o
    .port_o_1 (sum_mul_port_o_1)  //o
  );
  assign ph_0 = hi_mul_port_o_0;
  assign ph_1 = hi_mul_port_o_1;
  assign pl_0 = lo_mul_port_o_0;
  assign pl_1 = lo_mul_port_o_1;
  assign p_0 = sum_mul_port_o_0;
  assign p_1 = sum_mul_port_o_1;
  assign port_o_0 = (pl_0 ^ p_0);
  assign port_o_1 = (pl_1 ^ p_1);
  assign port_o_2 = (ph_0 ^ p_0);
  assign port_o_3 = (ph_1 ^ p_1);

endmodule

//GF_SQ_SCL_4 replaced by GF_SQ_SCL_4

module GF_SQ_SCL_4 (
  input      [0:0]    port_i_0,
  input      [0:0]    port_i_1,
  input      [0:0]    port_i_2,
  input      [0:0]    port_i_3,
  output     [0:0]    port_o_0,
  output     [0:0]    port_o_1,
  output     [0:0]    port_o_2,
  output     [0:0]    port_o_3
);

  wire       [0:0]    ab_sq_port_o_0;
  wire       [0:0]    ab_sq_port_o_1;
  wire       [0:0]    b_sq_port_o_0;
  wire       [0:0]    b_sq_port_o_1;
  wire       [0:0]    b_mulN2_port_o_0;
  wire       [0:0]    b_mulN2_port_o_1;
  wire       [0:0]    ax_0;
  wire       [0:0]    ax_1;
  wire       [0:0]    bx_0;
  wire       [0:0]    bx_1;
  wire       [0:0]    abx_0;
  wire       [0:0]    abx_1;
  wire       [0:0]    ab2x_0;
  wire       [0:0]    ab2x_1;
  wire       [0:0]    b2x_0;
  wire       [0:0]    b2x_1;
  wire       [0:0]    b2N2_0;
  wire       [0:0]    b2N2_1;

  GF_SQ_2 ab_sq (
    .port_i_0 (abx_0         ), //i
    .port_i_1 (abx_1         ), //i
    .port_o_0 (ab_sq_port_o_0), //o
    .port_o_1 (ab_sq_port_o_1)  //o
  );
  GF_SQ_2 b_sq (
    .port_i_0 (bx_0         ), //i
    .port_i_1 (bx_1         ), //i
    .port_o_0 (b_sq_port_o_0), //o
    .port_o_1 (b_sq_port_o_1)  //o
  );
  GF_SCLW_2 b_mulN2 (
    .port_i_0 (b2x_0           ), //i
    .port_i_1 (b2x_1           ), //i
    .port_o_0 (b_mulN2_port_o_0), //o
    .port_o_1 (b_mulN2_port_o_1)  //o
  );
  assign ax_0 = port_i_2;
  assign ax_1 = port_i_3;
  assign bx_0 = port_i_0;
  assign bx_1 = port_i_1;
  assign abx_0 = (ax_0 ^ bx_0);
  assign abx_1 = (ax_1 ^ bx_1);
  assign ab2x_0 = ab_sq_port_o_0;
  assign ab2x_1 = ab_sq_port_o_1;
  assign b2x_0 = b_sq_port_o_0;
  assign b2x_1 = b_sq_port_o_1;
  assign b2N2_0 = b_mulN2_port_o_0;
  assign b2N2_1 = b_mulN2_port_o_1;
  assign port_o_0 = b2N2_0;
  assign port_o_1 = b2N2_1;
  assign port_o_2 = ab2x_0;
  assign port_o_3 = ab2x_1;

endmodule

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_SCLW_2 replaced by GF_SCLW_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_SCLW_2 replaced by GF_SCLW_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_SCLW_2 replaced by GF_SCLW_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_SCLW_2 replaced by GF_SCLW_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_SCLW_2 replaced by GF_SCLW_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_SCLW_2 replaced by GF_SCLW_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_SCLW_2 replaced by GF_SCLW_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_SCLW_2 replaced by GF_SCLW_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_SCLW_2 replaced by GF_SCLW_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_SCLW_2 replaced by GF_SCLW_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_SCLW_2 replaced by GF_SCLW_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_SCLW_2 replaced by GF_SCLW_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_SCLW_2 replaced by GF_SCLW_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_SCLW_2 replaced by GF_SCLW_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_SCLW_2 replaced by GF_SCLW_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_SCLW_2 replaced by GF_SCLW_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_SCLW_2 replaced by GF_SCLW_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_SCLW_2 replaced by GF_SCLW_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_SCLW_2 replaced by GF_SCLW_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_SCLW_2 replaced by GF_SCLW_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_SCLW_2 replaced by GF_SCLW_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_SCLW_2 replaced by GF_SCLW_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_SCLW_2 replaced by GF_SCLW_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_SCLW_2 replaced by GF_SCLW_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_SCLW_2 replaced by GF_SCLW_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_SCLW_2 replaced by GF_SCLW_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_SCLW_2 replaced by GF_SCLW_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_SCLW_2 replaced by GF_SCLW_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_SCLW_2 replaced by GF_SCLW_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_SCLW_2 replaced by GF_SCLW_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_SCL_2 replaced by GF_MULS_SCL_2

//GF_MULS_2 replaced by GF_MULS_2

//GF_MULS_2 replaced by GF_MULS_2

module GF_MULS_SCL_2 (
  input      [0:0]    port_a_0,
  input      [0:0]    port_a_1,
  input      [0:0]    port_ab,
  input      [0:0]    port_b_0,
  input      [0:0]    port_b_1,
  input      [0:0]    port_cd,
  output     [0:0]    port_o_0,
  output     [0:0]    port_o_1
);

  wire       [0:0]    t;

  assign t = (~ (port_a_0 & port_b_0));
  assign port_o_0 = ((~ (port_a_1 & port_b_1)) ^ t);
  assign port_o_1 = ((~ (port_ab & port_cd)) ^ t);

endmodule

//GF_MULS_2 replaced by GF_MULS_2

module GF_MULS_2 (
  input      [0:0]    port_a_0,
  input      [0:0]    port_a_1,
  input      [0:0]    port_ab,
  input      [0:0]    port_b_0,
  input      [0:0]    port_b_1,
  input      [0:0]    port_cd,
  output     [0:0]    port_o_0,
  output     [0:0]    port_o_1
);

  wire       [0:0]    t;

  assign t = (~ (port_ab & port_cd));
  assign port_o_0 = ((~ (port_a_0 & port_b_0)) ^ t);
  assign port_o_1 = ((~ (port_a_1 & port_b_1)) ^ t);

endmodule

//GF_SCLW_2 replaced by GF_SCLW_2

//GF_SQ_2 replaced by GF_SQ_2

//GF_SQ_2 replaced by GF_SQ_2

module GF_SCLW_2 (
  input      [0:0]    port_i_0,
  input      [0:0]    port_i_1,
  output     [0:0]    port_o_0,
  output     [0:0]    port_o_1
);


  assign port_o_0 = port_i_1;
  assign port_o_1 = (port_i_0 ^ port_i_1);

endmodule

//GF_SQ_2 replaced by GF_SQ_2

module GF_SQ_2 (
  input      [0:0]    port_i_0,
  input      [0:0]    port_i_1,
  output     [0:0]    port_o_0,
  output     [0:0]    port_o_1
);


  assign port_o_0 = port_i_1;
  assign port_o_1 = port_i_0;

endmodule
