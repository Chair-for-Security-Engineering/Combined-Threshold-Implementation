// Generator : SpinalHDL v1.7.3    git head : aeaeece704fe43c766e0d36a93f2ecbb8a9f2003
// Component : AES_Round
// Git hash  : db593c14fe8e83f0a4a5d43cf13325e631d65148

`timescale 1ns/1ps

module Round_AES_CTI_d1_k1 (
  input      [2:0]    port_state_in_0_0_0,
  input      [2:0]    port_state_in_0_0_1,
  input      [2:0]    port_state_in_0_0_2,
  input      [2:0]    port_state_in_0_0_3,
  input      [2:0]    port_state_in_0_0_4,
  input      [2:0]    port_state_in_0_0_5,
  input      [2:0]    port_state_in_0_0_6,
  input      [2:0]    port_state_in_0_0_7,
  input      [2:0]    port_state_in_0_1_0,
  input      [2:0]    port_state_in_0_1_1,
  input      [2:0]    port_state_in_0_1_2,
  input      [2:0]    port_state_in_0_1_3,
  input      [2:0]    port_state_in_0_1_4,
  input      [2:0]    port_state_in_0_1_5,
  input      [2:0]    port_state_in_0_1_6,
  input      [2:0]    port_state_in_0_1_7,
  input      [2:0]    port_state_in_0_2_0,
  input      [2:0]    port_state_in_0_2_1,
  input      [2:0]    port_state_in_0_2_2,
  input      [2:0]    port_state_in_0_2_3,
  input      [2:0]    port_state_in_0_2_4,
  input      [2:0]    port_state_in_0_2_5,
  input      [2:0]    port_state_in_0_2_6,
  input      [2:0]    port_state_in_0_2_7,
  input      [2:0]    port_state_in_0_3_0,
  input      [2:0]    port_state_in_0_3_1,
  input      [2:0]    port_state_in_0_3_2,
  input      [2:0]    port_state_in_0_3_3,
  input      [2:0]    port_state_in_0_3_4,
  input      [2:0]    port_state_in_0_3_5,
  input      [2:0]    port_state_in_0_3_6,
  input      [2:0]    port_state_in_0_3_7,
  input      [2:0]    port_state_in_1_0_0,
  input      [2:0]    port_state_in_1_0_1,
  input      [2:0]    port_state_in_1_0_2,
  input      [2:0]    port_state_in_1_0_3,
  input      [2:0]    port_state_in_1_0_4,
  input      [2:0]    port_state_in_1_0_5,
  input      [2:0]    port_state_in_1_0_6,
  input      [2:0]    port_state_in_1_0_7,
  input      [2:0]    port_state_in_1_1_0,
  input      [2:0]    port_state_in_1_1_1,
  input      [2:0]    port_state_in_1_1_2,
  input      [2:0]    port_state_in_1_1_3,
  input      [2:0]    port_state_in_1_1_4,
  input      [2:0]    port_state_in_1_1_5,
  input      [2:0]    port_state_in_1_1_6,
  input      [2:0]    port_state_in_1_1_7,
  input      [2:0]    port_state_in_1_2_0,
  input      [2:0]    port_state_in_1_2_1,
  input      [2:0]    port_state_in_1_2_2,
  input      [2:0]    port_state_in_1_2_3,
  input      [2:0]    port_state_in_1_2_4,
  input      [2:0]    port_state_in_1_2_5,
  input      [2:0]    port_state_in_1_2_6,
  input      [2:0]    port_state_in_1_2_7,
  input      [2:0]    port_state_in_1_3_0,
  input      [2:0]    port_state_in_1_3_1,
  input      [2:0]    port_state_in_1_3_2,
  input      [2:0]    port_state_in_1_3_3,
  input      [2:0]    port_state_in_1_3_4,
  input      [2:0]    port_state_in_1_3_5,
  input      [2:0]    port_state_in_1_3_6,
  input      [2:0]    port_state_in_1_3_7,
  input      [2:0]    port_state_in_2_0_0,
  input      [2:0]    port_state_in_2_0_1,
  input      [2:0]    port_state_in_2_0_2,
  input      [2:0]    port_state_in_2_0_3,
  input      [2:0]    port_state_in_2_0_4,
  input      [2:0]    port_state_in_2_0_5,
  input      [2:0]    port_state_in_2_0_6,
  input      [2:0]    port_state_in_2_0_7,
  input      [2:0]    port_state_in_2_1_0,
  input      [2:0]    port_state_in_2_1_1,
  input      [2:0]    port_state_in_2_1_2,
  input      [2:0]    port_state_in_2_1_3,
  input      [2:0]    port_state_in_2_1_4,
  input      [2:0]    port_state_in_2_1_5,
  input      [2:0]    port_state_in_2_1_6,
  input      [2:0]    port_state_in_2_1_7,
  input      [2:0]    port_state_in_2_2_0,
  input      [2:0]    port_state_in_2_2_1,
  input      [2:0]    port_state_in_2_2_2,
  input      [2:0]    port_state_in_2_2_3,
  input      [2:0]    port_state_in_2_2_4,
  input      [2:0]    port_state_in_2_2_5,
  input      [2:0]    port_state_in_2_2_6,
  input      [2:0]    port_state_in_2_2_7,
  input      [2:0]    port_state_in_2_3_0,
  input      [2:0]    port_state_in_2_3_1,
  input      [2:0]    port_state_in_2_3_2,
  input      [2:0]    port_state_in_2_3_3,
  input      [2:0]    port_state_in_2_3_4,
  input      [2:0]    port_state_in_2_3_5,
  input      [2:0]    port_state_in_2_3_6,
  input      [2:0]    port_state_in_2_3_7,
  input      [2:0]    port_state_in_3_0_0,
  input      [2:0]    port_state_in_3_0_1,
  input      [2:0]    port_state_in_3_0_2,
  input      [2:0]    port_state_in_3_0_3,
  input      [2:0]    port_state_in_3_0_4,
  input      [2:0]    port_state_in_3_0_5,
  input      [2:0]    port_state_in_3_0_6,
  input      [2:0]    port_state_in_3_0_7,
  input      [2:0]    port_state_in_3_1_0,
  input      [2:0]    port_state_in_3_1_1,
  input      [2:0]    port_state_in_3_1_2,
  input      [2:0]    port_state_in_3_1_3,
  input      [2:0]    port_state_in_3_1_4,
  input      [2:0]    port_state_in_3_1_5,
  input      [2:0]    port_state_in_3_1_6,
  input      [2:0]    port_state_in_3_1_7,
  input      [2:0]    port_state_in_3_2_0,
  input      [2:0]    port_state_in_3_2_1,
  input      [2:0]    port_state_in_3_2_2,
  input      [2:0]    port_state_in_3_2_3,
  input      [2:0]    port_state_in_3_2_4,
  input      [2:0]    port_state_in_3_2_5,
  input      [2:0]    port_state_in_3_2_6,
  input      [2:0]    port_state_in_3_2_7,
  input      [2:0]    port_state_in_3_3_0,
  input      [2:0]    port_state_in_3_3_1,
  input      [2:0]    port_state_in_3_3_2,
  input      [2:0]    port_state_in_3_3_3,
  input      [2:0]    port_state_in_3_3_4,
  input      [2:0]    port_state_in_3_3_5,
  input      [2:0]    port_state_in_3_3_6,
  input      [2:0]    port_state_in_3_3_7,
  input      [2:0]    port_state_in_4_0_0,
  input      [2:0]    port_state_in_4_0_1,
  input      [2:0]    port_state_in_4_0_2,
  input      [2:0]    port_state_in_4_0_3,
  input      [2:0]    port_state_in_4_0_4,
  input      [2:0]    port_state_in_4_0_5,
  input      [2:0]    port_state_in_4_0_6,
  input      [2:0]    port_state_in_4_0_7,
  input      [2:0]    port_state_in_4_1_0,
  input      [2:0]    port_state_in_4_1_1,
  input      [2:0]    port_state_in_4_1_2,
  input      [2:0]    port_state_in_4_1_3,
  input      [2:0]    port_state_in_4_1_4,
  input      [2:0]    port_state_in_4_1_5,
  input      [2:0]    port_state_in_4_1_6,
  input      [2:0]    port_state_in_4_1_7,
  input      [2:0]    port_state_in_4_2_0,
  input      [2:0]    port_state_in_4_2_1,
  input      [2:0]    port_state_in_4_2_2,
  input      [2:0]    port_state_in_4_2_3,
  input      [2:0]    port_state_in_4_2_4,
  input      [2:0]    port_state_in_4_2_5,
  input      [2:0]    port_state_in_4_2_6,
  input      [2:0]    port_state_in_4_2_7,
  input      [2:0]    port_state_in_4_3_0,
  input      [2:0]    port_state_in_4_3_1,
  input      [2:0]    port_state_in_4_3_2,
  input      [2:0]    port_state_in_4_3_3,
  input      [2:0]    port_state_in_4_3_4,
  input      [2:0]    port_state_in_4_3_5,
  input      [2:0]    port_state_in_4_3_6,
  input      [2:0]    port_state_in_4_3_7,
  input      [2:0]    port_state_in_5_0_0,
  input      [2:0]    port_state_in_5_0_1,
  input      [2:0]    port_state_in_5_0_2,
  input      [2:0]    port_state_in_5_0_3,
  input      [2:0]    port_state_in_5_0_4,
  input      [2:0]    port_state_in_5_0_5,
  input      [2:0]    port_state_in_5_0_6,
  input      [2:0]    port_state_in_5_0_7,
  input      [2:0]    port_state_in_5_1_0,
  input      [2:0]    port_state_in_5_1_1,
  input      [2:0]    port_state_in_5_1_2,
  input      [2:0]    port_state_in_5_1_3,
  input      [2:0]    port_state_in_5_1_4,
  input      [2:0]    port_state_in_5_1_5,
  input      [2:0]    port_state_in_5_1_6,
  input      [2:0]    port_state_in_5_1_7,
  input      [2:0]    port_state_in_5_2_0,
  input      [2:0]    port_state_in_5_2_1,
  input      [2:0]    port_state_in_5_2_2,
  input      [2:0]    port_state_in_5_2_3,
  input      [2:0]    port_state_in_5_2_4,
  input      [2:0]    port_state_in_5_2_5,
  input      [2:0]    port_state_in_5_2_6,
  input      [2:0]    port_state_in_5_2_7,
  input      [2:0]    port_state_in_5_3_0,
  input      [2:0]    port_state_in_5_3_1,
  input      [2:0]    port_state_in_5_3_2,
  input      [2:0]    port_state_in_5_3_3,
  input      [2:0]    port_state_in_5_3_4,
  input      [2:0]    port_state_in_5_3_5,
  input      [2:0]    port_state_in_5_3_6,
  input      [2:0]    port_state_in_5_3_7,
  input      [2:0]    port_state_in_6_0_0,
  input      [2:0]    port_state_in_6_0_1,
  input      [2:0]    port_state_in_6_0_2,
  input      [2:0]    port_state_in_6_0_3,
  input      [2:0]    port_state_in_6_0_4,
  input      [2:0]    port_state_in_6_0_5,
  input      [2:0]    port_state_in_6_0_6,
  input      [2:0]    port_state_in_6_0_7,
  input      [2:0]    port_state_in_6_1_0,
  input      [2:0]    port_state_in_6_1_1,
  input      [2:0]    port_state_in_6_1_2,
  input      [2:0]    port_state_in_6_1_3,
  input      [2:0]    port_state_in_6_1_4,
  input      [2:0]    port_state_in_6_1_5,
  input      [2:0]    port_state_in_6_1_6,
  input      [2:0]    port_state_in_6_1_7,
  input      [2:0]    port_state_in_6_2_0,
  input      [2:0]    port_state_in_6_2_1,
  input      [2:0]    port_state_in_6_2_2,
  input      [2:0]    port_state_in_6_2_3,
  input      [2:0]    port_state_in_6_2_4,
  input      [2:0]    port_state_in_6_2_5,
  input      [2:0]    port_state_in_6_2_6,
  input      [2:0]    port_state_in_6_2_7,
  input      [2:0]    port_state_in_6_3_0,
  input      [2:0]    port_state_in_6_3_1,
  input      [2:0]    port_state_in_6_3_2,
  input      [2:0]    port_state_in_6_3_3,
  input      [2:0]    port_state_in_6_3_4,
  input      [2:0]    port_state_in_6_3_5,
  input      [2:0]    port_state_in_6_3_6,
  input      [2:0]    port_state_in_6_3_7,
  input      [2:0]    port_state_in_7_0_0,
  input      [2:0]    port_state_in_7_0_1,
  input      [2:0]    port_state_in_7_0_2,
  input      [2:0]    port_state_in_7_0_3,
  input      [2:0]    port_state_in_7_0_4,
  input      [2:0]    port_state_in_7_0_5,
  input      [2:0]    port_state_in_7_0_6,
  input      [2:0]    port_state_in_7_0_7,
  input      [2:0]    port_state_in_7_1_0,
  input      [2:0]    port_state_in_7_1_1,
  input      [2:0]    port_state_in_7_1_2,
  input      [2:0]    port_state_in_7_1_3,
  input      [2:0]    port_state_in_7_1_4,
  input      [2:0]    port_state_in_7_1_5,
  input      [2:0]    port_state_in_7_1_6,
  input      [2:0]    port_state_in_7_1_7,
  input      [2:0]    port_state_in_7_2_0,
  input      [2:0]    port_state_in_7_2_1,
  input      [2:0]    port_state_in_7_2_2,
  input      [2:0]    port_state_in_7_2_3,
  input      [2:0]    port_state_in_7_2_4,
  input      [2:0]    port_state_in_7_2_5,
  input      [2:0]    port_state_in_7_2_6,
  input      [2:0]    port_state_in_7_2_7,
  input      [2:0]    port_state_in_7_3_0,
  input      [2:0]    port_state_in_7_3_1,
  input      [2:0]    port_state_in_7_3_2,
  input      [2:0]    port_state_in_7_3_3,
  input      [2:0]    port_state_in_7_3_4,
  input      [2:0]    port_state_in_7_3_5,
  input      [2:0]    port_state_in_7_3_6,
  input      [2:0]    port_state_in_7_3_7,
  input      [2:0]    port_state_in_8_0_0,
  input      [2:0]    port_state_in_8_0_1,
  input      [2:0]    port_state_in_8_0_2,
  input      [2:0]    port_state_in_8_0_3,
  input      [2:0]    port_state_in_8_0_4,
  input      [2:0]    port_state_in_8_0_5,
  input      [2:0]    port_state_in_8_0_6,
  input      [2:0]    port_state_in_8_0_7,
  input      [2:0]    port_state_in_8_1_0,
  input      [2:0]    port_state_in_8_1_1,
  input      [2:0]    port_state_in_8_1_2,
  input      [2:0]    port_state_in_8_1_3,
  input      [2:0]    port_state_in_8_1_4,
  input      [2:0]    port_state_in_8_1_5,
  input      [2:0]    port_state_in_8_1_6,
  input      [2:0]    port_state_in_8_1_7,
  input      [2:0]    port_state_in_8_2_0,
  input      [2:0]    port_state_in_8_2_1,
  input      [2:0]    port_state_in_8_2_2,
  input      [2:0]    port_state_in_8_2_3,
  input      [2:0]    port_state_in_8_2_4,
  input      [2:0]    port_state_in_8_2_5,
  input      [2:0]    port_state_in_8_2_6,
  input      [2:0]    port_state_in_8_2_7,
  input      [2:0]    port_state_in_8_3_0,
  input      [2:0]    port_state_in_8_3_1,
  input      [2:0]    port_state_in_8_3_2,
  input      [2:0]    port_state_in_8_3_3,
  input      [2:0]    port_state_in_8_3_4,
  input      [2:0]    port_state_in_8_3_5,
  input      [2:0]    port_state_in_8_3_6,
  input      [2:0]    port_state_in_8_3_7,
  input      [2:0]    port_state_in_9_0_0,
  input      [2:0]    port_state_in_9_0_1,
  input      [2:0]    port_state_in_9_0_2,
  input      [2:0]    port_state_in_9_0_3,
  input      [2:0]    port_state_in_9_0_4,
  input      [2:0]    port_state_in_9_0_5,
  input      [2:0]    port_state_in_9_0_6,
  input      [2:0]    port_state_in_9_0_7,
  input      [2:0]    port_state_in_9_1_0,
  input      [2:0]    port_state_in_9_1_1,
  input      [2:0]    port_state_in_9_1_2,
  input      [2:0]    port_state_in_9_1_3,
  input      [2:0]    port_state_in_9_1_4,
  input      [2:0]    port_state_in_9_1_5,
  input      [2:0]    port_state_in_9_1_6,
  input      [2:0]    port_state_in_9_1_7,
  input      [2:0]    port_state_in_9_2_0,
  input      [2:0]    port_state_in_9_2_1,
  input      [2:0]    port_state_in_9_2_2,
  input      [2:0]    port_state_in_9_2_3,
  input      [2:0]    port_state_in_9_2_4,
  input      [2:0]    port_state_in_9_2_5,
  input      [2:0]    port_state_in_9_2_6,
  input      [2:0]    port_state_in_9_2_7,
  input      [2:0]    port_state_in_9_3_0,
  input      [2:0]    port_state_in_9_3_1,
  input      [2:0]    port_state_in_9_3_2,
  input      [2:0]    port_state_in_9_3_3,
  input      [2:0]    port_state_in_9_3_4,
  input      [2:0]    port_state_in_9_3_5,
  input      [2:0]    port_state_in_9_3_6,
  input      [2:0]    port_state_in_9_3_7,
  input      [2:0]    port_state_in_10_0_0,
  input      [2:0]    port_state_in_10_0_1,
  input      [2:0]    port_state_in_10_0_2,
  input      [2:0]    port_state_in_10_0_3,
  input      [2:0]    port_state_in_10_0_4,
  input      [2:0]    port_state_in_10_0_5,
  input      [2:0]    port_state_in_10_0_6,
  input      [2:0]    port_state_in_10_0_7,
  input      [2:0]    port_state_in_10_1_0,
  input      [2:0]    port_state_in_10_1_1,
  input      [2:0]    port_state_in_10_1_2,
  input      [2:0]    port_state_in_10_1_3,
  input      [2:0]    port_state_in_10_1_4,
  input      [2:0]    port_state_in_10_1_5,
  input      [2:0]    port_state_in_10_1_6,
  input      [2:0]    port_state_in_10_1_7,
  input      [2:0]    port_state_in_10_2_0,
  input      [2:0]    port_state_in_10_2_1,
  input      [2:0]    port_state_in_10_2_2,
  input      [2:0]    port_state_in_10_2_3,
  input      [2:0]    port_state_in_10_2_4,
  input      [2:0]    port_state_in_10_2_5,
  input      [2:0]    port_state_in_10_2_6,
  input      [2:0]    port_state_in_10_2_7,
  input      [2:0]    port_state_in_10_3_0,
  input      [2:0]    port_state_in_10_3_1,
  input      [2:0]    port_state_in_10_3_2,
  input      [2:0]    port_state_in_10_3_3,
  input      [2:0]    port_state_in_10_3_4,
  input      [2:0]    port_state_in_10_3_5,
  input      [2:0]    port_state_in_10_3_6,
  input      [2:0]    port_state_in_10_3_7,
  input      [2:0]    port_state_in_11_0_0,
  input      [2:0]    port_state_in_11_0_1,
  input      [2:0]    port_state_in_11_0_2,
  input      [2:0]    port_state_in_11_0_3,
  input      [2:0]    port_state_in_11_0_4,
  input      [2:0]    port_state_in_11_0_5,
  input      [2:0]    port_state_in_11_0_6,
  input      [2:0]    port_state_in_11_0_7,
  input      [2:0]    port_state_in_11_1_0,
  input      [2:0]    port_state_in_11_1_1,
  input      [2:0]    port_state_in_11_1_2,
  input      [2:0]    port_state_in_11_1_3,
  input      [2:0]    port_state_in_11_1_4,
  input      [2:0]    port_state_in_11_1_5,
  input      [2:0]    port_state_in_11_1_6,
  input      [2:0]    port_state_in_11_1_7,
  input      [2:0]    port_state_in_11_2_0,
  input      [2:0]    port_state_in_11_2_1,
  input      [2:0]    port_state_in_11_2_2,
  input      [2:0]    port_state_in_11_2_3,
  input      [2:0]    port_state_in_11_2_4,
  input      [2:0]    port_state_in_11_2_5,
  input      [2:0]    port_state_in_11_2_6,
  input      [2:0]    port_state_in_11_2_7,
  input      [2:0]    port_state_in_11_3_0,
  input      [2:0]    port_state_in_11_3_1,
  input      [2:0]    port_state_in_11_3_2,
  input      [2:0]    port_state_in_11_3_3,
  input      [2:0]    port_state_in_11_3_4,
  input      [2:0]    port_state_in_11_3_5,
  input      [2:0]    port_state_in_11_3_6,
  input      [2:0]    port_state_in_11_3_7,
  input      [2:0]    port_state_in_12_0_0,
  input      [2:0]    port_state_in_12_0_1,
  input      [2:0]    port_state_in_12_0_2,
  input      [2:0]    port_state_in_12_0_3,
  input      [2:0]    port_state_in_12_0_4,
  input      [2:0]    port_state_in_12_0_5,
  input      [2:0]    port_state_in_12_0_6,
  input      [2:0]    port_state_in_12_0_7,
  input      [2:0]    port_state_in_12_1_0,
  input      [2:0]    port_state_in_12_1_1,
  input      [2:0]    port_state_in_12_1_2,
  input      [2:0]    port_state_in_12_1_3,
  input      [2:0]    port_state_in_12_1_4,
  input      [2:0]    port_state_in_12_1_5,
  input      [2:0]    port_state_in_12_1_6,
  input      [2:0]    port_state_in_12_1_7,
  input      [2:0]    port_state_in_12_2_0,
  input      [2:0]    port_state_in_12_2_1,
  input      [2:0]    port_state_in_12_2_2,
  input      [2:0]    port_state_in_12_2_3,
  input      [2:0]    port_state_in_12_2_4,
  input      [2:0]    port_state_in_12_2_5,
  input      [2:0]    port_state_in_12_2_6,
  input      [2:0]    port_state_in_12_2_7,
  input      [2:0]    port_state_in_12_3_0,
  input      [2:0]    port_state_in_12_3_1,
  input      [2:0]    port_state_in_12_3_2,
  input      [2:0]    port_state_in_12_3_3,
  input      [2:0]    port_state_in_12_3_4,
  input      [2:0]    port_state_in_12_3_5,
  input      [2:0]    port_state_in_12_3_6,
  input      [2:0]    port_state_in_12_3_7,
  input      [2:0]    port_state_in_13_0_0,
  input      [2:0]    port_state_in_13_0_1,
  input      [2:0]    port_state_in_13_0_2,
  input      [2:0]    port_state_in_13_0_3,
  input      [2:0]    port_state_in_13_0_4,
  input      [2:0]    port_state_in_13_0_5,
  input      [2:0]    port_state_in_13_0_6,
  input      [2:0]    port_state_in_13_0_7,
  input      [2:0]    port_state_in_13_1_0,
  input      [2:0]    port_state_in_13_1_1,
  input      [2:0]    port_state_in_13_1_2,
  input      [2:0]    port_state_in_13_1_3,
  input      [2:0]    port_state_in_13_1_4,
  input      [2:0]    port_state_in_13_1_5,
  input      [2:0]    port_state_in_13_1_6,
  input      [2:0]    port_state_in_13_1_7,
  input      [2:0]    port_state_in_13_2_0,
  input      [2:0]    port_state_in_13_2_1,
  input      [2:0]    port_state_in_13_2_2,
  input      [2:0]    port_state_in_13_2_3,
  input      [2:0]    port_state_in_13_2_4,
  input      [2:0]    port_state_in_13_2_5,
  input      [2:0]    port_state_in_13_2_6,
  input      [2:0]    port_state_in_13_2_7,
  input      [2:0]    port_state_in_13_3_0,
  input      [2:0]    port_state_in_13_3_1,
  input      [2:0]    port_state_in_13_3_2,
  input      [2:0]    port_state_in_13_3_3,
  input      [2:0]    port_state_in_13_3_4,
  input      [2:0]    port_state_in_13_3_5,
  input      [2:0]    port_state_in_13_3_6,
  input      [2:0]    port_state_in_13_3_7,
  input      [2:0]    port_state_in_14_0_0,
  input      [2:0]    port_state_in_14_0_1,
  input      [2:0]    port_state_in_14_0_2,
  input      [2:0]    port_state_in_14_0_3,
  input      [2:0]    port_state_in_14_0_4,
  input      [2:0]    port_state_in_14_0_5,
  input      [2:0]    port_state_in_14_0_6,
  input      [2:0]    port_state_in_14_0_7,
  input      [2:0]    port_state_in_14_1_0,
  input      [2:0]    port_state_in_14_1_1,
  input      [2:0]    port_state_in_14_1_2,
  input      [2:0]    port_state_in_14_1_3,
  input      [2:0]    port_state_in_14_1_4,
  input      [2:0]    port_state_in_14_1_5,
  input      [2:0]    port_state_in_14_1_6,
  input      [2:0]    port_state_in_14_1_7,
  input      [2:0]    port_state_in_14_2_0,
  input      [2:0]    port_state_in_14_2_1,
  input      [2:0]    port_state_in_14_2_2,
  input      [2:0]    port_state_in_14_2_3,
  input      [2:0]    port_state_in_14_2_4,
  input      [2:0]    port_state_in_14_2_5,
  input      [2:0]    port_state_in_14_2_6,
  input      [2:0]    port_state_in_14_2_7,
  input      [2:0]    port_state_in_14_3_0,
  input      [2:0]    port_state_in_14_3_1,
  input      [2:0]    port_state_in_14_3_2,
  input      [2:0]    port_state_in_14_3_3,
  input      [2:0]    port_state_in_14_3_4,
  input      [2:0]    port_state_in_14_3_5,
  input      [2:0]    port_state_in_14_3_6,
  input      [2:0]    port_state_in_14_3_7,
  input      [2:0]    port_state_in_15_0_0,
  input      [2:0]    port_state_in_15_0_1,
  input      [2:0]    port_state_in_15_0_2,
  input      [2:0]    port_state_in_15_0_3,
  input      [2:0]    port_state_in_15_0_4,
  input      [2:0]    port_state_in_15_0_5,
  input      [2:0]    port_state_in_15_0_6,
  input      [2:0]    port_state_in_15_0_7,
  input      [2:0]    port_state_in_15_1_0,
  input      [2:0]    port_state_in_15_1_1,
  input      [2:0]    port_state_in_15_1_2,
  input      [2:0]    port_state_in_15_1_3,
  input      [2:0]    port_state_in_15_1_4,
  input      [2:0]    port_state_in_15_1_5,
  input      [2:0]    port_state_in_15_1_6,
  input      [2:0]    port_state_in_15_1_7,
  input      [2:0]    port_state_in_15_2_0,
  input      [2:0]    port_state_in_15_2_1,
  input      [2:0]    port_state_in_15_2_2,
  input      [2:0]    port_state_in_15_2_3,
  input      [2:0]    port_state_in_15_2_4,
  input      [2:0]    port_state_in_15_2_5,
  input      [2:0]    port_state_in_15_2_6,
  input      [2:0]    port_state_in_15_2_7,
  input      [2:0]    port_state_in_15_3_0,
  input      [2:0]    port_state_in_15_3_1,
  input      [2:0]    port_state_in_15_3_2,
  input      [2:0]    port_state_in_15_3_3,
  input      [2:0]    port_state_in_15_3_4,
  input      [2:0]    port_state_in_15_3_5,
  input      [2:0]    port_state_in_15_3_6,
  input      [2:0]    port_state_in_15_3_7,
  input      [2:0]    port_key_0_0_0,
  input      [2:0]    port_key_0_0_1,
  input      [2:0]    port_key_0_0_2,
  input      [2:0]    port_key_0_0_3,
  input      [2:0]    port_key_0_0_4,
  input      [2:0]    port_key_0_0_5,
  input      [2:0]    port_key_0_0_6,
  input      [2:0]    port_key_0_0_7,
  input      [2:0]    port_key_0_1_0,
  input      [2:0]    port_key_0_1_1,
  input      [2:0]    port_key_0_1_2,
  input      [2:0]    port_key_0_1_3,
  input      [2:0]    port_key_0_1_4,
  input      [2:0]    port_key_0_1_5,
  input      [2:0]    port_key_0_1_6,
  input      [2:0]    port_key_0_1_7,
  input      [2:0]    port_key_0_2_0,
  input      [2:0]    port_key_0_2_1,
  input      [2:0]    port_key_0_2_2,
  input      [2:0]    port_key_0_2_3,
  input      [2:0]    port_key_0_2_4,
  input      [2:0]    port_key_0_2_5,
  input      [2:0]    port_key_0_2_6,
  input      [2:0]    port_key_0_2_7,
  input      [2:0]    port_key_0_3_0,
  input      [2:0]    port_key_0_3_1,
  input      [2:0]    port_key_0_3_2,
  input      [2:0]    port_key_0_3_3,
  input      [2:0]    port_key_0_3_4,
  input      [2:0]    port_key_0_3_5,
  input      [2:0]    port_key_0_3_6,
  input      [2:0]    port_key_0_3_7,
  input      [2:0]    port_key_1_0_0,
  input      [2:0]    port_key_1_0_1,
  input      [2:0]    port_key_1_0_2,
  input      [2:0]    port_key_1_0_3,
  input      [2:0]    port_key_1_0_4,
  input      [2:0]    port_key_1_0_5,
  input      [2:0]    port_key_1_0_6,
  input      [2:0]    port_key_1_0_7,
  input      [2:0]    port_key_1_1_0,
  input      [2:0]    port_key_1_1_1,
  input      [2:0]    port_key_1_1_2,
  input      [2:0]    port_key_1_1_3,
  input      [2:0]    port_key_1_1_4,
  input      [2:0]    port_key_1_1_5,
  input      [2:0]    port_key_1_1_6,
  input      [2:0]    port_key_1_1_7,
  input      [2:0]    port_key_1_2_0,
  input      [2:0]    port_key_1_2_1,
  input      [2:0]    port_key_1_2_2,
  input      [2:0]    port_key_1_2_3,
  input      [2:0]    port_key_1_2_4,
  input      [2:0]    port_key_1_2_5,
  input      [2:0]    port_key_1_2_6,
  input      [2:0]    port_key_1_2_7,
  input      [2:0]    port_key_1_3_0,
  input      [2:0]    port_key_1_3_1,
  input      [2:0]    port_key_1_3_2,
  input      [2:0]    port_key_1_3_3,
  input      [2:0]    port_key_1_3_4,
  input      [2:0]    port_key_1_3_5,
  input      [2:0]    port_key_1_3_6,
  input      [2:0]    port_key_1_3_7,
  input      [2:0]    port_key_2_0_0,
  input      [2:0]    port_key_2_0_1,
  input      [2:0]    port_key_2_0_2,
  input      [2:0]    port_key_2_0_3,
  input      [2:0]    port_key_2_0_4,
  input      [2:0]    port_key_2_0_5,
  input      [2:0]    port_key_2_0_6,
  input      [2:0]    port_key_2_0_7,
  input      [2:0]    port_key_2_1_0,
  input      [2:0]    port_key_2_1_1,
  input      [2:0]    port_key_2_1_2,
  input      [2:0]    port_key_2_1_3,
  input      [2:0]    port_key_2_1_4,
  input      [2:0]    port_key_2_1_5,
  input      [2:0]    port_key_2_1_6,
  input      [2:0]    port_key_2_1_7,
  input      [2:0]    port_key_2_2_0,
  input      [2:0]    port_key_2_2_1,
  input      [2:0]    port_key_2_2_2,
  input      [2:0]    port_key_2_2_3,
  input      [2:0]    port_key_2_2_4,
  input      [2:0]    port_key_2_2_5,
  input      [2:0]    port_key_2_2_6,
  input      [2:0]    port_key_2_2_7,
  input      [2:0]    port_key_2_3_0,
  input      [2:0]    port_key_2_3_1,
  input      [2:0]    port_key_2_3_2,
  input      [2:0]    port_key_2_3_3,
  input      [2:0]    port_key_2_3_4,
  input      [2:0]    port_key_2_3_5,
  input      [2:0]    port_key_2_3_6,
  input      [2:0]    port_key_2_3_7,
  input      [2:0]    port_key_3_0_0,
  input      [2:0]    port_key_3_0_1,
  input      [2:0]    port_key_3_0_2,
  input      [2:0]    port_key_3_0_3,
  input      [2:0]    port_key_3_0_4,
  input      [2:0]    port_key_3_0_5,
  input      [2:0]    port_key_3_0_6,
  input      [2:0]    port_key_3_0_7,
  input      [2:0]    port_key_3_1_0,
  input      [2:0]    port_key_3_1_1,
  input      [2:0]    port_key_3_1_2,
  input      [2:0]    port_key_3_1_3,
  input      [2:0]    port_key_3_1_4,
  input      [2:0]    port_key_3_1_5,
  input      [2:0]    port_key_3_1_6,
  input      [2:0]    port_key_3_1_7,
  input      [2:0]    port_key_3_2_0,
  input      [2:0]    port_key_3_2_1,
  input      [2:0]    port_key_3_2_2,
  input      [2:0]    port_key_3_2_3,
  input      [2:0]    port_key_3_2_4,
  input      [2:0]    port_key_3_2_5,
  input      [2:0]    port_key_3_2_6,
  input      [2:0]    port_key_3_2_7,
  input      [2:0]    port_key_3_3_0,
  input      [2:0]    port_key_3_3_1,
  input      [2:0]    port_key_3_3_2,
  input      [2:0]    port_key_3_3_3,
  input      [2:0]    port_key_3_3_4,
  input      [2:0]    port_key_3_3_5,
  input      [2:0]    port_key_3_3_6,
  input      [2:0]    port_key_3_3_7,
  input      [2:0]    port_key_4_0_0,
  input      [2:0]    port_key_4_0_1,
  input      [2:0]    port_key_4_0_2,
  input      [2:0]    port_key_4_0_3,
  input      [2:0]    port_key_4_0_4,
  input      [2:0]    port_key_4_0_5,
  input      [2:0]    port_key_4_0_6,
  input      [2:0]    port_key_4_0_7,
  input      [2:0]    port_key_4_1_0,
  input      [2:0]    port_key_4_1_1,
  input      [2:0]    port_key_4_1_2,
  input      [2:0]    port_key_4_1_3,
  input      [2:0]    port_key_4_1_4,
  input      [2:0]    port_key_4_1_5,
  input      [2:0]    port_key_4_1_6,
  input      [2:0]    port_key_4_1_7,
  input      [2:0]    port_key_4_2_0,
  input      [2:0]    port_key_4_2_1,
  input      [2:0]    port_key_4_2_2,
  input      [2:0]    port_key_4_2_3,
  input      [2:0]    port_key_4_2_4,
  input      [2:0]    port_key_4_2_5,
  input      [2:0]    port_key_4_2_6,
  input      [2:0]    port_key_4_2_7,
  input      [2:0]    port_key_4_3_0,
  input      [2:0]    port_key_4_3_1,
  input      [2:0]    port_key_4_3_2,
  input      [2:0]    port_key_4_3_3,
  input      [2:0]    port_key_4_3_4,
  input      [2:0]    port_key_4_3_5,
  input      [2:0]    port_key_4_3_6,
  input      [2:0]    port_key_4_3_7,
  input      [2:0]    port_key_5_0_0,
  input      [2:0]    port_key_5_0_1,
  input      [2:0]    port_key_5_0_2,
  input      [2:0]    port_key_5_0_3,
  input      [2:0]    port_key_5_0_4,
  input      [2:0]    port_key_5_0_5,
  input      [2:0]    port_key_5_0_6,
  input      [2:0]    port_key_5_0_7,
  input      [2:0]    port_key_5_1_0,
  input      [2:0]    port_key_5_1_1,
  input      [2:0]    port_key_5_1_2,
  input      [2:0]    port_key_5_1_3,
  input      [2:0]    port_key_5_1_4,
  input      [2:0]    port_key_5_1_5,
  input      [2:0]    port_key_5_1_6,
  input      [2:0]    port_key_5_1_7,
  input      [2:0]    port_key_5_2_0,
  input      [2:0]    port_key_5_2_1,
  input      [2:0]    port_key_5_2_2,
  input      [2:0]    port_key_5_2_3,
  input      [2:0]    port_key_5_2_4,
  input      [2:0]    port_key_5_2_5,
  input      [2:0]    port_key_5_2_6,
  input      [2:0]    port_key_5_2_7,
  input      [2:0]    port_key_5_3_0,
  input      [2:0]    port_key_5_3_1,
  input      [2:0]    port_key_5_3_2,
  input      [2:0]    port_key_5_3_3,
  input      [2:0]    port_key_5_3_4,
  input      [2:0]    port_key_5_3_5,
  input      [2:0]    port_key_5_3_6,
  input      [2:0]    port_key_5_3_7,
  input      [2:0]    port_key_6_0_0,
  input      [2:0]    port_key_6_0_1,
  input      [2:0]    port_key_6_0_2,
  input      [2:0]    port_key_6_0_3,
  input      [2:0]    port_key_6_0_4,
  input      [2:0]    port_key_6_0_5,
  input      [2:0]    port_key_6_0_6,
  input      [2:0]    port_key_6_0_7,
  input      [2:0]    port_key_6_1_0,
  input      [2:0]    port_key_6_1_1,
  input      [2:0]    port_key_6_1_2,
  input      [2:0]    port_key_6_1_3,
  input      [2:0]    port_key_6_1_4,
  input      [2:0]    port_key_6_1_5,
  input      [2:0]    port_key_6_1_6,
  input      [2:0]    port_key_6_1_7,
  input      [2:0]    port_key_6_2_0,
  input      [2:0]    port_key_6_2_1,
  input      [2:0]    port_key_6_2_2,
  input      [2:0]    port_key_6_2_3,
  input      [2:0]    port_key_6_2_4,
  input      [2:0]    port_key_6_2_5,
  input      [2:0]    port_key_6_2_6,
  input      [2:0]    port_key_6_2_7,
  input      [2:0]    port_key_6_3_0,
  input      [2:0]    port_key_6_3_1,
  input      [2:0]    port_key_6_3_2,
  input      [2:0]    port_key_6_3_3,
  input      [2:0]    port_key_6_3_4,
  input      [2:0]    port_key_6_3_5,
  input      [2:0]    port_key_6_3_6,
  input      [2:0]    port_key_6_3_7,
  input      [2:0]    port_key_7_0_0,
  input      [2:0]    port_key_7_0_1,
  input      [2:0]    port_key_7_0_2,
  input      [2:0]    port_key_7_0_3,
  input      [2:0]    port_key_7_0_4,
  input      [2:0]    port_key_7_0_5,
  input      [2:0]    port_key_7_0_6,
  input      [2:0]    port_key_7_0_7,
  input      [2:0]    port_key_7_1_0,
  input      [2:0]    port_key_7_1_1,
  input      [2:0]    port_key_7_1_2,
  input      [2:0]    port_key_7_1_3,
  input      [2:0]    port_key_7_1_4,
  input      [2:0]    port_key_7_1_5,
  input      [2:0]    port_key_7_1_6,
  input      [2:0]    port_key_7_1_7,
  input      [2:0]    port_key_7_2_0,
  input      [2:0]    port_key_7_2_1,
  input      [2:0]    port_key_7_2_2,
  input      [2:0]    port_key_7_2_3,
  input      [2:0]    port_key_7_2_4,
  input      [2:0]    port_key_7_2_5,
  input      [2:0]    port_key_7_2_6,
  input      [2:0]    port_key_7_2_7,
  input      [2:0]    port_key_7_3_0,
  input      [2:0]    port_key_7_3_1,
  input      [2:0]    port_key_7_3_2,
  input      [2:0]    port_key_7_3_3,
  input      [2:0]    port_key_7_3_4,
  input      [2:0]    port_key_7_3_5,
  input      [2:0]    port_key_7_3_6,
  input      [2:0]    port_key_7_3_7,
  input      [2:0]    port_key_8_0_0,
  input      [2:0]    port_key_8_0_1,
  input      [2:0]    port_key_8_0_2,
  input      [2:0]    port_key_8_0_3,
  input      [2:0]    port_key_8_0_4,
  input      [2:0]    port_key_8_0_5,
  input      [2:0]    port_key_8_0_6,
  input      [2:0]    port_key_8_0_7,
  input      [2:0]    port_key_8_1_0,
  input      [2:0]    port_key_8_1_1,
  input      [2:0]    port_key_8_1_2,
  input      [2:0]    port_key_8_1_3,
  input      [2:0]    port_key_8_1_4,
  input      [2:0]    port_key_8_1_5,
  input      [2:0]    port_key_8_1_6,
  input      [2:0]    port_key_8_1_7,
  input      [2:0]    port_key_8_2_0,
  input      [2:0]    port_key_8_2_1,
  input      [2:0]    port_key_8_2_2,
  input      [2:0]    port_key_8_2_3,
  input      [2:0]    port_key_8_2_4,
  input      [2:0]    port_key_8_2_5,
  input      [2:0]    port_key_8_2_6,
  input      [2:0]    port_key_8_2_7,
  input      [2:0]    port_key_8_3_0,
  input      [2:0]    port_key_8_3_1,
  input      [2:0]    port_key_8_3_2,
  input      [2:0]    port_key_8_3_3,
  input      [2:0]    port_key_8_3_4,
  input      [2:0]    port_key_8_3_5,
  input      [2:0]    port_key_8_3_6,
  input      [2:0]    port_key_8_3_7,
  input      [2:0]    port_key_9_0_0,
  input      [2:0]    port_key_9_0_1,
  input      [2:0]    port_key_9_0_2,
  input      [2:0]    port_key_9_0_3,
  input      [2:0]    port_key_9_0_4,
  input      [2:0]    port_key_9_0_5,
  input      [2:0]    port_key_9_0_6,
  input      [2:0]    port_key_9_0_7,
  input      [2:0]    port_key_9_1_0,
  input      [2:0]    port_key_9_1_1,
  input      [2:0]    port_key_9_1_2,
  input      [2:0]    port_key_9_1_3,
  input      [2:0]    port_key_9_1_4,
  input      [2:0]    port_key_9_1_5,
  input      [2:0]    port_key_9_1_6,
  input      [2:0]    port_key_9_1_7,
  input      [2:0]    port_key_9_2_0,
  input      [2:0]    port_key_9_2_1,
  input      [2:0]    port_key_9_2_2,
  input      [2:0]    port_key_9_2_3,
  input      [2:0]    port_key_9_2_4,
  input      [2:0]    port_key_9_2_5,
  input      [2:0]    port_key_9_2_6,
  input      [2:0]    port_key_9_2_7,
  input      [2:0]    port_key_9_3_0,
  input      [2:0]    port_key_9_3_1,
  input      [2:0]    port_key_9_3_2,
  input      [2:0]    port_key_9_3_3,
  input      [2:0]    port_key_9_3_4,
  input      [2:0]    port_key_9_3_5,
  input      [2:0]    port_key_9_3_6,
  input      [2:0]    port_key_9_3_7,
  input      [2:0]    port_key_10_0_0,
  input      [2:0]    port_key_10_0_1,
  input      [2:0]    port_key_10_0_2,
  input      [2:0]    port_key_10_0_3,
  input      [2:0]    port_key_10_0_4,
  input      [2:0]    port_key_10_0_5,
  input      [2:0]    port_key_10_0_6,
  input      [2:0]    port_key_10_0_7,
  input      [2:0]    port_key_10_1_0,
  input      [2:0]    port_key_10_1_1,
  input      [2:0]    port_key_10_1_2,
  input      [2:0]    port_key_10_1_3,
  input      [2:0]    port_key_10_1_4,
  input      [2:0]    port_key_10_1_5,
  input      [2:0]    port_key_10_1_6,
  input      [2:0]    port_key_10_1_7,
  input      [2:0]    port_key_10_2_0,
  input      [2:0]    port_key_10_2_1,
  input      [2:0]    port_key_10_2_2,
  input      [2:0]    port_key_10_2_3,
  input      [2:0]    port_key_10_2_4,
  input      [2:0]    port_key_10_2_5,
  input      [2:0]    port_key_10_2_6,
  input      [2:0]    port_key_10_2_7,
  input      [2:0]    port_key_10_3_0,
  input      [2:0]    port_key_10_3_1,
  input      [2:0]    port_key_10_3_2,
  input      [2:0]    port_key_10_3_3,
  input      [2:0]    port_key_10_3_4,
  input      [2:0]    port_key_10_3_5,
  input      [2:0]    port_key_10_3_6,
  input      [2:0]    port_key_10_3_7,
  input      [2:0]    port_key_11_0_0,
  input      [2:0]    port_key_11_0_1,
  input      [2:0]    port_key_11_0_2,
  input      [2:0]    port_key_11_0_3,
  input      [2:0]    port_key_11_0_4,
  input      [2:0]    port_key_11_0_5,
  input      [2:0]    port_key_11_0_6,
  input      [2:0]    port_key_11_0_7,
  input      [2:0]    port_key_11_1_0,
  input      [2:0]    port_key_11_1_1,
  input      [2:0]    port_key_11_1_2,
  input      [2:0]    port_key_11_1_3,
  input      [2:0]    port_key_11_1_4,
  input      [2:0]    port_key_11_1_5,
  input      [2:0]    port_key_11_1_6,
  input      [2:0]    port_key_11_1_7,
  input      [2:0]    port_key_11_2_0,
  input      [2:0]    port_key_11_2_1,
  input      [2:0]    port_key_11_2_2,
  input      [2:0]    port_key_11_2_3,
  input      [2:0]    port_key_11_2_4,
  input      [2:0]    port_key_11_2_5,
  input      [2:0]    port_key_11_2_6,
  input      [2:0]    port_key_11_2_7,
  input      [2:0]    port_key_11_3_0,
  input      [2:0]    port_key_11_3_1,
  input      [2:0]    port_key_11_3_2,
  input      [2:0]    port_key_11_3_3,
  input      [2:0]    port_key_11_3_4,
  input      [2:0]    port_key_11_3_5,
  input      [2:0]    port_key_11_3_6,
  input      [2:0]    port_key_11_3_7,
  input      [2:0]    port_key_12_0_0,
  input      [2:0]    port_key_12_0_1,
  input      [2:0]    port_key_12_0_2,
  input      [2:0]    port_key_12_0_3,
  input      [2:0]    port_key_12_0_4,
  input      [2:0]    port_key_12_0_5,
  input      [2:0]    port_key_12_0_6,
  input      [2:0]    port_key_12_0_7,
  input      [2:0]    port_key_12_1_0,
  input      [2:0]    port_key_12_1_1,
  input      [2:0]    port_key_12_1_2,
  input      [2:0]    port_key_12_1_3,
  input      [2:0]    port_key_12_1_4,
  input      [2:0]    port_key_12_1_5,
  input      [2:0]    port_key_12_1_6,
  input      [2:0]    port_key_12_1_7,
  input      [2:0]    port_key_12_2_0,
  input      [2:0]    port_key_12_2_1,
  input      [2:0]    port_key_12_2_2,
  input      [2:0]    port_key_12_2_3,
  input      [2:0]    port_key_12_2_4,
  input      [2:0]    port_key_12_2_5,
  input      [2:0]    port_key_12_2_6,
  input      [2:0]    port_key_12_2_7,
  input      [2:0]    port_key_12_3_0,
  input      [2:0]    port_key_12_3_1,
  input      [2:0]    port_key_12_3_2,
  input      [2:0]    port_key_12_3_3,
  input      [2:0]    port_key_12_3_4,
  input      [2:0]    port_key_12_3_5,
  input      [2:0]    port_key_12_3_6,
  input      [2:0]    port_key_12_3_7,
  input      [2:0]    port_key_13_0_0,
  input      [2:0]    port_key_13_0_1,
  input      [2:0]    port_key_13_0_2,
  input      [2:0]    port_key_13_0_3,
  input      [2:0]    port_key_13_0_4,
  input      [2:0]    port_key_13_0_5,
  input      [2:0]    port_key_13_0_6,
  input      [2:0]    port_key_13_0_7,
  input      [2:0]    port_key_13_1_0,
  input      [2:0]    port_key_13_1_1,
  input      [2:0]    port_key_13_1_2,
  input      [2:0]    port_key_13_1_3,
  input      [2:0]    port_key_13_1_4,
  input      [2:0]    port_key_13_1_5,
  input      [2:0]    port_key_13_1_6,
  input      [2:0]    port_key_13_1_7,
  input      [2:0]    port_key_13_2_0,
  input      [2:0]    port_key_13_2_1,
  input      [2:0]    port_key_13_2_2,
  input      [2:0]    port_key_13_2_3,
  input      [2:0]    port_key_13_2_4,
  input      [2:0]    port_key_13_2_5,
  input      [2:0]    port_key_13_2_6,
  input      [2:0]    port_key_13_2_7,
  input      [2:0]    port_key_13_3_0,
  input      [2:0]    port_key_13_3_1,
  input      [2:0]    port_key_13_3_2,
  input      [2:0]    port_key_13_3_3,
  input      [2:0]    port_key_13_3_4,
  input      [2:0]    port_key_13_3_5,
  input      [2:0]    port_key_13_3_6,
  input      [2:0]    port_key_13_3_7,
  input      [2:0]    port_key_14_0_0,
  input      [2:0]    port_key_14_0_1,
  input      [2:0]    port_key_14_0_2,
  input      [2:0]    port_key_14_0_3,
  input      [2:0]    port_key_14_0_4,
  input      [2:0]    port_key_14_0_5,
  input      [2:0]    port_key_14_0_6,
  input      [2:0]    port_key_14_0_7,
  input      [2:0]    port_key_14_1_0,
  input      [2:0]    port_key_14_1_1,
  input      [2:0]    port_key_14_1_2,
  input      [2:0]    port_key_14_1_3,
  input      [2:0]    port_key_14_1_4,
  input      [2:0]    port_key_14_1_5,
  input      [2:0]    port_key_14_1_6,
  input      [2:0]    port_key_14_1_7,
  input      [2:0]    port_key_14_2_0,
  input      [2:0]    port_key_14_2_1,
  input      [2:0]    port_key_14_2_2,
  input      [2:0]    port_key_14_2_3,
  input      [2:0]    port_key_14_2_4,
  input      [2:0]    port_key_14_2_5,
  input      [2:0]    port_key_14_2_6,
  input      [2:0]    port_key_14_2_7,
  input      [2:0]    port_key_14_3_0,
  input      [2:0]    port_key_14_3_1,
  input      [2:0]    port_key_14_3_2,
  input      [2:0]    port_key_14_3_3,
  input      [2:0]    port_key_14_3_4,
  input      [2:0]    port_key_14_3_5,
  input      [2:0]    port_key_14_3_6,
  input      [2:0]    port_key_14_3_7,
  input      [2:0]    port_key_15_0_0,
  input      [2:0]    port_key_15_0_1,
  input      [2:0]    port_key_15_0_2,
  input      [2:0]    port_key_15_0_3,
  input      [2:0]    port_key_15_0_4,
  input      [2:0]    port_key_15_0_5,
  input      [2:0]    port_key_15_0_6,
  input      [2:0]    port_key_15_0_7,
  input      [2:0]    port_key_15_1_0,
  input      [2:0]    port_key_15_1_1,
  input      [2:0]    port_key_15_1_2,
  input      [2:0]    port_key_15_1_3,
  input      [2:0]    port_key_15_1_4,
  input      [2:0]    port_key_15_1_5,
  input      [2:0]    port_key_15_1_6,
  input      [2:0]    port_key_15_1_7,
  input      [2:0]    port_key_15_2_0,
  input      [2:0]    port_key_15_2_1,
  input      [2:0]    port_key_15_2_2,
  input      [2:0]    port_key_15_2_3,
  input      [2:0]    port_key_15_2_4,
  input      [2:0]    port_key_15_2_5,
  input      [2:0]    port_key_15_2_6,
  input      [2:0]    port_key_15_2_7,
  input      [2:0]    port_key_15_3_0,
  input      [2:0]    port_key_15_3_1,
  input      [2:0]    port_key_15_3_2,
  input      [2:0]    port_key_15_3_3,
  input      [2:0]    port_key_15_3_4,
  input      [2:0]    port_key_15_3_5,
  input      [2:0]    port_key_15_3_6,
  input      [2:0]    port_key_15_3_7,
  output     [2:0]    port_state_out_0_0_0,
  output     [2:0]    port_state_out_0_0_1,
  output     [2:0]    port_state_out_0_0_2,
  output     [2:0]    port_state_out_0_0_3,
  output     [2:0]    port_state_out_0_0_4,
  output     [2:0]    port_state_out_0_0_5,
  output     [2:0]    port_state_out_0_0_6,
  output     [2:0]    port_state_out_0_0_7,
  output     [2:0]    port_state_out_0_1_0,
  output     [2:0]    port_state_out_0_1_1,
  output     [2:0]    port_state_out_0_1_2,
  output     [2:0]    port_state_out_0_1_3,
  output     [2:0]    port_state_out_0_1_4,
  output     [2:0]    port_state_out_0_1_5,
  output     [2:0]    port_state_out_0_1_6,
  output     [2:0]    port_state_out_0_1_7,
  output     [2:0]    port_state_out_0_2_0,
  output     [2:0]    port_state_out_0_2_1,
  output     [2:0]    port_state_out_0_2_2,
  output     [2:0]    port_state_out_0_2_3,
  output     [2:0]    port_state_out_0_2_4,
  output     [2:0]    port_state_out_0_2_5,
  output     [2:0]    port_state_out_0_2_6,
  output     [2:0]    port_state_out_0_2_7,
  output     [2:0]    port_state_out_0_3_0,
  output     [2:0]    port_state_out_0_3_1,
  output     [2:0]    port_state_out_0_3_2,
  output     [2:0]    port_state_out_0_3_3,
  output     [2:0]    port_state_out_0_3_4,
  output     [2:0]    port_state_out_0_3_5,
  output     [2:0]    port_state_out_0_3_6,
  output     [2:0]    port_state_out_0_3_7,
  output     [2:0]    port_state_out_1_0_0,
  output     [2:0]    port_state_out_1_0_1,
  output     [2:0]    port_state_out_1_0_2,
  output     [2:0]    port_state_out_1_0_3,
  output     [2:0]    port_state_out_1_0_4,
  output     [2:0]    port_state_out_1_0_5,
  output     [2:0]    port_state_out_1_0_6,
  output     [2:0]    port_state_out_1_0_7,
  output     [2:0]    port_state_out_1_1_0,
  output     [2:0]    port_state_out_1_1_1,
  output     [2:0]    port_state_out_1_1_2,
  output     [2:0]    port_state_out_1_1_3,
  output     [2:0]    port_state_out_1_1_4,
  output     [2:0]    port_state_out_1_1_5,
  output     [2:0]    port_state_out_1_1_6,
  output     [2:0]    port_state_out_1_1_7,
  output     [2:0]    port_state_out_1_2_0,
  output     [2:0]    port_state_out_1_2_1,
  output     [2:0]    port_state_out_1_2_2,
  output     [2:0]    port_state_out_1_2_3,
  output     [2:0]    port_state_out_1_2_4,
  output     [2:0]    port_state_out_1_2_5,
  output     [2:0]    port_state_out_1_2_6,
  output     [2:0]    port_state_out_1_2_7,
  output     [2:0]    port_state_out_1_3_0,
  output     [2:0]    port_state_out_1_3_1,
  output     [2:0]    port_state_out_1_3_2,
  output     [2:0]    port_state_out_1_3_3,
  output     [2:0]    port_state_out_1_3_4,
  output     [2:0]    port_state_out_1_3_5,
  output     [2:0]    port_state_out_1_3_6,
  output     [2:0]    port_state_out_1_3_7,
  output     [2:0]    port_state_out_2_0_0,
  output     [2:0]    port_state_out_2_0_1,
  output     [2:0]    port_state_out_2_0_2,
  output     [2:0]    port_state_out_2_0_3,
  output     [2:0]    port_state_out_2_0_4,
  output     [2:0]    port_state_out_2_0_5,
  output     [2:0]    port_state_out_2_0_6,
  output     [2:0]    port_state_out_2_0_7,
  output     [2:0]    port_state_out_2_1_0,
  output     [2:0]    port_state_out_2_1_1,
  output     [2:0]    port_state_out_2_1_2,
  output     [2:0]    port_state_out_2_1_3,
  output     [2:0]    port_state_out_2_1_4,
  output     [2:0]    port_state_out_2_1_5,
  output     [2:0]    port_state_out_2_1_6,
  output     [2:0]    port_state_out_2_1_7,
  output     [2:0]    port_state_out_2_2_0,
  output     [2:0]    port_state_out_2_2_1,
  output     [2:0]    port_state_out_2_2_2,
  output     [2:0]    port_state_out_2_2_3,
  output     [2:0]    port_state_out_2_2_4,
  output     [2:0]    port_state_out_2_2_5,
  output     [2:0]    port_state_out_2_2_6,
  output     [2:0]    port_state_out_2_2_7,
  output     [2:0]    port_state_out_2_3_0,
  output     [2:0]    port_state_out_2_3_1,
  output     [2:0]    port_state_out_2_3_2,
  output     [2:0]    port_state_out_2_3_3,
  output     [2:0]    port_state_out_2_3_4,
  output     [2:0]    port_state_out_2_3_5,
  output     [2:0]    port_state_out_2_3_6,
  output     [2:0]    port_state_out_2_3_7,
  output     [2:0]    port_state_out_3_0_0,
  output     [2:0]    port_state_out_3_0_1,
  output     [2:0]    port_state_out_3_0_2,
  output     [2:0]    port_state_out_3_0_3,
  output     [2:0]    port_state_out_3_0_4,
  output     [2:0]    port_state_out_3_0_5,
  output     [2:0]    port_state_out_3_0_6,
  output     [2:0]    port_state_out_3_0_7,
  output     [2:0]    port_state_out_3_1_0,
  output     [2:0]    port_state_out_3_1_1,
  output     [2:0]    port_state_out_3_1_2,
  output     [2:0]    port_state_out_3_1_3,
  output     [2:0]    port_state_out_3_1_4,
  output     [2:0]    port_state_out_3_1_5,
  output     [2:0]    port_state_out_3_1_6,
  output     [2:0]    port_state_out_3_1_7,
  output     [2:0]    port_state_out_3_2_0,
  output     [2:0]    port_state_out_3_2_1,
  output     [2:0]    port_state_out_3_2_2,
  output     [2:0]    port_state_out_3_2_3,
  output     [2:0]    port_state_out_3_2_4,
  output     [2:0]    port_state_out_3_2_5,
  output     [2:0]    port_state_out_3_2_6,
  output     [2:0]    port_state_out_3_2_7,
  output     [2:0]    port_state_out_3_3_0,
  output     [2:0]    port_state_out_3_3_1,
  output     [2:0]    port_state_out_3_3_2,
  output     [2:0]    port_state_out_3_3_3,
  output     [2:0]    port_state_out_3_3_4,
  output     [2:0]    port_state_out_3_3_5,
  output     [2:0]    port_state_out_3_3_6,
  output     [2:0]    port_state_out_3_3_7,
  output     [2:0]    port_state_out_4_0_0,
  output     [2:0]    port_state_out_4_0_1,
  output     [2:0]    port_state_out_4_0_2,
  output     [2:0]    port_state_out_4_0_3,
  output     [2:0]    port_state_out_4_0_4,
  output     [2:0]    port_state_out_4_0_5,
  output     [2:0]    port_state_out_4_0_6,
  output     [2:0]    port_state_out_4_0_7,
  output     [2:0]    port_state_out_4_1_0,
  output     [2:0]    port_state_out_4_1_1,
  output     [2:0]    port_state_out_4_1_2,
  output     [2:0]    port_state_out_4_1_3,
  output     [2:0]    port_state_out_4_1_4,
  output     [2:0]    port_state_out_4_1_5,
  output     [2:0]    port_state_out_4_1_6,
  output     [2:0]    port_state_out_4_1_7,
  output     [2:0]    port_state_out_4_2_0,
  output     [2:0]    port_state_out_4_2_1,
  output     [2:0]    port_state_out_4_2_2,
  output     [2:0]    port_state_out_4_2_3,
  output     [2:0]    port_state_out_4_2_4,
  output     [2:0]    port_state_out_4_2_5,
  output     [2:0]    port_state_out_4_2_6,
  output     [2:0]    port_state_out_4_2_7,
  output     [2:0]    port_state_out_4_3_0,
  output     [2:0]    port_state_out_4_3_1,
  output     [2:0]    port_state_out_4_3_2,
  output     [2:0]    port_state_out_4_3_3,
  output     [2:0]    port_state_out_4_3_4,
  output     [2:0]    port_state_out_4_3_5,
  output     [2:0]    port_state_out_4_3_6,
  output     [2:0]    port_state_out_4_3_7,
  output     [2:0]    port_state_out_5_0_0,
  output     [2:0]    port_state_out_5_0_1,
  output     [2:0]    port_state_out_5_0_2,
  output     [2:0]    port_state_out_5_0_3,
  output     [2:0]    port_state_out_5_0_4,
  output     [2:0]    port_state_out_5_0_5,
  output     [2:0]    port_state_out_5_0_6,
  output     [2:0]    port_state_out_5_0_7,
  output     [2:0]    port_state_out_5_1_0,
  output     [2:0]    port_state_out_5_1_1,
  output     [2:0]    port_state_out_5_1_2,
  output     [2:0]    port_state_out_5_1_3,
  output     [2:0]    port_state_out_5_1_4,
  output     [2:0]    port_state_out_5_1_5,
  output     [2:0]    port_state_out_5_1_6,
  output     [2:0]    port_state_out_5_1_7,
  output     [2:0]    port_state_out_5_2_0,
  output     [2:0]    port_state_out_5_2_1,
  output     [2:0]    port_state_out_5_2_2,
  output     [2:0]    port_state_out_5_2_3,
  output     [2:0]    port_state_out_5_2_4,
  output     [2:0]    port_state_out_5_2_5,
  output     [2:0]    port_state_out_5_2_6,
  output     [2:0]    port_state_out_5_2_7,
  output     [2:0]    port_state_out_5_3_0,
  output     [2:0]    port_state_out_5_3_1,
  output     [2:0]    port_state_out_5_3_2,
  output     [2:0]    port_state_out_5_3_3,
  output     [2:0]    port_state_out_5_3_4,
  output     [2:0]    port_state_out_5_3_5,
  output     [2:0]    port_state_out_5_3_6,
  output     [2:0]    port_state_out_5_3_7,
  output     [2:0]    port_state_out_6_0_0,
  output     [2:0]    port_state_out_6_0_1,
  output     [2:0]    port_state_out_6_0_2,
  output     [2:0]    port_state_out_6_0_3,
  output     [2:0]    port_state_out_6_0_4,
  output     [2:0]    port_state_out_6_0_5,
  output     [2:0]    port_state_out_6_0_6,
  output     [2:0]    port_state_out_6_0_7,
  output     [2:0]    port_state_out_6_1_0,
  output     [2:0]    port_state_out_6_1_1,
  output     [2:0]    port_state_out_6_1_2,
  output     [2:0]    port_state_out_6_1_3,
  output     [2:0]    port_state_out_6_1_4,
  output     [2:0]    port_state_out_6_1_5,
  output     [2:0]    port_state_out_6_1_6,
  output     [2:0]    port_state_out_6_1_7,
  output     [2:0]    port_state_out_6_2_0,
  output     [2:0]    port_state_out_6_2_1,
  output     [2:0]    port_state_out_6_2_2,
  output     [2:0]    port_state_out_6_2_3,
  output     [2:0]    port_state_out_6_2_4,
  output     [2:0]    port_state_out_6_2_5,
  output     [2:0]    port_state_out_6_2_6,
  output     [2:0]    port_state_out_6_2_7,
  output     [2:0]    port_state_out_6_3_0,
  output     [2:0]    port_state_out_6_3_1,
  output     [2:0]    port_state_out_6_3_2,
  output     [2:0]    port_state_out_6_3_3,
  output     [2:0]    port_state_out_6_3_4,
  output     [2:0]    port_state_out_6_3_5,
  output     [2:0]    port_state_out_6_3_6,
  output     [2:0]    port_state_out_6_3_7,
  output     [2:0]    port_state_out_7_0_0,
  output     [2:0]    port_state_out_7_0_1,
  output     [2:0]    port_state_out_7_0_2,
  output     [2:0]    port_state_out_7_0_3,
  output     [2:0]    port_state_out_7_0_4,
  output     [2:0]    port_state_out_7_0_5,
  output     [2:0]    port_state_out_7_0_6,
  output     [2:0]    port_state_out_7_0_7,
  output     [2:0]    port_state_out_7_1_0,
  output     [2:0]    port_state_out_7_1_1,
  output     [2:0]    port_state_out_7_1_2,
  output     [2:0]    port_state_out_7_1_3,
  output     [2:0]    port_state_out_7_1_4,
  output     [2:0]    port_state_out_7_1_5,
  output     [2:0]    port_state_out_7_1_6,
  output     [2:0]    port_state_out_7_1_7,
  output     [2:0]    port_state_out_7_2_0,
  output     [2:0]    port_state_out_7_2_1,
  output     [2:0]    port_state_out_7_2_2,
  output     [2:0]    port_state_out_7_2_3,
  output     [2:0]    port_state_out_7_2_4,
  output     [2:0]    port_state_out_7_2_5,
  output     [2:0]    port_state_out_7_2_6,
  output     [2:0]    port_state_out_7_2_7,
  output     [2:0]    port_state_out_7_3_0,
  output     [2:0]    port_state_out_7_3_1,
  output     [2:0]    port_state_out_7_3_2,
  output     [2:0]    port_state_out_7_3_3,
  output     [2:0]    port_state_out_7_3_4,
  output     [2:0]    port_state_out_7_3_5,
  output     [2:0]    port_state_out_7_3_6,
  output     [2:0]    port_state_out_7_3_7,
  output     [2:0]    port_state_out_8_0_0,
  output     [2:0]    port_state_out_8_0_1,
  output     [2:0]    port_state_out_8_0_2,
  output     [2:0]    port_state_out_8_0_3,
  output     [2:0]    port_state_out_8_0_4,
  output     [2:0]    port_state_out_8_0_5,
  output     [2:0]    port_state_out_8_0_6,
  output     [2:0]    port_state_out_8_0_7,
  output     [2:0]    port_state_out_8_1_0,
  output     [2:0]    port_state_out_8_1_1,
  output     [2:0]    port_state_out_8_1_2,
  output     [2:0]    port_state_out_8_1_3,
  output     [2:0]    port_state_out_8_1_4,
  output     [2:0]    port_state_out_8_1_5,
  output     [2:0]    port_state_out_8_1_6,
  output     [2:0]    port_state_out_8_1_7,
  output     [2:0]    port_state_out_8_2_0,
  output     [2:0]    port_state_out_8_2_1,
  output     [2:0]    port_state_out_8_2_2,
  output     [2:0]    port_state_out_8_2_3,
  output     [2:0]    port_state_out_8_2_4,
  output     [2:0]    port_state_out_8_2_5,
  output     [2:0]    port_state_out_8_2_6,
  output     [2:0]    port_state_out_8_2_7,
  output     [2:0]    port_state_out_8_3_0,
  output     [2:0]    port_state_out_8_3_1,
  output     [2:0]    port_state_out_8_3_2,
  output     [2:0]    port_state_out_8_3_3,
  output     [2:0]    port_state_out_8_3_4,
  output     [2:0]    port_state_out_8_3_5,
  output     [2:0]    port_state_out_8_3_6,
  output     [2:0]    port_state_out_8_3_7,
  output     [2:0]    port_state_out_9_0_0,
  output     [2:0]    port_state_out_9_0_1,
  output     [2:0]    port_state_out_9_0_2,
  output     [2:0]    port_state_out_9_0_3,
  output     [2:0]    port_state_out_9_0_4,
  output     [2:0]    port_state_out_9_0_5,
  output     [2:0]    port_state_out_9_0_6,
  output     [2:0]    port_state_out_9_0_7,
  output     [2:0]    port_state_out_9_1_0,
  output     [2:0]    port_state_out_9_1_1,
  output     [2:0]    port_state_out_9_1_2,
  output     [2:0]    port_state_out_9_1_3,
  output     [2:0]    port_state_out_9_1_4,
  output     [2:0]    port_state_out_9_1_5,
  output     [2:0]    port_state_out_9_1_6,
  output     [2:0]    port_state_out_9_1_7,
  output     [2:0]    port_state_out_9_2_0,
  output     [2:0]    port_state_out_9_2_1,
  output     [2:0]    port_state_out_9_2_2,
  output     [2:0]    port_state_out_9_2_3,
  output     [2:0]    port_state_out_9_2_4,
  output     [2:0]    port_state_out_9_2_5,
  output     [2:0]    port_state_out_9_2_6,
  output     [2:0]    port_state_out_9_2_7,
  output     [2:0]    port_state_out_9_3_0,
  output     [2:0]    port_state_out_9_3_1,
  output     [2:0]    port_state_out_9_3_2,
  output     [2:0]    port_state_out_9_3_3,
  output     [2:0]    port_state_out_9_3_4,
  output     [2:0]    port_state_out_9_3_5,
  output     [2:0]    port_state_out_9_3_6,
  output     [2:0]    port_state_out_9_3_7,
  output     [2:0]    port_state_out_10_0_0,
  output     [2:0]    port_state_out_10_0_1,
  output     [2:0]    port_state_out_10_0_2,
  output     [2:0]    port_state_out_10_0_3,
  output     [2:0]    port_state_out_10_0_4,
  output     [2:0]    port_state_out_10_0_5,
  output     [2:0]    port_state_out_10_0_6,
  output     [2:0]    port_state_out_10_0_7,
  output     [2:0]    port_state_out_10_1_0,
  output     [2:0]    port_state_out_10_1_1,
  output     [2:0]    port_state_out_10_1_2,
  output     [2:0]    port_state_out_10_1_3,
  output     [2:0]    port_state_out_10_1_4,
  output     [2:0]    port_state_out_10_1_5,
  output     [2:0]    port_state_out_10_1_6,
  output     [2:0]    port_state_out_10_1_7,
  output     [2:0]    port_state_out_10_2_0,
  output     [2:0]    port_state_out_10_2_1,
  output     [2:0]    port_state_out_10_2_2,
  output     [2:0]    port_state_out_10_2_3,
  output     [2:0]    port_state_out_10_2_4,
  output     [2:0]    port_state_out_10_2_5,
  output     [2:0]    port_state_out_10_2_6,
  output     [2:0]    port_state_out_10_2_7,
  output     [2:0]    port_state_out_10_3_0,
  output     [2:0]    port_state_out_10_3_1,
  output     [2:0]    port_state_out_10_3_2,
  output     [2:0]    port_state_out_10_3_3,
  output     [2:0]    port_state_out_10_3_4,
  output     [2:0]    port_state_out_10_3_5,
  output     [2:0]    port_state_out_10_3_6,
  output     [2:0]    port_state_out_10_3_7,
  output     [2:0]    port_state_out_11_0_0,
  output     [2:0]    port_state_out_11_0_1,
  output     [2:0]    port_state_out_11_0_2,
  output     [2:0]    port_state_out_11_0_3,
  output     [2:0]    port_state_out_11_0_4,
  output     [2:0]    port_state_out_11_0_5,
  output     [2:0]    port_state_out_11_0_6,
  output     [2:0]    port_state_out_11_0_7,
  output     [2:0]    port_state_out_11_1_0,
  output     [2:0]    port_state_out_11_1_1,
  output     [2:0]    port_state_out_11_1_2,
  output     [2:0]    port_state_out_11_1_3,
  output     [2:0]    port_state_out_11_1_4,
  output     [2:0]    port_state_out_11_1_5,
  output     [2:0]    port_state_out_11_1_6,
  output     [2:0]    port_state_out_11_1_7,
  output     [2:0]    port_state_out_11_2_0,
  output     [2:0]    port_state_out_11_2_1,
  output     [2:0]    port_state_out_11_2_2,
  output     [2:0]    port_state_out_11_2_3,
  output     [2:0]    port_state_out_11_2_4,
  output     [2:0]    port_state_out_11_2_5,
  output     [2:0]    port_state_out_11_2_6,
  output     [2:0]    port_state_out_11_2_7,
  output     [2:0]    port_state_out_11_3_0,
  output     [2:0]    port_state_out_11_3_1,
  output     [2:0]    port_state_out_11_3_2,
  output     [2:0]    port_state_out_11_3_3,
  output     [2:0]    port_state_out_11_3_4,
  output     [2:0]    port_state_out_11_3_5,
  output     [2:0]    port_state_out_11_3_6,
  output     [2:0]    port_state_out_11_3_7,
  output     [2:0]    port_state_out_12_0_0,
  output     [2:0]    port_state_out_12_0_1,
  output     [2:0]    port_state_out_12_0_2,
  output     [2:0]    port_state_out_12_0_3,
  output     [2:0]    port_state_out_12_0_4,
  output     [2:0]    port_state_out_12_0_5,
  output     [2:0]    port_state_out_12_0_6,
  output     [2:0]    port_state_out_12_0_7,
  output     [2:0]    port_state_out_12_1_0,
  output     [2:0]    port_state_out_12_1_1,
  output     [2:0]    port_state_out_12_1_2,
  output     [2:0]    port_state_out_12_1_3,
  output     [2:0]    port_state_out_12_1_4,
  output     [2:0]    port_state_out_12_1_5,
  output     [2:0]    port_state_out_12_1_6,
  output     [2:0]    port_state_out_12_1_7,
  output     [2:0]    port_state_out_12_2_0,
  output     [2:0]    port_state_out_12_2_1,
  output     [2:0]    port_state_out_12_2_2,
  output     [2:0]    port_state_out_12_2_3,
  output     [2:0]    port_state_out_12_2_4,
  output     [2:0]    port_state_out_12_2_5,
  output     [2:0]    port_state_out_12_2_6,
  output     [2:0]    port_state_out_12_2_7,
  output     [2:0]    port_state_out_12_3_0,
  output     [2:0]    port_state_out_12_3_1,
  output     [2:0]    port_state_out_12_3_2,
  output     [2:0]    port_state_out_12_3_3,
  output     [2:0]    port_state_out_12_3_4,
  output     [2:0]    port_state_out_12_3_5,
  output     [2:0]    port_state_out_12_3_6,
  output     [2:0]    port_state_out_12_3_7,
  output     [2:0]    port_state_out_13_0_0,
  output     [2:0]    port_state_out_13_0_1,
  output     [2:0]    port_state_out_13_0_2,
  output     [2:0]    port_state_out_13_0_3,
  output     [2:0]    port_state_out_13_0_4,
  output     [2:0]    port_state_out_13_0_5,
  output     [2:0]    port_state_out_13_0_6,
  output     [2:0]    port_state_out_13_0_7,
  output     [2:0]    port_state_out_13_1_0,
  output     [2:0]    port_state_out_13_1_1,
  output     [2:0]    port_state_out_13_1_2,
  output     [2:0]    port_state_out_13_1_3,
  output     [2:0]    port_state_out_13_1_4,
  output     [2:0]    port_state_out_13_1_5,
  output     [2:0]    port_state_out_13_1_6,
  output     [2:0]    port_state_out_13_1_7,
  output     [2:0]    port_state_out_13_2_0,
  output     [2:0]    port_state_out_13_2_1,
  output     [2:0]    port_state_out_13_2_2,
  output     [2:0]    port_state_out_13_2_3,
  output     [2:0]    port_state_out_13_2_4,
  output     [2:0]    port_state_out_13_2_5,
  output     [2:0]    port_state_out_13_2_6,
  output     [2:0]    port_state_out_13_2_7,
  output     [2:0]    port_state_out_13_3_0,
  output     [2:0]    port_state_out_13_3_1,
  output     [2:0]    port_state_out_13_3_2,
  output     [2:0]    port_state_out_13_3_3,
  output     [2:0]    port_state_out_13_3_4,
  output     [2:0]    port_state_out_13_3_5,
  output     [2:0]    port_state_out_13_3_6,
  output     [2:0]    port_state_out_13_3_7,
  output     [2:0]    port_state_out_14_0_0,
  output     [2:0]    port_state_out_14_0_1,
  output     [2:0]    port_state_out_14_0_2,
  output     [2:0]    port_state_out_14_0_3,
  output     [2:0]    port_state_out_14_0_4,
  output     [2:0]    port_state_out_14_0_5,
  output     [2:0]    port_state_out_14_0_6,
  output     [2:0]    port_state_out_14_0_7,
  output     [2:0]    port_state_out_14_1_0,
  output     [2:0]    port_state_out_14_1_1,
  output     [2:0]    port_state_out_14_1_2,
  output     [2:0]    port_state_out_14_1_3,
  output     [2:0]    port_state_out_14_1_4,
  output     [2:0]    port_state_out_14_1_5,
  output     [2:0]    port_state_out_14_1_6,
  output     [2:0]    port_state_out_14_1_7,
  output     [2:0]    port_state_out_14_2_0,
  output     [2:0]    port_state_out_14_2_1,
  output     [2:0]    port_state_out_14_2_2,
  output     [2:0]    port_state_out_14_2_3,
  output     [2:0]    port_state_out_14_2_4,
  output     [2:0]    port_state_out_14_2_5,
  output     [2:0]    port_state_out_14_2_6,
  output     [2:0]    port_state_out_14_2_7,
  output     [2:0]    port_state_out_14_3_0,
  output     [2:0]    port_state_out_14_3_1,
  output     [2:0]    port_state_out_14_3_2,
  output     [2:0]    port_state_out_14_3_3,
  output     [2:0]    port_state_out_14_3_4,
  output     [2:0]    port_state_out_14_3_5,
  output     [2:0]    port_state_out_14_3_6,
  output     [2:0]    port_state_out_14_3_7,
  output     [2:0]    port_state_out_15_0_0,
  output     [2:0]    port_state_out_15_0_1,
  output     [2:0]    port_state_out_15_0_2,
  output     [2:0]    port_state_out_15_0_3,
  output     [2:0]    port_state_out_15_0_4,
  output     [2:0]    port_state_out_15_0_5,
  output     [2:0]    port_state_out_15_0_6,
  output     [2:0]    port_state_out_15_0_7,
  output     [2:0]    port_state_out_15_1_0,
  output     [2:0]    port_state_out_15_1_1,
  output     [2:0]    port_state_out_15_1_2,
  output     [2:0]    port_state_out_15_1_3,
  output     [2:0]    port_state_out_15_1_4,
  output     [2:0]    port_state_out_15_1_5,
  output     [2:0]    port_state_out_15_1_6,
  output     [2:0]    port_state_out_15_1_7,
  output     [2:0]    port_state_out_15_2_0,
  output     [2:0]    port_state_out_15_2_1,
  output     [2:0]    port_state_out_15_2_2,
  output     [2:0]    port_state_out_15_2_3,
  output     [2:0]    port_state_out_15_2_4,
  output     [2:0]    port_state_out_15_2_5,
  output     [2:0]    port_state_out_15_2_6,
  output     [2:0]    port_state_out_15_2_7,
  output     [2:0]    port_state_out_15_3_0,
  output     [2:0]    port_state_out_15_3_1,
  output     [2:0]    port_state_out_15_3_2,
  output     [2:0]    port_state_out_15_3_3,
  output     [2:0]    port_state_out_15_3_4,
  output     [2:0]    port_state_out_15_3_5,
  output     [2:0]    port_state_out_15_3_6,
  output     [2:0]    port_state_out_15_3_7,
  input               clk,
  input               reset
);

  wire       [2:0]    keyAdd_port_state_out_0_0_0;
  wire       [2:0]    keyAdd_port_state_out_0_0_1;
  wire       [2:0]    keyAdd_port_state_out_0_0_2;
  wire       [2:0]    keyAdd_port_state_out_0_0_3;
  wire       [2:0]    keyAdd_port_state_out_0_0_4;
  wire       [2:0]    keyAdd_port_state_out_0_0_5;
  wire       [2:0]    keyAdd_port_state_out_0_0_6;
  wire       [2:0]    keyAdd_port_state_out_0_0_7;
  wire       [2:0]    keyAdd_port_state_out_0_1_0;
  wire       [2:0]    keyAdd_port_state_out_0_1_1;
  wire       [2:0]    keyAdd_port_state_out_0_1_2;
  wire       [2:0]    keyAdd_port_state_out_0_1_3;
  wire       [2:0]    keyAdd_port_state_out_0_1_4;
  wire       [2:0]    keyAdd_port_state_out_0_1_5;
  wire       [2:0]    keyAdd_port_state_out_0_1_6;
  wire       [2:0]    keyAdd_port_state_out_0_1_7;
  wire       [2:0]    keyAdd_port_state_out_0_2_0;
  wire       [2:0]    keyAdd_port_state_out_0_2_1;
  wire       [2:0]    keyAdd_port_state_out_0_2_2;
  wire       [2:0]    keyAdd_port_state_out_0_2_3;
  wire       [2:0]    keyAdd_port_state_out_0_2_4;
  wire       [2:0]    keyAdd_port_state_out_0_2_5;
  wire       [2:0]    keyAdd_port_state_out_0_2_6;
  wire       [2:0]    keyAdd_port_state_out_0_2_7;
  wire       [2:0]    keyAdd_port_state_out_0_3_0;
  wire       [2:0]    keyAdd_port_state_out_0_3_1;
  wire       [2:0]    keyAdd_port_state_out_0_3_2;
  wire       [2:0]    keyAdd_port_state_out_0_3_3;
  wire       [2:0]    keyAdd_port_state_out_0_3_4;
  wire       [2:0]    keyAdd_port_state_out_0_3_5;
  wire       [2:0]    keyAdd_port_state_out_0_3_6;
  wire       [2:0]    keyAdd_port_state_out_0_3_7;
  wire       [2:0]    keyAdd_port_state_out_1_0_0;
  wire       [2:0]    keyAdd_port_state_out_1_0_1;
  wire       [2:0]    keyAdd_port_state_out_1_0_2;
  wire       [2:0]    keyAdd_port_state_out_1_0_3;
  wire       [2:0]    keyAdd_port_state_out_1_0_4;
  wire       [2:0]    keyAdd_port_state_out_1_0_5;
  wire       [2:0]    keyAdd_port_state_out_1_0_6;
  wire       [2:0]    keyAdd_port_state_out_1_0_7;
  wire       [2:0]    keyAdd_port_state_out_1_1_0;
  wire       [2:0]    keyAdd_port_state_out_1_1_1;
  wire       [2:0]    keyAdd_port_state_out_1_1_2;
  wire       [2:0]    keyAdd_port_state_out_1_1_3;
  wire       [2:0]    keyAdd_port_state_out_1_1_4;
  wire       [2:0]    keyAdd_port_state_out_1_1_5;
  wire       [2:0]    keyAdd_port_state_out_1_1_6;
  wire       [2:0]    keyAdd_port_state_out_1_1_7;
  wire       [2:0]    keyAdd_port_state_out_1_2_0;
  wire       [2:0]    keyAdd_port_state_out_1_2_1;
  wire       [2:0]    keyAdd_port_state_out_1_2_2;
  wire       [2:0]    keyAdd_port_state_out_1_2_3;
  wire       [2:0]    keyAdd_port_state_out_1_2_4;
  wire       [2:0]    keyAdd_port_state_out_1_2_5;
  wire       [2:0]    keyAdd_port_state_out_1_2_6;
  wire       [2:0]    keyAdd_port_state_out_1_2_7;
  wire       [2:0]    keyAdd_port_state_out_1_3_0;
  wire       [2:0]    keyAdd_port_state_out_1_3_1;
  wire       [2:0]    keyAdd_port_state_out_1_3_2;
  wire       [2:0]    keyAdd_port_state_out_1_3_3;
  wire       [2:0]    keyAdd_port_state_out_1_3_4;
  wire       [2:0]    keyAdd_port_state_out_1_3_5;
  wire       [2:0]    keyAdd_port_state_out_1_3_6;
  wire       [2:0]    keyAdd_port_state_out_1_3_7;
  wire       [2:0]    keyAdd_port_state_out_2_0_0;
  wire       [2:0]    keyAdd_port_state_out_2_0_1;
  wire       [2:0]    keyAdd_port_state_out_2_0_2;
  wire       [2:0]    keyAdd_port_state_out_2_0_3;
  wire       [2:0]    keyAdd_port_state_out_2_0_4;
  wire       [2:0]    keyAdd_port_state_out_2_0_5;
  wire       [2:0]    keyAdd_port_state_out_2_0_6;
  wire       [2:0]    keyAdd_port_state_out_2_0_7;
  wire       [2:0]    keyAdd_port_state_out_2_1_0;
  wire       [2:0]    keyAdd_port_state_out_2_1_1;
  wire       [2:0]    keyAdd_port_state_out_2_1_2;
  wire       [2:0]    keyAdd_port_state_out_2_1_3;
  wire       [2:0]    keyAdd_port_state_out_2_1_4;
  wire       [2:0]    keyAdd_port_state_out_2_1_5;
  wire       [2:0]    keyAdd_port_state_out_2_1_6;
  wire       [2:0]    keyAdd_port_state_out_2_1_7;
  wire       [2:0]    keyAdd_port_state_out_2_2_0;
  wire       [2:0]    keyAdd_port_state_out_2_2_1;
  wire       [2:0]    keyAdd_port_state_out_2_2_2;
  wire       [2:0]    keyAdd_port_state_out_2_2_3;
  wire       [2:0]    keyAdd_port_state_out_2_2_4;
  wire       [2:0]    keyAdd_port_state_out_2_2_5;
  wire       [2:0]    keyAdd_port_state_out_2_2_6;
  wire       [2:0]    keyAdd_port_state_out_2_2_7;
  wire       [2:0]    keyAdd_port_state_out_2_3_0;
  wire       [2:0]    keyAdd_port_state_out_2_3_1;
  wire       [2:0]    keyAdd_port_state_out_2_3_2;
  wire       [2:0]    keyAdd_port_state_out_2_3_3;
  wire       [2:0]    keyAdd_port_state_out_2_3_4;
  wire       [2:0]    keyAdd_port_state_out_2_3_5;
  wire       [2:0]    keyAdd_port_state_out_2_3_6;
  wire       [2:0]    keyAdd_port_state_out_2_3_7;
  wire       [2:0]    keyAdd_port_state_out_3_0_0;
  wire       [2:0]    keyAdd_port_state_out_3_0_1;
  wire       [2:0]    keyAdd_port_state_out_3_0_2;
  wire       [2:0]    keyAdd_port_state_out_3_0_3;
  wire       [2:0]    keyAdd_port_state_out_3_0_4;
  wire       [2:0]    keyAdd_port_state_out_3_0_5;
  wire       [2:0]    keyAdd_port_state_out_3_0_6;
  wire       [2:0]    keyAdd_port_state_out_3_0_7;
  wire       [2:0]    keyAdd_port_state_out_3_1_0;
  wire       [2:0]    keyAdd_port_state_out_3_1_1;
  wire       [2:0]    keyAdd_port_state_out_3_1_2;
  wire       [2:0]    keyAdd_port_state_out_3_1_3;
  wire       [2:0]    keyAdd_port_state_out_3_1_4;
  wire       [2:0]    keyAdd_port_state_out_3_1_5;
  wire       [2:0]    keyAdd_port_state_out_3_1_6;
  wire       [2:0]    keyAdd_port_state_out_3_1_7;
  wire       [2:0]    keyAdd_port_state_out_3_2_0;
  wire       [2:0]    keyAdd_port_state_out_3_2_1;
  wire       [2:0]    keyAdd_port_state_out_3_2_2;
  wire       [2:0]    keyAdd_port_state_out_3_2_3;
  wire       [2:0]    keyAdd_port_state_out_3_2_4;
  wire       [2:0]    keyAdd_port_state_out_3_2_5;
  wire       [2:0]    keyAdd_port_state_out_3_2_6;
  wire       [2:0]    keyAdd_port_state_out_3_2_7;
  wire       [2:0]    keyAdd_port_state_out_3_3_0;
  wire       [2:0]    keyAdd_port_state_out_3_3_1;
  wire       [2:0]    keyAdd_port_state_out_3_3_2;
  wire       [2:0]    keyAdd_port_state_out_3_3_3;
  wire       [2:0]    keyAdd_port_state_out_3_3_4;
  wire       [2:0]    keyAdd_port_state_out_3_3_5;
  wire       [2:0]    keyAdd_port_state_out_3_3_6;
  wire       [2:0]    keyAdd_port_state_out_3_3_7;
  wire       [2:0]    keyAdd_port_state_out_4_0_0;
  wire       [2:0]    keyAdd_port_state_out_4_0_1;
  wire       [2:0]    keyAdd_port_state_out_4_0_2;
  wire       [2:0]    keyAdd_port_state_out_4_0_3;
  wire       [2:0]    keyAdd_port_state_out_4_0_4;
  wire       [2:0]    keyAdd_port_state_out_4_0_5;
  wire       [2:0]    keyAdd_port_state_out_4_0_6;
  wire       [2:0]    keyAdd_port_state_out_4_0_7;
  wire       [2:0]    keyAdd_port_state_out_4_1_0;
  wire       [2:0]    keyAdd_port_state_out_4_1_1;
  wire       [2:0]    keyAdd_port_state_out_4_1_2;
  wire       [2:0]    keyAdd_port_state_out_4_1_3;
  wire       [2:0]    keyAdd_port_state_out_4_1_4;
  wire       [2:0]    keyAdd_port_state_out_4_1_5;
  wire       [2:0]    keyAdd_port_state_out_4_1_6;
  wire       [2:0]    keyAdd_port_state_out_4_1_7;
  wire       [2:0]    keyAdd_port_state_out_4_2_0;
  wire       [2:0]    keyAdd_port_state_out_4_2_1;
  wire       [2:0]    keyAdd_port_state_out_4_2_2;
  wire       [2:0]    keyAdd_port_state_out_4_2_3;
  wire       [2:0]    keyAdd_port_state_out_4_2_4;
  wire       [2:0]    keyAdd_port_state_out_4_2_5;
  wire       [2:0]    keyAdd_port_state_out_4_2_6;
  wire       [2:0]    keyAdd_port_state_out_4_2_7;
  wire       [2:0]    keyAdd_port_state_out_4_3_0;
  wire       [2:0]    keyAdd_port_state_out_4_3_1;
  wire       [2:0]    keyAdd_port_state_out_4_3_2;
  wire       [2:0]    keyAdd_port_state_out_4_3_3;
  wire       [2:0]    keyAdd_port_state_out_4_3_4;
  wire       [2:0]    keyAdd_port_state_out_4_3_5;
  wire       [2:0]    keyAdd_port_state_out_4_3_6;
  wire       [2:0]    keyAdd_port_state_out_4_3_7;
  wire       [2:0]    keyAdd_port_state_out_5_0_0;
  wire       [2:0]    keyAdd_port_state_out_5_0_1;
  wire       [2:0]    keyAdd_port_state_out_5_0_2;
  wire       [2:0]    keyAdd_port_state_out_5_0_3;
  wire       [2:0]    keyAdd_port_state_out_5_0_4;
  wire       [2:0]    keyAdd_port_state_out_5_0_5;
  wire       [2:0]    keyAdd_port_state_out_5_0_6;
  wire       [2:0]    keyAdd_port_state_out_5_0_7;
  wire       [2:0]    keyAdd_port_state_out_5_1_0;
  wire       [2:0]    keyAdd_port_state_out_5_1_1;
  wire       [2:0]    keyAdd_port_state_out_5_1_2;
  wire       [2:0]    keyAdd_port_state_out_5_1_3;
  wire       [2:0]    keyAdd_port_state_out_5_1_4;
  wire       [2:0]    keyAdd_port_state_out_5_1_5;
  wire       [2:0]    keyAdd_port_state_out_5_1_6;
  wire       [2:0]    keyAdd_port_state_out_5_1_7;
  wire       [2:0]    keyAdd_port_state_out_5_2_0;
  wire       [2:0]    keyAdd_port_state_out_5_2_1;
  wire       [2:0]    keyAdd_port_state_out_5_2_2;
  wire       [2:0]    keyAdd_port_state_out_5_2_3;
  wire       [2:0]    keyAdd_port_state_out_5_2_4;
  wire       [2:0]    keyAdd_port_state_out_5_2_5;
  wire       [2:0]    keyAdd_port_state_out_5_2_6;
  wire       [2:0]    keyAdd_port_state_out_5_2_7;
  wire       [2:0]    keyAdd_port_state_out_5_3_0;
  wire       [2:0]    keyAdd_port_state_out_5_3_1;
  wire       [2:0]    keyAdd_port_state_out_5_3_2;
  wire       [2:0]    keyAdd_port_state_out_5_3_3;
  wire       [2:0]    keyAdd_port_state_out_5_3_4;
  wire       [2:0]    keyAdd_port_state_out_5_3_5;
  wire       [2:0]    keyAdd_port_state_out_5_3_6;
  wire       [2:0]    keyAdd_port_state_out_5_3_7;
  wire       [2:0]    keyAdd_port_state_out_6_0_0;
  wire       [2:0]    keyAdd_port_state_out_6_0_1;
  wire       [2:0]    keyAdd_port_state_out_6_0_2;
  wire       [2:0]    keyAdd_port_state_out_6_0_3;
  wire       [2:0]    keyAdd_port_state_out_6_0_4;
  wire       [2:0]    keyAdd_port_state_out_6_0_5;
  wire       [2:0]    keyAdd_port_state_out_6_0_6;
  wire       [2:0]    keyAdd_port_state_out_6_0_7;
  wire       [2:0]    keyAdd_port_state_out_6_1_0;
  wire       [2:0]    keyAdd_port_state_out_6_1_1;
  wire       [2:0]    keyAdd_port_state_out_6_1_2;
  wire       [2:0]    keyAdd_port_state_out_6_1_3;
  wire       [2:0]    keyAdd_port_state_out_6_1_4;
  wire       [2:0]    keyAdd_port_state_out_6_1_5;
  wire       [2:0]    keyAdd_port_state_out_6_1_6;
  wire       [2:0]    keyAdd_port_state_out_6_1_7;
  wire       [2:0]    keyAdd_port_state_out_6_2_0;
  wire       [2:0]    keyAdd_port_state_out_6_2_1;
  wire       [2:0]    keyAdd_port_state_out_6_2_2;
  wire       [2:0]    keyAdd_port_state_out_6_2_3;
  wire       [2:0]    keyAdd_port_state_out_6_2_4;
  wire       [2:0]    keyAdd_port_state_out_6_2_5;
  wire       [2:0]    keyAdd_port_state_out_6_2_6;
  wire       [2:0]    keyAdd_port_state_out_6_2_7;
  wire       [2:0]    keyAdd_port_state_out_6_3_0;
  wire       [2:0]    keyAdd_port_state_out_6_3_1;
  wire       [2:0]    keyAdd_port_state_out_6_3_2;
  wire       [2:0]    keyAdd_port_state_out_6_3_3;
  wire       [2:0]    keyAdd_port_state_out_6_3_4;
  wire       [2:0]    keyAdd_port_state_out_6_3_5;
  wire       [2:0]    keyAdd_port_state_out_6_3_6;
  wire       [2:0]    keyAdd_port_state_out_6_3_7;
  wire       [2:0]    keyAdd_port_state_out_7_0_0;
  wire       [2:0]    keyAdd_port_state_out_7_0_1;
  wire       [2:0]    keyAdd_port_state_out_7_0_2;
  wire       [2:0]    keyAdd_port_state_out_7_0_3;
  wire       [2:0]    keyAdd_port_state_out_7_0_4;
  wire       [2:0]    keyAdd_port_state_out_7_0_5;
  wire       [2:0]    keyAdd_port_state_out_7_0_6;
  wire       [2:0]    keyAdd_port_state_out_7_0_7;
  wire       [2:0]    keyAdd_port_state_out_7_1_0;
  wire       [2:0]    keyAdd_port_state_out_7_1_1;
  wire       [2:0]    keyAdd_port_state_out_7_1_2;
  wire       [2:0]    keyAdd_port_state_out_7_1_3;
  wire       [2:0]    keyAdd_port_state_out_7_1_4;
  wire       [2:0]    keyAdd_port_state_out_7_1_5;
  wire       [2:0]    keyAdd_port_state_out_7_1_6;
  wire       [2:0]    keyAdd_port_state_out_7_1_7;
  wire       [2:0]    keyAdd_port_state_out_7_2_0;
  wire       [2:0]    keyAdd_port_state_out_7_2_1;
  wire       [2:0]    keyAdd_port_state_out_7_2_2;
  wire       [2:0]    keyAdd_port_state_out_7_2_3;
  wire       [2:0]    keyAdd_port_state_out_7_2_4;
  wire       [2:0]    keyAdd_port_state_out_7_2_5;
  wire       [2:0]    keyAdd_port_state_out_7_2_6;
  wire       [2:0]    keyAdd_port_state_out_7_2_7;
  wire       [2:0]    keyAdd_port_state_out_7_3_0;
  wire       [2:0]    keyAdd_port_state_out_7_3_1;
  wire       [2:0]    keyAdd_port_state_out_7_3_2;
  wire       [2:0]    keyAdd_port_state_out_7_3_3;
  wire       [2:0]    keyAdd_port_state_out_7_3_4;
  wire       [2:0]    keyAdd_port_state_out_7_3_5;
  wire       [2:0]    keyAdd_port_state_out_7_3_6;
  wire       [2:0]    keyAdd_port_state_out_7_3_7;
  wire       [2:0]    keyAdd_port_state_out_8_0_0;
  wire       [2:0]    keyAdd_port_state_out_8_0_1;
  wire       [2:0]    keyAdd_port_state_out_8_0_2;
  wire       [2:0]    keyAdd_port_state_out_8_0_3;
  wire       [2:0]    keyAdd_port_state_out_8_0_4;
  wire       [2:0]    keyAdd_port_state_out_8_0_5;
  wire       [2:0]    keyAdd_port_state_out_8_0_6;
  wire       [2:0]    keyAdd_port_state_out_8_0_7;
  wire       [2:0]    keyAdd_port_state_out_8_1_0;
  wire       [2:0]    keyAdd_port_state_out_8_1_1;
  wire       [2:0]    keyAdd_port_state_out_8_1_2;
  wire       [2:0]    keyAdd_port_state_out_8_1_3;
  wire       [2:0]    keyAdd_port_state_out_8_1_4;
  wire       [2:0]    keyAdd_port_state_out_8_1_5;
  wire       [2:0]    keyAdd_port_state_out_8_1_6;
  wire       [2:0]    keyAdd_port_state_out_8_1_7;
  wire       [2:0]    keyAdd_port_state_out_8_2_0;
  wire       [2:0]    keyAdd_port_state_out_8_2_1;
  wire       [2:0]    keyAdd_port_state_out_8_2_2;
  wire       [2:0]    keyAdd_port_state_out_8_2_3;
  wire       [2:0]    keyAdd_port_state_out_8_2_4;
  wire       [2:0]    keyAdd_port_state_out_8_2_5;
  wire       [2:0]    keyAdd_port_state_out_8_2_6;
  wire       [2:0]    keyAdd_port_state_out_8_2_7;
  wire       [2:0]    keyAdd_port_state_out_8_3_0;
  wire       [2:0]    keyAdd_port_state_out_8_3_1;
  wire       [2:0]    keyAdd_port_state_out_8_3_2;
  wire       [2:0]    keyAdd_port_state_out_8_3_3;
  wire       [2:0]    keyAdd_port_state_out_8_3_4;
  wire       [2:0]    keyAdd_port_state_out_8_3_5;
  wire       [2:0]    keyAdd_port_state_out_8_3_6;
  wire       [2:0]    keyAdd_port_state_out_8_3_7;
  wire       [2:0]    keyAdd_port_state_out_9_0_0;
  wire       [2:0]    keyAdd_port_state_out_9_0_1;
  wire       [2:0]    keyAdd_port_state_out_9_0_2;
  wire       [2:0]    keyAdd_port_state_out_9_0_3;
  wire       [2:0]    keyAdd_port_state_out_9_0_4;
  wire       [2:0]    keyAdd_port_state_out_9_0_5;
  wire       [2:0]    keyAdd_port_state_out_9_0_6;
  wire       [2:0]    keyAdd_port_state_out_9_0_7;
  wire       [2:0]    keyAdd_port_state_out_9_1_0;
  wire       [2:0]    keyAdd_port_state_out_9_1_1;
  wire       [2:0]    keyAdd_port_state_out_9_1_2;
  wire       [2:0]    keyAdd_port_state_out_9_1_3;
  wire       [2:0]    keyAdd_port_state_out_9_1_4;
  wire       [2:0]    keyAdd_port_state_out_9_1_5;
  wire       [2:0]    keyAdd_port_state_out_9_1_6;
  wire       [2:0]    keyAdd_port_state_out_9_1_7;
  wire       [2:0]    keyAdd_port_state_out_9_2_0;
  wire       [2:0]    keyAdd_port_state_out_9_2_1;
  wire       [2:0]    keyAdd_port_state_out_9_2_2;
  wire       [2:0]    keyAdd_port_state_out_9_2_3;
  wire       [2:0]    keyAdd_port_state_out_9_2_4;
  wire       [2:0]    keyAdd_port_state_out_9_2_5;
  wire       [2:0]    keyAdd_port_state_out_9_2_6;
  wire       [2:0]    keyAdd_port_state_out_9_2_7;
  wire       [2:0]    keyAdd_port_state_out_9_3_0;
  wire       [2:0]    keyAdd_port_state_out_9_3_1;
  wire       [2:0]    keyAdd_port_state_out_9_3_2;
  wire       [2:0]    keyAdd_port_state_out_9_3_3;
  wire       [2:0]    keyAdd_port_state_out_9_3_4;
  wire       [2:0]    keyAdd_port_state_out_9_3_5;
  wire       [2:0]    keyAdd_port_state_out_9_3_6;
  wire       [2:0]    keyAdd_port_state_out_9_3_7;
  wire       [2:0]    keyAdd_port_state_out_10_0_0;
  wire       [2:0]    keyAdd_port_state_out_10_0_1;
  wire       [2:0]    keyAdd_port_state_out_10_0_2;
  wire       [2:0]    keyAdd_port_state_out_10_0_3;
  wire       [2:0]    keyAdd_port_state_out_10_0_4;
  wire       [2:0]    keyAdd_port_state_out_10_0_5;
  wire       [2:0]    keyAdd_port_state_out_10_0_6;
  wire       [2:0]    keyAdd_port_state_out_10_0_7;
  wire       [2:0]    keyAdd_port_state_out_10_1_0;
  wire       [2:0]    keyAdd_port_state_out_10_1_1;
  wire       [2:0]    keyAdd_port_state_out_10_1_2;
  wire       [2:0]    keyAdd_port_state_out_10_1_3;
  wire       [2:0]    keyAdd_port_state_out_10_1_4;
  wire       [2:0]    keyAdd_port_state_out_10_1_5;
  wire       [2:0]    keyAdd_port_state_out_10_1_6;
  wire       [2:0]    keyAdd_port_state_out_10_1_7;
  wire       [2:0]    keyAdd_port_state_out_10_2_0;
  wire       [2:0]    keyAdd_port_state_out_10_2_1;
  wire       [2:0]    keyAdd_port_state_out_10_2_2;
  wire       [2:0]    keyAdd_port_state_out_10_2_3;
  wire       [2:0]    keyAdd_port_state_out_10_2_4;
  wire       [2:0]    keyAdd_port_state_out_10_2_5;
  wire       [2:0]    keyAdd_port_state_out_10_2_6;
  wire       [2:0]    keyAdd_port_state_out_10_2_7;
  wire       [2:0]    keyAdd_port_state_out_10_3_0;
  wire       [2:0]    keyAdd_port_state_out_10_3_1;
  wire       [2:0]    keyAdd_port_state_out_10_3_2;
  wire       [2:0]    keyAdd_port_state_out_10_3_3;
  wire       [2:0]    keyAdd_port_state_out_10_3_4;
  wire       [2:0]    keyAdd_port_state_out_10_3_5;
  wire       [2:0]    keyAdd_port_state_out_10_3_6;
  wire       [2:0]    keyAdd_port_state_out_10_3_7;
  wire       [2:0]    keyAdd_port_state_out_11_0_0;
  wire       [2:0]    keyAdd_port_state_out_11_0_1;
  wire       [2:0]    keyAdd_port_state_out_11_0_2;
  wire       [2:0]    keyAdd_port_state_out_11_0_3;
  wire       [2:0]    keyAdd_port_state_out_11_0_4;
  wire       [2:0]    keyAdd_port_state_out_11_0_5;
  wire       [2:0]    keyAdd_port_state_out_11_0_6;
  wire       [2:0]    keyAdd_port_state_out_11_0_7;
  wire       [2:0]    keyAdd_port_state_out_11_1_0;
  wire       [2:0]    keyAdd_port_state_out_11_1_1;
  wire       [2:0]    keyAdd_port_state_out_11_1_2;
  wire       [2:0]    keyAdd_port_state_out_11_1_3;
  wire       [2:0]    keyAdd_port_state_out_11_1_4;
  wire       [2:0]    keyAdd_port_state_out_11_1_5;
  wire       [2:0]    keyAdd_port_state_out_11_1_6;
  wire       [2:0]    keyAdd_port_state_out_11_1_7;
  wire       [2:0]    keyAdd_port_state_out_11_2_0;
  wire       [2:0]    keyAdd_port_state_out_11_2_1;
  wire       [2:0]    keyAdd_port_state_out_11_2_2;
  wire       [2:0]    keyAdd_port_state_out_11_2_3;
  wire       [2:0]    keyAdd_port_state_out_11_2_4;
  wire       [2:0]    keyAdd_port_state_out_11_2_5;
  wire       [2:0]    keyAdd_port_state_out_11_2_6;
  wire       [2:0]    keyAdd_port_state_out_11_2_7;
  wire       [2:0]    keyAdd_port_state_out_11_3_0;
  wire       [2:0]    keyAdd_port_state_out_11_3_1;
  wire       [2:0]    keyAdd_port_state_out_11_3_2;
  wire       [2:0]    keyAdd_port_state_out_11_3_3;
  wire       [2:0]    keyAdd_port_state_out_11_3_4;
  wire       [2:0]    keyAdd_port_state_out_11_3_5;
  wire       [2:0]    keyAdd_port_state_out_11_3_6;
  wire       [2:0]    keyAdd_port_state_out_11_3_7;
  wire       [2:0]    keyAdd_port_state_out_12_0_0;
  wire       [2:0]    keyAdd_port_state_out_12_0_1;
  wire       [2:0]    keyAdd_port_state_out_12_0_2;
  wire       [2:0]    keyAdd_port_state_out_12_0_3;
  wire       [2:0]    keyAdd_port_state_out_12_0_4;
  wire       [2:0]    keyAdd_port_state_out_12_0_5;
  wire       [2:0]    keyAdd_port_state_out_12_0_6;
  wire       [2:0]    keyAdd_port_state_out_12_0_7;
  wire       [2:0]    keyAdd_port_state_out_12_1_0;
  wire       [2:0]    keyAdd_port_state_out_12_1_1;
  wire       [2:0]    keyAdd_port_state_out_12_1_2;
  wire       [2:0]    keyAdd_port_state_out_12_1_3;
  wire       [2:0]    keyAdd_port_state_out_12_1_4;
  wire       [2:0]    keyAdd_port_state_out_12_1_5;
  wire       [2:0]    keyAdd_port_state_out_12_1_6;
  wire       [2:0]    keyAdd_port_state_out_12_1_7;
  wire       [2:0]    keyAdd_port_state_out_12_2_0;
  wire       [2:0]    keyAdd_port_state_out_12_2_1;
  wire       [2:0]    keyAdd_port_state_out_12_2_2;
  wire       [2:0]    keyAdd_port_state_out_12_2_3;
  wire       [2:0]    keyAdd_port_state_out_12_2_4;
  wire       [2:0]    keyAdd_port_state_out_12_2_5;
  wire       [2:0]    keyAdd_port_state_out_12_2_6;
  wire       [2:0]    keyAdd_port_state_out_12_2_7;
  wire       [2:0]    keyAdd_port_state_out_12_3_0;
  wire       [2:0]    keyAdd_port_state_out_12_3_1;
  wire       [2:0]    keyAdd_port_state_out_12_3_2;
  wire       [2:0]    keyAdd_port_state_out_12_3_3;
  wire       [2:0]    keyAdd_port_state_out_12_3_4;
  wire       [2:0]    keyAdd_port_state_out_12_3_5;
  wire       [2:0]    keyAdd_port_state_out_12_3_6;
  wire       [2:0]    keyAdd_port_state_out_12_3_7;
  wire       [2:0]    keyAdd_port_state_out_13_0_0;
  wire       [2:0]    keyAdd_port_state_out_13_0_1;
  wire       [2:0]    keyAdd_port_state_out_13_0_2;
  wire       [2:0]    keyAdd_port_state_out_13_0_3;
  wire       [2:0]    keyAdd_port_state_out_13_0_4;
  wire       [2:0]    keyAdd_port_state_out_13_0_5;
  wire       [2:0]    keyAdd_port_state_out_13_0_6;
  wire       [2:0]    keyAdd_port_state_out_13_0_7;
  wire       [2:0]    keyAdd_port_state_out_13_1_0;
  wire       [2:0]    keyAdd_port_state_out_13_1_1;
  wire       [2:0]    keyAdd_port_state_out_13_1_2;
  wire       [2:0]    keyAdd_port_state_out_13_1_3;
  wire       [2:0]    keyAdd_port_state_out_13_1_4;
  wire       [2:0]    keyAdd_port_state_out_13_1_5;
  wire       [2:0]    keyAdd_port_state_out_13_1_6;
  wire       [2:0]    keyAdd_port_state_out_13_1_7;
  wire       [2:0]    keyAdd_port_state_out_13_2_0;
  wire       [2:0]    keyAdd_port_state_out_13_2_1;
  wire       [2:0]    keyAdd_port_state_out_13_2_2;
  wire       [2:0]    keyAdd_port_state_out_13_2_3;
  wire       [2:0]    keyAdd_port_state_out_13_2_4;
  wire       [2:0]    keyAdd_port_state_out_13_2_5;
  wire       [2:0]    keyAdd_port_state_out_13_2_6;
  wire       [2:0]    keyAdd_port_state_out_13_2_7;
  wire       [2:0]    keyAdd_port_state_out_13_3_0;
  wire       [2:0]    keyAdd_port_state_out_13_3_1;
  wire       [2:0]    keyAdd_port_state_out_13_3_2;
  wire       [2:0]    keyAdd_port_state_out_13_3_3;
  wire       [2:0]    keyAdd_port_state_out_13_3_4;
  wire       [2:0]    keyAdd_port_state_out_13_3_5;
  wire       [2:0]    keyAdd_port_state_out_13_3_6;
  wire       [2:0]    keyAdd_port_state_out_13_3_7;
  wire       [2:0]    keyAdd_port_state_out_14_0_0;
  wire       [2:0]    keyAdd_port_state_out_14_0_1;
  wire       [2:0]    keyAdd_port_state_out_14_0_2;
  wire       [2:0]    keyAdd_port_state_out_14_0_3;
  wire       [2:0]    keyAdd_port_state_out_14_0_4;
  wire       [2:0]    keyAdd_port_state_out_14_0_5;
  wire       [2:0]    keyAdd_port_state_out_14_0_6;
  wire       [2:0]    keyAdd_port_state_out_14_0_7;
  wire       [2:0]    keyAdd_port_state_out_14_1_0;
  wire       [2:0]    keyAdd_port_state_out_14_1_1;
  wire       [2:0]    keyAdd_port_state_out_14_1_2;
  wire       [2:0]    keyAdd_port_state_out_14_1_3;
  wire       [2:0]    keyAdd_port_state_out_14_1_4;
  wire       [2:0]    keyAdd_port_state_out_14_1_5;
  wire       [2:0]    keyAdd_port_state_out_14_1_6;
  wire       [2:0]    keyAdd_port_state_out_14_1_7;
  wire       [2:0]    keyAdd_port_state_out_14_2_0;
  wire       [2:0]    keyAdd_port_state_out_14_2_1;
  wire       [2:0]    keyAdd_port_state_out_14_2_2;
  wire       [2:0]    keyAdd_port_state_out_14_2_3;
  wire       [2:0]    keyAdd_port_state_out_14_2_4;
  wire       [2:0]    keyAdd_port_state_out_14_2_5;
  wire       [2:0]    keyAdd_port_state_out_14_2_6;
  wire       [2:0]    keyAdd_port_state_out_14_2_7;
  wire       [2:0]    keyAdd_port_state_out_14_3_0;
  wire       [2:0]    keyAdd_port_state_out_14_3_1;
  wire       [2:0]    keyAdd_port_state_out_14_3_2;
  wire       [2:0]    keyAdd_port_state_out_14_3_3;
  wire       [2:0]    keyAdd_port_state_out_14_3_4;
  wire       [2:0]    keyAdd_port_state_out_14_3_5;
  wire       [2:0]    keyAdd_port_state_out_14_3_6;
  wire       [2:0]    keyAdd_port_state_out_14_3_7;
  wire       [2:0]    keyAdd_port_state_out_15_0_0;
  wire       [2:0]    keyAdd_port_state_out_15_0_1;
  wire       [2:0]    keyAdd_port_state_out_15_0_2;
  wire       [2:0]    keyAdd_port_state_out_15_0_3;
  wire       [2:0]    keyAdd_port_state_out_15_0_4;
  wire       [2:0]    keyAdd_port_state_out_15_0_5;
  wire       [2:0]    keyAdd_port_state_out_15_0_6;
  wire       [2:0]    keyAdd_port_state_out_15_0_7;
  wire       [2:0]    keyAdd_port_state_out_15_1_0;
  wire       [2:0]    keyAdd_port_state_out_15_1_1;
  wire       [2:0]    keyAdd_port_state_out_15_1_2;
  wire       [2:0]    keyAdd_port_state_out_15_1_3;
  wire       [2:0]    keyAdd_port_state_out_15_1_4;
  wire       [2:0]    keyAdd_port_state_out_15_1_5;
  wire       [2:0]    keyAdd_port_state_out_15_1_6;
  wire       [2:0]    keyAdd_port_state_out_15_1_7;
  wire       [2:0]    keyAdd_port_state_out_15_2_0;
  wire       [2:0]    keyAdd_port_state_out_15_2_1;
  wire       [2:0]    keyAdd_port_state_out_15_2_2;
  wire       [2:0]    keyAdd_port_state_out_15_2_3;
  wire       [2:0]    keyAdd_port_state_out_15_2_4;
  wire       [2:0]    keyAdd_port_state_out_15_2_5;
  wire       [2:0]    keyAdd_port_state_out_15_2_6;
  wire       [2:0]    keyAdd_port_state_out_15_2_7;
  wire       [2:0]    keyAdd_port_state_out_15_3_0;
  wire       [2:0]    keyAdd_port_state_out_15_3_1;
  wire       [2:0]    keyAdd_port_state_out_15_3_2;
  wire       [2:0]    keyAdd_port_state_out_15_3_3;
  wire       [2:0]    keyAdd_port_state_out_15_3_4;
  wire       [2:0]    keyAdd_port_state_out_15_3_5;
  wire       [2:0]    keyAdd_port_state_out_15_3_6;
  wire       [2:0]    keyAdd_port_state_out_15_3_7;
  wire       [2:0]    sbox_AES_BoyarPeralta_16_port_o_0_0;
  wire       [2:0]    sbox_AES_BoyarPeralta_16_port_o_0_1;
  wire       [2:0]    sbox_AES_BoyarPeralta_16_port_o_0_2;
  wire       [2:0]    sbox_AES_BoyarPeralta_16_port_o_0_3;
  wire       [2:0]    sbox_AES_BoyarPeralta_16_port_o_0_4;
  wire       [2:0]    sbox_AES_BoyarPeralta_16_port_o_0_5;
  wire       [2:0]    sbox_AES_BoyarPeralta_16_port_o_0_6;
  wire       [2:0]    sbox_AES_BoyarPeralta_16_port_o_0_7;
  wire       [2:0]    sbox_AES_BoyarPeralta_16_port_o_1_0;
  wire       [2:0]    sbox_AES_BoyarPeralta_16_port_o_1_1;
  wire       [2:0]    sbox_AES_BoyarPeralta_16_port_o_1_2;
  wire       [2:0]    sbox_AES_BoyarPeralta_16_port_o_1_3;
  wire       [2:0]    sbox_AES_BoyarPeralta_16_port_o_1_4;
  wire       [2:0]    sbox_AES_BoyarPeralta_16_port_o_1_5;
  wire       [2:0]    sbox_AES_BoyarPeralta_16_port_o_1_6;
  wire       [2:0]    sbox_AES_BoyarPeralta_16_port_o_1_7;
  wire       [2:0]    sbox_AES_BoyarPeralta_16_port_o_2_0;
  wire       [2:0]    sbox_AES_BoyarPeralta_16_port_o_2_1;
  wire       [2:0]    sbox_AES_BoyarPeralta_16_port_o_2_2;
  wire       [2:0]    sbox_AES_BoyarPeralta_16_port_o_2_3;
  wire       [2:0]    sbox_AES_BoyarPeralta_16_port_o_2_4;
  wire       [2:0]    sbox_AES_BoyarPeralta_16_port_o_2_5;
  wire       [2:0]    sbox_AES_BoyarPeralta_16_port_o_2_6;
  wire       [2:0]    sbox_AES_BoyarPeralta_16_port_o_2_7;
  wire       [2:0]    sbox_AES_BoyarPeralta_16_port_o_3_0;
  wire       [2:0]    sbox_AES_BoyarPeralta_16_port_o_3_1;
  wire       [2:0]    sbox_AES_BoyarPeralta_16_port_o_3_2;
  wire       [2:0]    sbox_AES_BoyarPeralta_16_port_o_3_3;
  wire       [2:0]    sbox_AES_BoyarPeralta_16_port_o_3_4;
  wire       [2:0]    sbox_AES_BoyarPeralta_16_port_o_3_5;
  wire       [2:0]    sbox_AES_BoyarPeralta_16_port_o_3_6;
  wire       [2:0]    sbox_AES_BoyarPeralta_16_port_o_3_7;
  wire       [2:0]    sbox_AES_BoyarPeralta_17_port_o_0_0;
  wire       [2:0]    sbox_AES_BoyarPeralta_17_port_o_0_1;
  wire       [2:0]    sbox_AES_BoyarPeralta_17_port_o_0_2;
  wire       [2:0]    sbox_AES_BoyarPeralta_17_port_o_0_3;
  wire       [2:0]    sbox_AES_BoyarPeralta_17_port_o_0_4;
  wire       [2:0]    sbox_AES_BoyarPeralta_17_port_o_0_5;
  wire       [2:0]    sbox_AES_BoyarPeralta_17_port_o_0_6;
  wire       [2:0]    sbox_AES_BoyarPeralta_17_port_o_0_7;
  wire       [2:0]    sbox_AES_BoyarPeralta_17_port_o_1_0;
  wire       [2:0]    sbox_AES_BoyarPeralta_17_port_o_1_1;
  wire       [2:0]    sbox_AES_BoyarPeralta_17_port_o_1_2;
  wire       [2:0]    sbox_AES_BoyarPeralta_17_port_o_1_3;
  wire       [2:0]    sbox_AES_BoyarPeralta_17_port_o_1_4;
  wire       [2:0]    sbox_AES_BoyarPeralta_17_port_o_1_5;
  wire       [2:0]    sbox_AES_BoyarPeralta_17_port_o_1_6;
  wire       [2:0]    sbox_AES_BoyarPeralta_17_port_o_1_7;
  wire       [2:0]    sbox_AES_BoyarPeralta_17_port_o_2_0;
  wire       [2:0]    sbox_AES_BoyarPeralta_17_port_o_2_1;
  wire       [2:0]    sbox_AES_BoyarPeralta_17_port_o_2_2;
  wire       [2:0]    sbox_AES_BoyarPeralta_17_port_o_2_3;
  wire       [2:0]    sbox_AES_BoyarPeralta_17_port_o_2_4;
  wire       [2:0]    sbox_AES_BoyarPeralta_17_port_o_2_5;
  wire       [2:0]    sbox_AES_BoyarPeralta_17_port_o_2_6;
  wire       [2:0]    sbox_AES_BoyarPeralta_17_port_o_2_7;
  wire       [2:0]    sbox_AES_BoyarPeralta_17_port_o_3_0;
  wire       [2:0]    sbox_AES_BoyarPeralta_17_port_o_3_1;
  wire       [2:0]    sbox_AES_BoyarPeralta_17_port_o_3_2;
  wire       [2:0]    sbox_AES_BoyarPeralta_17_port_o_3_3;
  wire       [2:0]    sbox_AES_BoyarPeralta_17_port_o_3_4;
  wire       [2:0]    sbox_AES_BoyarPeralta_17_port_o_3_5;
  wire       [2:0]    sbox_AES_BoyarPeralta_17_port_o_3_6;
  wire       [2:0]    sbox_AES_BoyarPeralta_17_port_o_3_7;
  wire       [2:0]    sbox_AES_BoyarPeralta_18_port_o_0_0;
  wire       [2:0]    sbox_AES_BoyarPeralta_18_port_o_0_1;
  wire       [2:0]    sbox_AES_BoyarPeralta_18_port_o_0_2;
  wire       [2:0]    sbox_AES_BoyarPeralta_18_port_o_0_3;
  wire       [2:0]    sbox_AES_BoyarPeralta_18_port_o_0_4;
  wire       [2:0]    sbox_AES_BoyarPeralta_18_port_o_0_5;
  wire       [2:0]    sbox_AES_BoyarPeralta_18_port_o_0_6;
  wire       [2:0]    sbox_AES_BoyarPeralta_18_port_o_0_7;
  wire       [2:0]    sbox_AES_BoyarPeralta_18_port_o_1_0;
  wire       [2:0]    sbox_AES_BoyarPeralta_18_port_o_1_1;
  wire       [2:0]    sbox_AES_BoyarPeralta_18_port_o_1_2;
  wire       [2:0]    sbox_AES_BoyarPeralta_18_port_o_1_3;
  wire       [2:0]    sbox_AES_BoyarPeralta_18_port_o_1_4;
  wire       [2:0]    sbox_AES_BoyarPeralta_18_port_o_1_5;
  wire       [2:0]    sbox_AES_BoyarPeralta_18_port_o_1_6;
  wire       [2:0]    sbox_AES_BoyarPeralta_18_port_o_1_7;
  wire       [2:0]    sbox_AES_BoyarPeralta_18_port_o_2_0;
  wire       [2:0]    sbox_AES_BoyarPeralta_18_port_o_2_1;
  wire       [2:0]    sbox_AES_BoyarPeralta_18_port_o_2_2;
  wire       [2:0]    sbox_AES_BoyarPeralta_18_port_o_2_3;
  wire       [2:0]    sbox_AES_BoyarPeralta_18_port_o_2_4;
  wire       [2:0]    sbox_AES_BoyarPeralta_18_port_o_2_5;
  wire       [2:0]    sbox_AES_BoyarPeralta_18_port_o_2_6;
  wire       [2:0]    sbox_AES_BoyarPeralta_18_port_o_2_7;
  wire       [2:0]    sbox_AES_BoyarPeralta_18_port_o_3_0;
  wire       [2:0]    sbox_AES_BoyarPeralta_18_port_o_3_1;
  wire       [2:0]    sbox_AES_BoyarPeralta_18_port_o_3_2;
  wire       [2:0]    sbox_AES_BoyarPeralta_18_port_o_3_3;
  wire       [2:0]    sbox_AES_BoyarPeralta_18_port_o_3_4;
  wire       [2:0]    sbox_AES_BoyarPeralta_18_port_o_3_5;
  wire       [2:0]    sbox_AES_BoyarPeralta_18_port_o_3_6;
  wire       [2:0]    sbox_AES_BoyarPeralta_18_port_o_3_7;
  wire       [2:0]    sbox_AES_BoyarPeralta_19_port_o_0_0;
  wire       [2:0]    sbox_AES_BoyarPeralta_19_port_o_0_1;
  wire       [2:0]    sbox_AES_BoyarPeralta_19_port_o_0_2;
  wire       [2:0]    sbox_AES_BoyarPeralta_19_port_o_0_3;
  wire       [2:0]    sbox_AES_BoyarPeralta_19_port_o_0_4;
  wire       [2:0]    sbox_AES_BoyarPeralta_19_port_o_0_5;
  wire       [2:0]    sbox_AES_BoyarPeralta_19_port_o_0_6;
  wire       [2:0]    sbox_AES_BoyarPeralta_19_port_o_0_7;
  wire       [2:0]    sbox_AES_BoyarPeralta_19_port_o_1_0;
  wire       [2:0]    sbox_AES_BoyarPeralta_19_port_o_1_1;
  wire       [2:0]    sbox_AES_BoyarPeralta_19_port_o_1_2;
  wire       [2:0]    sbox_AES_BoyarPeralta_19_port_o_1_3;
  wire       [2:0]    sbox_AES_BoyarPeralta_19_port_o_1_4;
  wire       [2:0]    sbox_AES_BoyarPeralta_19_port_o_1_5;
  wire       [2:0]    sbox_AES_BoyarPeralta_19_port_o_1_6;
  wire       [2:0]    sbox_AES_BoyarPeralta_19_port_o_1_7;
  wire       [2:0]    sbox_AES_BoyarPeralta_19_port_o_2_0;
  wire       [2:0]    sbox_AES_BoyarPeralta_19_port_o_2_1;
  wire       [2:0]    sbox_AES_BoyarPeralta_19_port_o_2_2;
  wire       [2:0]    sbox_AES_BoyarPeralta_19_port_o_2_3;
  wire       [2:0]    sbox_AES_BoyarPeralta_19_port_o_2_4;
  wire       [2:0]    sbox_AES_BoyarPeralta_19_port_o_2_5;
  wire       [2:0]    sbox_AES_BoyarPeralta_19_port_o_2_6;
  wire       [2:0]    sbox_AES_BoyarPeralta_19_port_o_2_7;
  wire       [2:0]    sbox_AES_BoyarPeralta_19_port_o_3_0;
  wire       [2:0]    sbox_AES_BoyarPeralta_19_port_o_3_1;
  wire       [2:0]    sbox_AES_BoyarPeralta_19_port_o_3_2;
  wire       [2:0]    sbox_AES_BoyarPeralta_19_port_o_3_3;
  wire       [2:0]    sbox_AES_BoyarPeralta_19_port_o_3_4;
  wire       [2:0]    sbox_AES_BoyarPeralta_19_port_o_3_5;
  wire       [2:0]    sbox_AES_BoyarPeralta_19_port_o_3_6;
  wire       [2:0]    sbox_AES_BoyarPeralta_19_port_o_3_7;
  wire       [2:0]    sbox_AES_BoyarPeralta_20_port_o_0_0;
  wire       [2:0]    sbox_AES_BoyarPeralta_20_port_o_0_1;
  wire       [2:0]    sbox_AES_BoyarPeralta_20_port_o_0_2;
  wire       [2:0]    sbox_AES_BoyarPeralta_20_port_o_0_3;
  wire       [2:0]    sbox_AES_BoyarPeralta_20_port_o_0_4;
  wire       [2:0]    sbox_AES_BoyarPeralta_20_port_o_0_5;
  wire       [2:0]    sbox_AES_BoyarPeralta_20_port_o_0_6;
  wire       [2:0]    sbox_AES_BoyarPeralta_20_port_o_0_7;
  wire       [2:0]    sbox_AES_BoyarPeralta_20_port_o_1_0;
  wire       [2:0]    sbox_AES_BoyarPeralta_20_port_o_1_1;
  wire       [2:0]    sbox_AES_BoyarPeralta_20_port_o_1_2;
  wire       [2:0]    sbox_AES_BoyarPeralta_20_port_o_1_3;
  wire       [2:0]    sbox_AES_BoyarPeralta_20_port_o_1_4;
  wire       [2:0]    sbox_AES_BoyarPeralta_20_port_o_1_5;
  wire       [2:0]    sbox_AES_BoyarPeralta_20_port_o_1_6;
  wire       [2:0]    sbox_AES_BoyarPeralta_20_port_o_1_7;
  wire       [2:0]    sbox_AES_BoyarPeralta_20_port_o_2_0;
  wire       [2:0]    sbox_AES_BoyarPeralta_20_port_o_2_1;
  wire       [2:0]    sbox_AES_BoyarPeralta_20_port_o_2_2;
  wire       [2:0]    sbox_AES_BoyarPeralta_20_port_o_2_3;
  wire       [2:0]    sbox_AES_BoyarPeralta_20_port_o_2_4;
  wire       [2:0]    sbox_AES_BoyarPeralta_20_port_o_2_5;
  wire       [2:0]    sbox_AES_BoyarPeralta_20_port_o_2_6;
  wire       [2:0]    sbox_AES_BoyarPeralta_20_port_o_2_7;
  wire       [2:0]    sbox_AES_BoyarPeralta_20_port_o_3_0;
  wire       [2:0]    sbox_AES_BoyarPeralta_20_port_o_3_1;
  wire       [2:0]    sbox_AES_BoyarPeralta_20_port_o_3_2;
  wire       [2:0]    sbox_AES_BoyarPeralta_20_port_o_3_3;
  wire       [2:0]    sbox_AES_BoyarPeralta_20_port_o_3_4;
  wire       [2:0]    sbox_AES_BoyarPeralta_20_port_o_3_5;
  wire       [2:0]    sbox_AES_BoyarPeralta_20_port_o_3_6;
  wire       [2:0]    sbox_AES_BoyarPeralta_20_port_o_3_7;
  wire       [2:0]    sbox_AES_BoyarPeralta_21_port_o_0_0;
  wire       [2:0]    sbox_AES_BoyarPeralta_21_port_o_0_1;
  wire       [2:0]    sbox_AES_BoyarPeralta_21_port_o_0_2;
  wire       [2:0]    sbox_AES_BoyarPeralta_21_port_o_0_3;
  wire       [2:0]    sbox_AES_BoyarPeralta_21_port_o_0_4;
  wire       [2:0]    sbox_AES_BoyarPeralta_21_port_o_0_5;
  wire       [2:0]    sbox_AES_BoyarPeralta_21_port_o_0_6;
  wire       [2:0]    sbox_AES_BoyarPeralta_21_port_o_0_7;
  wire       [2:0]    sbox_AES_BoyarPeralta_21_port_o_1_0;
  wire       [2:0]    sbox_AES_BoyarPeralta_21_port_o_1_1;
  wire       [2:0]    sbox_AES_BoyarPeralta_21_port_o_1_2;
  wire       [2:0]    sbox_AES_BoyarPeralta_21_port_o_1_3;
  wire       [2:0]    sbox_AES_BoyarPeralta_21_port_o_1_4;
  wire       [2:0]    sbox_AES_BoyarPeralta_21_port_o_1_5;
  wire       [2:0]    sbox_AES_BoyarPeralta_21_port_o_1_6;
  wire       [2:0]    sbox_AES_BoyarPeralta_21_port_o_1_7;
  wire       [2:0]    sbox_AES_BoyarPeralta_21_port_o_2_0;
  wire       [2:0]    sbox_AES_BoyarPeralta_21_port_o_2_1;
  wire       [2:0]    sbox_AES_BoyarPeralta_21_port_o_2_2;
  wire       [2:0]    sbox_AES_BoyarPeralta_21_port_o_2_3;
  wire       [2:0]    sbox_AES_BoyarPeralta_21_port_o_2_4;
  wire       [2:0]    sbox_AES_BoyarPeralta_21_port_o_2_5;
  wire       [2:0]    sbox_AES_BoyarPeralta_21_port_o_2_6;
  wire       [2:0]    sbox_AES_BoyarPeralta_21_port_o_2_7;
  wire       [2:0]    sbox_AES_BoyarPeralta_21_port_o_3_0;
  wire       [2:0]    sbox_AES_BoyarPeralta_21_port_o_3_1;
  wire       [2:0]    sbox_AES_BoyarPeralta_21_port_o_3_2;
  wire       [2:0]    sbox_AES_BoyarPeralta_21_port_o_3_3;
  wire       [2:0]    sbox_AES_BoyarPeralta_21_port_o_3_4;
  wire       [2:0]    sbox_AES_BoyarPeralta_21_port_o_3_5;
  wire       [2:0]    sbox_AES_BoyarPeralta_21_port_o_3_6;
  wire       [2:0]    sbox_AES_BoyarPeralta_21_port_o_3_7;
  wire       [2:0]    sbox_AES_BoyarPeralta_22_port_o_0_0;
  wire       [2:0]    sbox_AES_BoyarPeralta_22_port_o_0_1;
  wire       [2:0]    sbox_AES_BoyarPeralta_22_port_o_0_2;
  wire       [2:0]    sbox_AES_BoyarPeralta_22_port_o_0_3;
  wire       [2:0]    sbox_AES_BoyarPeralta_22_port_o_0_4;
  wire       [2:0]    sbox_AES_BoyarPeralta_22_port_o_0_5;
  wire       [2:0]    sbox_AES_BoyarPeralta_22_port_o_0_6;
  wire       [2:0]    sbox_AES_BoyarPeralta_22_port_o_0_7;
  wire       [2:0]    sbox_AES_BoyarPeralta_22_port_o_1_0;
  wire       [2:0]    sbox_AES_BoyarPeralta_22_port_o_1_1;
  wire       [2:0]    sbox_AES_BoyarPeralta_22_port_o_1_2;
  wire       [2:0]    sbox_AES_BoyarPeralta_22_port_o_1_3;
  wire       [2:0]    sbox_AES_BoyarPeralta_22_port_o_1_4;
  wire       [2:0]    sbox_AES_BoyarPeralta_22_port_o_1_5;
  wire       [2:0]    sbox_AES_BoyarPeralta_22_port_o_1_6;
  wire       [2:0]    sbox_AES_BoyarPeralta_22_port_o_1_7;
  wire       [2:0]    sbox_AES_BoyarPeralta_22_port_o_2_0;
  wire       [2:0]    sbox_AES_BoyarPeralta_22_port_o_2_1;
  wire       [2:0]    sbox_AES_BoyarPeralta_22_port_o_2_2;
  wire       [2:0]    sbox_AES_BoyarPeralta_22_port_o_2_3;
  wire       [2:0]    sbox_AES_BoyarPeralta_22_port_o_2_4;
  wire       [2:0]    sbox_AES_BoyarPeralta_22_port_o_2_5;
  wire       [2:0]    sbox_AES_BoyarPeralta_22_port_o_2_6;
  wire       [2:0]    sbox_AES_BoyarPeralta_22_port_o_2_7;
  wire       [2:0]    sbox_AES_BoyarPeralta_22_port_o_3_0;
  wire       [2:0]    sbox_AES_BoyarPeralta_22_port_o_3_1;
  wire       [2:0]    sbox_AES_BoyarPeralta_22_port_o_3_2;
  wire       [2:0]    sbox_AES_BoyarPeralta_22_port_o_3_3;
  wire       [2:0]    sbox_AES_BoyarPeralta_22_port_o_3_4;
  wire       [2:0]    sbox_AES_BoyarPeralta_22_port_o_3_5;
  wire       [2:0]    sbox_AES_BoyarPeralta_22_port_o_3_6;
  wire       [2:0]    sbox_AES_BoyarPeralta_22_port_o_3_7;
  wire       [2:0]    sbox_AES_BoyarPeralta_23_port_o_0_0;
  wire       [2:0]    sbox_AES_BoyarPeralta_23_port_o_0_1;
  wire       [2:0]    sbox_AES_BoyarPeralta_23_port_o_0_2;
  wire       [2:0]    sbox_AES_BoyarPeralta_23_port_o_0_3;
  wire       [2:0]    sbox_AES_BoyarPeralta_23_port_o_0_4;
  wire       [2:0]    sbox_AES_BoyarPeralta_23_port_o_0_5;
  wire       [2:0]    sbox_AES_BoyarPeralta_23_port_o_0_6;
  wire       [2:0]    sbox_AES_BoyarPeralta_23_port_o_0_7;
  wire       [2:0]    sbox_AES_BoyarPeralta_23_port_o_1_0;
  wire       [2:0]    sbox_AES_BoyarPeralta_23_port_o_1_1;
  wire       [2:0]    sbox_AES_BoyarPeralta_23_port_o_1_2;
  wire       [2:0]    sbox_AES_BoyarPeralta_23_port_o_1_3;
  wire       [2:0]    sbox_AES_BoyarPeralta_23_port_o_1_4;
  wire       [2:0]    sbox_AES_BoyarPeralta_23_port_o_1_5;
  wire       [2:0]    sbox_AES_BoyarPeralta_23_port_o_1_6;
  wire       [2:0]    sbox_AES_BoyarPeralta_23_port_o_1_7;
  wire       [2:0]    sbox_AES_BoyarPeralta_23_port_o_2_0;
  wire       [2:0]    sbox_AES_BoyarPeralta_23_port_o_2_1;
  wire       [2:0]    sbox_AES_BoyarPeralta_23_port_o_2_2;
  wire       [2:0]    sbox_AES_BoyarPeralta_23_port_o_2_3;
  wire       [2:0]    sbox_AES_BoyarPeralta_23_port_o_2_4;
  wire       [2:0]    sbox_AES_BoyarPeralta_23_port_o_2_5;
  wire       [2:0]    sbox_AES_BoyarPeralta_23_port_o_2_6;
  wire       [2:0]    sbox_AES_BoyarPeralta_23_port_o_2_7;
  wire       [2:0]    sbox_AES_BoyarPeralta_23_port_o_3_0;
  wire       [2:0]    sbox_AES_BoyarPeralta_23_port_o_3_1;
  wire       [2:0]    sbox_AES_BoyarPeralta_23_port_o_3_2;
  wire       [2:0]    sbox_AES_BoyarPeralta_23_port_o_3_3;
  wire       [2:0]    sbox_AES_BoyarPeralta_23_port_o_3_4;
  wire       [2:0]    sbox_AES_BoyarPeralta_23_port_o_3_5;
  wire       [2:0]    sbox_AES_BoyarPeralta_23_port_o_3_6;
  wire       [2:0]    sbox_AES_BoyarPeralta_23_port_o_3_7;
  wire       [2:0]    sbox_AES_BoyarPeralta_24_port_o_0_0;
  wire       [2:0]    sbox_AES_BoyarPeralta_24_port_o_0_1;
  wire       [2:0]    sbox_AES_BoyarPeralta_24_port_o_0_2;
  wire       [2:0]    sbox_AES_BoyarPeralta_24_port_o_0_3;
  wire       [2:0]    sbox_AES_BoyarPeralta_24_port_o_0_4;
  wire       [2:0]    sbox_AES_BoyarPeralta_24_port_o_0_5;
  wire       [2:0]    sbox_AES_BoyarPeralta_24_port_o_0_6;
  wire       [2:0]    sbox_AES_BoyarPeralta_24_port_o_0_7;
  wire       [2:0]    sbox_AES_BoyarPeralta_24_port_o_1_0;
  wire       [2:0]    sbox_AES_BoyarPeralta_24_port_o_1_1;
  wire       [2:0]    sbox_AES_BoyarPeralta_24_port_o_1_2;
  wire       [2:0]    sbox_AES_BoyarPeralta_24_port_o_1_3;
  wire       [2:0]    sbox_AES_BoyarPeralta_24_port_o_1_4;
  wire       [2:0]    sbox_AES_BoyarPeralta_24_port_o_1_5;
  wire       [2:0]    sbox_AES_BoyarPeralta_24_port_o_1_6;
  wire       [2:0]    sbox_AES_BoyarPeralta_24_port_o_1_7;
  wire       [2:0]    sbox_AES_BoyarPeralta_24_port_o_2_0;
  wire       [2:0]    sbox_AES_BoyarPeralta_24_port_o_2_1;
  wire       [2:0]    sbox_AES_BoyarPeralta_24_port_o_2_2;
  wire       [2:0]    sbox_AES_BoyarPeralta_24_port_o_2_3;
  wire       [2:0]    sbox_AES_BoyarPeralta_24_port_o_2_4;
  wire       [2:0]    sbox_AES_BoyarPeralta_24_port_o_2_5;
  wire       [2:0]    sbox_AES_BoyarPeralta_24_port_o_2_6;
  wire       [2:0]    sbox_AES_BoyarPeralta_24_port_o_2_7;
  wire       [2:0]    sbox_AES_BoyarPeralta_24_port_o_3_0;
  wire       [2:0]    sbox_AES_BoyarPeralta_24_port_o_3_1;
  wire       [2:0]    sbox_AES_BoyarPeralta_24_port_o_3_2;
  wire       [2:0]    sbox_AES_BoyarPeralta_24_port_o_3_3;
  wire       [2:0]    sbox_AES_BoyarPeralta_24_port_o_3_4;
  wire       [2:0]    sbox_AES_BoyarPeralta_24_port_o_3_5;
  wire       [2:0]    sbox_AES_BoyarPeralta_24_port_o_3_6;
  wire       [2:0]    sbox_AES_BoyarPeralta_24_port_o_3_7;
  wire       [2:0]    sbox_AES_BoyarPeralta_25_port_o_0_0;
  wire       [2:0]    sbox_AES_BoyarPeralta_25_port_o_0_1;
  wire       [2:0]    sbox_AES_BoyarPeralta_25_port_o_0_2;
  wire       [2:0]    sbox_AES_BoyarPeralta_25_port_o_0_3;
  wire       [2:0]    sbox_AES_BoyarPeralta_25_port_o_0_4;
  wire       [2:0]    sbox_AES_BoyarPeralta_25_port_o_0_5;
  wire       [2:0]    sbox_AES_BoyarPeralta_25_port_o_0_6;
  wire       [2:0]    sbox_AES_BoyarPeralta_25_port_o_0_7;
  wire       [2:0]    sbox_AES_BoyarPeralta_25_port_o_1_0;
  wire       [2:0]    sbox_AES_BoyarPeralta_25_port_o_1_1;
  wire       [2:0]    sbox_AES_BoyarPeralta_25_port_o_1_2;
  wire       [2:0]    sbox_AES_BoyarPeralta_25_port_o_1_3;
  wire       [2:0]    sbox_AES_BoyarPeralta_25_port_o_1_4;
  wire       [2:0]    sbox_AES_BoyarPeralta_25_port_o_1_5;
  wire       [2:0]    sbox_AES_BoyarPeralta_25_port_o_1_6;
  wire       [2:0]    sbox_AES_BoyarPeralta_25_port_o_1_7;
  wire       [2:0]    sbox_AES_BoyarPeralta_25_port_o_2_0;
  wire       [2:0]    sbox_AES_BoyarPeralta_25_port_o_2_1;
  wire       [2:0]    sbox_AES_BoyarPeralta_25_port_o_2_2;
  wire       [2:0]    sbox_AES_BoyarPeralta_25_port_o_2_3;
  wire       [2:0]    sbox_AES_BoyarPeralta_25_port_o_2_4;
  wire       [2:0]    sbox_AES_BoyarPeralta_25_port_o_2_5;
  wire       [2:0]    sbox_AES_BoyarPeralta_25_port_o_2_6;
  wire       [2:0]    sbox_AES_BoyarPeralta_25_port_o_2_7;
  wire       [2:0]    sbox_AES_BoyarPeralta_25_port_o_3_0;
  wire       [2:0]    sbox_AES_BoyarPeralta_25_port_o_3_1;
  wire       [2:0]    sbox_AES_BoyarPeralta_25_port_o_3_2;
  wire       [2:0]    sbox_AES_BoyarPeralta_25_port_o_3_3;
  wire       [2:0]    sbox_AES_BoyarPeralta_25_port_o_3_4;
  wire       [2:0]    sbox_AES_BoyarPeralta_25_port_o_3_5;
  wire       [2:0]    sbox_AES_BoyarPeralta_25_port_o_3_6;
  wire       [2:0]    sbox_AES_BoyarPeralta_25_port_o_3_7;
  wire       [2:0]    sbox_AES_BoyarPeralta_26_port_o_0_0;
  wire       [2:0]    sbox_AES_BoyarPeralta_26_port_o_0_1;
  wire       [2:0]    sbox_AES_BoyarPeralta_26_port_o_0_2;
  wire       [2:0]    sbox_AES_BoyarPeralta_26_port_o_0_3;
  wire       [2:0]    sbox_AES_BoyarPeralta_26_port_o_0_4;
  wire       [2:0]    sbox_AES_BoyarPeralta_26_port_o_0_5;
  wire       [2:0]    sbox_AES_BoyarPeralta_26_port_o_0_6;
  wire       [2:0]    sbox_AES_BoyarPeralta_26_port_o_0_7;
  wire       [2:0]    sbox_AES_BoyarPeralta_26_port_o_1_0;
  wire       [2:0]    sbox_AES_BoyarPeralta_26_port_o_1_1;
  wire       [2:0]    sbox_AES_BoyarPeralta_26_port_o_1_2;
  wire       [2:0]    sbox_AES_BoyarPeralta_26_port_o_1_3;
  wire       [2:0]    sbox_AES_BoyarPeralta_26_port_o_1_4;
  wire       [2:0]    sbox_AES_BoyarPeralta_26_port_o_1_5;
  wire       [2:0]    sbox_AES_BoyarPeralta_26_port_o_1_6;
  wire       [2:0]    sbox_AES_BoyarPeralta_26_port_o_1_7;
  wire       [2:0]    sbox_AES_BoyarPeralta_26_port_o_2_0;
  wire       [2:0]    sbox_AES_BoyarPeralta_26_port_o_2_1;
  wire       [2:0]    sbox_AES_BoyarPeralta_26_port_o_2_2;
  wire       [2:0]    sbox_AES_BoyarPeralta_26_port_o_2_3;
  wire       [2:0]    sbox_AES_BoyarPeralta_26_port_o_2_4;
  wire       [2:0]    sbox_AES_BoyarPeralta_26_port_o_2_5;
  wire       [2:0]    sbox_AES_BoyarPeralta_26_port_o_2_6;
  wire       [2:0]    sbox_AES_BoyarPeralta_26_port_o_2_7;
  wire       [2:0]    sbox_AES_BoyarPeralta_26_port_o_3_0;
  wire       [2:0]    sbox_AES_BoyarPeralta_26_port_o_3_1;
  wire       [2:0]    sbox_AES_BoyarPeralta_26_port_o_3_2;
  wire       [2:0]    sbox_AES_BoyarPeralta_26_port_o_3_3;
  wire       [2:0]    sbox_AES_BoyarPeralta_26_port_o_3_4;
  wire       [2:0]    sbox_AES_BoyarPeralta_26_port_o_3_5;
  wire       [2:0]    sbox_AES_BoyarPeralta_26_port_o_3_6;
  wire       [2:0]    sbox_AES_BoyarPeralta_26_port_o_3_7;
  wire       [2:0]    sbox_AES_BoyarPeralta_27_port_o_0_0;
  wire       [2:0]    sbox_AES_BoyarPeralta_27_port_o_0_1;
  wire       [2:0]    sbox_AES_BoyarPeralta_27_port_o_0_2;
  wire       [2:0]    sbox_AES_BoyarPeralta_27_port_o_0_3;
  wire       [2:0]    sbox_AES_BoyarPeralta_27_port_o_0_4;
  wire       [2:0]    sbox_AES_BoyarPeralta_27_port_o_0_5;
  wire       [2:0]    sbox_AES_BoyarPeralta_27_port_o_0_6;
  wire       [2:0]    sbox_AES_BoyarPeralta_27_port_o_0_7;
  wire       [2:0]    sbox_AES_BoyarPeralta_27_port_o_1_0;
  wire       [2:0]    sbox_AES_BoyarPeralta_27_port_o_1_1;
  wire       [2:0]    sbox_AES_BoyarPeralta_27_port_o_1_2;
  wire       [2:0]    sbox_AES_BoyarPeralta_27_port_o_1_3;
  wire       [2:0]    sbox_AES_BoyarPeralta_27_port_o_1_4;
  wire       [2:0]    sbox_AES_BoyarPeralta_27_port_o_1_5;
  wire       [2:0]    sbox_AES_BoyarPeralta_27_port_o_1_6;
  wire       [2:0]    sbox_AES_BoyarPeralta_27_port_o_1_7;
  wire       [2:0]    sbox_AES_BoyarPeralta_27_port_o_2_0;
  wire       [2:0]    sbox_AES_BoyarPeralta_27_port_o_2_1;
  wire       [2:0]    sbox_AES_BoyarPeralta_27_port_o_2_2;
  wire       [2:0]    sbox_AES_BoyarPeralta_27_port_o_2_3;
  wire       [2:0]    sbox_AES_BoyarPeralta_27_port_o_2_4;
  wire       [2:0]    sbox_AES_BoyarPeralta_27_port_o_2_5;
  wire       [2:0]    sbox_AES_BoyarPeralta_27_port_o_2_6;
  wire       [2:0]    sbox_AES_BoyarPeralta_27_port_o_2_7;
  wire       [2:0]    sbox_AES_BoyarPeralta_27_port_o_3_0;
  wire       [2:0]    sbox_AES_BoyarPeralta_27_port_o_3_1;
  wire       [2:0]    sbox_AES_BoyarPeralta_27_port_o_3_2;
  wire       [2:0]    sbox_AES_BoyarPeralta_27_port_o_3_3;
  wire       [2:0]    sbox_AES_BoyarPeralta_27_port_o_3_4;
  wire       [2:0]    sbox_AES_BoyarPeralta_27_port_o_3_5;
  wire       [2:0]    sbox_AES_BoyarPeralta_27_port_o_3_6;
  wire       [2:0]    sbox_AES_BoyarPeralta_27_port_o_3_7;
  wire       [2:0]    sbox_AES_BoyarPeralta_28_port_o_0_0;
  wire       [2:0]    sbox_AES_BoyarPeralta_28_port_o_0_1;
  wire       [2:0]    sbox_AES_BoyarPeralta_28_port_o_0_2;
  wire       [2:0]    sbox_AES_BoyarPeralta_28_port_o_0_3;
  wire       [2:0]    sbox_AES_BoyarPeralta_28_port_o_0_4;
  wire       [2:0]    sbox_AES_BoyarPeralta_28_port_o_0_5;
  wire       [2:0]    sbox_AES_BoyarPeralta_28_port_o_0_6;
  wire       [2:0]    sbox_AES_BoyarPeralta_28_port_o_0_7;
  wire       [2:0]    sbox_AES_BoyarPeralta_28_port_o_1_0;
  wire       [2:0]    sbox_AES_BoyarPeralta_28_port_o_1_1;
  wire       [2:0]    sbox_AES_BoyarPeralta_28_port_o_1_2;
  wire       [2:0]    sbox_AES_BoyarPeralta_28_port_o_1_3;
  wire       [2:0]    sbox_AES_BoyarPeralta_28_port_o_1_4;
  wire       [2:0]    sbox_AES_BoyarPeralta_28_port_o_1_5;
  wire       [2:0]    sbox_AES_BoyarPeralta_28_port_o_1_6;
  wire       [2:0]    sbox_AES_BoyarPeralta_28_port_o_1_7;
  wire       [2:0]    sbox_AES_BoyarPeralta_28_port_o_2_0;
  wire       [2:0]    sbox_AES_BoyarPeralta_28_port_o_2_1;
  wire       [2:0]    sbox_AES_BoyarPeralta_28_port_o_2_2;
  wire       [2:0]    sbox_AES_BoyarPeralta_28_port_o_2_3;
  wire       [2:0]    sbox_AES_BoyarPeralta_28_port_o_2_4;
  wire       [2:0]    sbox_AES_BoyarPeralta_28_port_o_2_5;
  wire       [2:0]    sbox_AES_BoyarPeralta_28_port_o_2_6;
  wire       [2:0]    sbox_AES_BoyarPeralta_28_port_o_2_7;
  wire       [2:0]    sbox_AES_BoyarPeralta_28_port_o_3_0;
  wire       [2:0]    sbox_AES_BoyarPeralta_28_port_o_3_1;
  wire       [2:0]    sbox_AES_BoyarPeralta_28_port_o_3_2;
  wire       [2:0]    sbox_AES_BoyarPeralta_28_port_o_3_3;
  wire       [2:0]    sbox_AES_BoyarPeralta_28_port_o_3_4;
  wire       [2:0]    sbox_AES_BoyarPeralta_28_port_o_3_5;
  wire       [2:0]    sbox_AES_BoyarPeralta_28_port_o_3_6;
  wire       [2:0]    sbox_AES_BoyarPeralta_28_port_o_3_7;
  wire       [2:0]    sbox_AES_BoyarPeralta_29_port_o_0_0;
  wire       [2:0]    sbox_AES_BoyarPeralta_29_port_o_0_1;
  wire       [2:0]    sbox_AES_BoyarPeralta_29_port_o_0_2;
  wire       [2:0]    sbox_AES_BoyarPeralta_29_port_o_0_3;
  wire       [2:0]    sbox_AES_BoyarPeralta_29_port_o_0_4;
  wire       [2:0]    sbox_AES_BoyarPeralta_29_port_o_0_5;
  wire       [2:0]    sbox_AES_BoyarPeralta_29_port_o_0_6;
  wire       [2:0]    sbox_AES_BoyarPeralta_29_port_o_0_7;
  wire       [2:0]    sbox_AES_BoyarPeralta_29_port_o_1_0;
  wire       [2:0]    sbox_AES_BoyarPeralta_29_port_o_1_1;
  wire       [2:0]    sbox_AES_BoyarPeralta_29_port_o_1_2;
  wire       [2:0]    sbox_AES_BoyarPeralta_29_port_o_1_3;
  wire       [2:0]    sbox_AES_BoyarPeralta_29_port_o_1_4;
  wire       [2:0]    sbox_AES_BoyarPeralta_29_port_o_1_5;
  wire       [2:0]    sbox_AES_BoyarPeralta_29_port_o_1_6;
  wire       [2:0]    sbox_AES_BoyarPeralta_29_port_o_1_7;
  wire       [2:0]    sbox_AES_BoyarPeralta_29_port_o_2_0;
  wire       [2:0]    sbox_AES_BoyarPeralta_29_port_o_2_1;
  wire       [2:0]    sbox_AES_BoyarPeralta_29_port_o_2_2;
  wire       [2:0]    sbox_AES_BoyarPeralta_29_port_o_2_3;
  wire       [2:0]    sbox_AES_BoyarPeralta_29_port_o_2_4;
  wire       [2:0]    sbox_AES_BoyarPeralta_29_port_o_2_5;
  wire       [2:0]    sbox_AES_BoyarPeralta_29_port_o_2_6;
  wire       [2:0]    sbox_AES_BoyarPeralta_29_port_o_2_7;
  wire       [2:0]    sbox_AES_BoyarPeralta_29_port_o_3_0;
  wire       [2:0]    sbox_AES_BoyarPeralta_29_port_o_3_1;
  wire       [2:0]    sbox_AES_BoyarPeralta_29_port_o_3_2;
  wire       [2:0]    sbox_AES_BoyarPeralta_29_port_o_3_3;
  wire       [2:0]    sbox_AES_BoyarPeralta_29_port_o_3_4;
  wire       [2:0]    sbox_AES_BoyarPeralta_29_port_o_3_5;
  wire       [2:0]    sbox_AES_BoyarPeralta_29_port_o_3_6;
  wire       [2:0]    sbox_AES_BoyarPeralta_29_port_o_3_7;
  wire       [2:0]    sbox_AES_BoyarPeralta_30_port_o_0_0;
  wire       [2:0]    sbox_AES_BoyarPeralta_30_port_o_0_1;
  wire       [2:0]    sbox_AES_BoyarPeralta_30_port_o_0_2;
  wire       [2:0]    sbox_AES_BoyarPeralta_30_port_o_0_3;
  wire       [2:0]    sbox_AES_BoyarPeralta_30_port_o_0_4;
  wire       [2:0]    sbox_AES_BoyarPeralta_30_port_o_0_5;
  wire       [2:0]    sbox_AES_BoyarPeralta_30_port_o_0_6;
  wire       [2:0]    sbox_AES_BoyarPeralta_30_port_o_0_7;
  wire       [2:0]    sbox_AES_BoyarPeralta_30_port_o_1_0;
  wire       [2:0]    sbox_AES_BoyarPeralta_30_port_o_1_1;
  wire       [2:0]    sbox_AES_BoyarPeralta_30_port_o_1_2;
  wire       [2:0]    sbox_AES_BoyarPeralta_30_port_o_1_3;
  wire       [2:0]    sbox_AES_BoyarPeralta_30_port_o_1_4;
  wire       [2:0]    sbox_AES_BoyarPeralta_30_port_o_1_5;
  wire       [2:0]    sbox_AES_BoyarPeralta_30_port_o_1_6;
  wire       [2:0]    sbox_AES_BoyarPeralta_30_port_o_1_7;
  wire       [2:0]    sbox_AES_BoyarPeralta_30_port_o_2_0;
  wire       [2:0]    sbox_AES_BoyarPeralta_30_port_o_2_1;
  wire       [2:0]    sbox_AES_BoyarPeralta_30_port_o_2_2;
  wire       [2:0]    sbox_AES_BoyarPeralta_30_port_o_2_3;
  wire       [2:0]    sbox_AES_BoyarPeralta_30_port_o_2_4;
  wire       [2:0]    sbox_AES_BoyarPeralta_30_port_o_2_5;
  wire       [2:0]    sbox_AES_BoyarPeralta_30_port_o_2_6;
  wire       [2:0]    sbox_AES_BoyarPeralta_30_port_o_2_7;
  wire       [2:0]    sbox_AES_BoyarPeralta_30_port_o_3_0;
  wire       [2:0]    sbox_AES_BoyarPeralta_30_port_o_3_1;
  wire       [2:0]    sbox_AES_BoyarPeralta_30_port_o_3_2;
  wire       [2:0]    sbox_AES_BoyarPeralta_30_port_o_3_3;
  wire       [2:0]    sbox_AES_BoyarPeralta_30_port_o_3_4;
  wire       [2:0]    sbox_AES_BoyarPeralta_30_port_o_3_5;
  wire       [2:0]    sbox_AES_BoyarPeralta_30_port_o_3_6;
  wire       [2:0]    sbox_AES_BoyarPeralta_30_port_o_3_7;
  wire       [2:0]    sbox_AES_BoyarPeralta_31_port_o_0_0;
  wire       [2:0]    sbox_AES_BoyarPeralta_31_port_o_0_1;
  wire       [2:0]    sbox_AES_BoyarPeralta_31_port_o_0_2;
  wire       [2:0]    sbox_AES_BoyarPeralta_31_port_o_0_3;
  wire       [2:0]    sbox_AES_BoyarPeralta_31_port_o_0_4;
  wire       [2:0]    sbox_AES_BoyarPeralta_31_port_o_0_5;
  wire       [2:0]    sbox_AES_BoyarPeralta_31_port_o_0_6;
  wire       [2:0]    sbox_AES_BoyarPeralta_31_port_o_0_7;
  wire       [2:0]    sbox_AES_BoyarPeralta_31_port_o_1_0;
  wire       [2:0]    sbox_AES_BoyarPeralta_31_port_o_1_1;
  wire       [2:0]    sbox_AES_BoyarPeralta_31_port_o_1_2;
  wire       [2:0]    sbox_AES_BoyarPeralta_31_port_o_1_3;
  wire       [2:0]    sbox_AES_BoyarPeralta_31_port_o_1_4;
  wire       [2:0]    sbox_AES_BoyarPeralta_31_port_o_1_5;
  wire       [2:0]    sbox_AES_BoyarPeralta_31_port_o_1_6;
  wire       [2:0]    sbox_AES_BoyarPeralta_31_port_o_1_7;
  wire       [2:0]    sbox_AES_BoyarPeralta_31_port_o_2_0;
  wire       [2:0]    sbox_AES_BoyarPeralta_31_port_o_2_1;
  wire       [2:0]    sbox_AES_BoyarPeralta_31_port_o_2_2;
  wire       [2:0]    sbox_AES_BoyarPeralta_31_port_o_2_3;
  wire       [2:0]    sbox_AES_BoyarPeralta_31_port_o_2_4;
  wire       [2:0]    sbox_AES_BoyarPeralta_31_port_o_2_5;
  wire       [2:0]    sbox_AES_BoyarPeralta_31_port_o_2_6;
  wire       [2:0]    sbox_AES_BoyarPeralta_31_port_o_2_7;
  wire       [2:0]    sbox_AES_BoyarPeralta_31_port_o_3_0;
  wire       [2:0]    sbox_AES_BoyarPeralta_31_port_o_3_1;
  wire       [2:0]    sbox_AES_BoyarPeralta_31_port_o_3_2;
  wire       [2:0]    sbox_AES_BoyarPeralta_31_port_o_3_3;
  wire       [2:0]    sbox_AES_BoyarPeralta_31_port_o_3_4;
  wire       [2:0]    sbox_AES_BoyarPeralta_31_port_o_3_5;
  wire       [2:0]    sbox_AES_BoyarPeralta_31_port_o_3_6;
  wire       [2:0]    sbox_AES_BoyarPeralta_31_port_o_3_7;
  wire       [2:0]    shiftRows_port_state_out_0_0_0;
  wire       [2:0]    shiftRows_port_state_out_0_0_1;
  wire       [2:0]    shiftRows_port_state_out_0_0_2;
  wire       [2:0]    shiftRows_port_state_out_0_0_3;
  wire       [2:0]    shiftRows_port_state_out_0_0_4;
  wire       [2:0]    shiftRows_port_state_out_0_0_5;
  wire       [2:0]    shiftRows_port_state_out_0_0_6;
  wire       [2:0]    shiftRows_port_state_out_0_0_7;
  wire       [2:0]    shiftRows_port_state_out_0_1_0;
  wire       [2:0]    shiftRows_port_state_out_0_1_1;
  wire       [2:0]    shiftRows_port_state_out_0_1_2;
  wire       [2:0]    shiftRows_port_state_out_0_1_3;
  wire       [2:0]    shiftRows_port_state_out_0_1_4;
  wire       [2:0]    shiftRows_port_state_out_0_1_5;
  wire       [2:0]    shiftRows_port_state_out_0_1_6;
  wire       [2:0]    shiftRows_port_state_out_0_1_7;
  wire       [2:0]    shiftRows_port_state_out_0_2_0;
  wire       [2:0]    shiftRows_port_state_out_0_2_1;
  wire       [2:0]    shiftRows_port_state_out_0_2_2;
  wire       [2:0]    shiftRows_port_state_out_0_2_3;
  wire       [2:0]    shiftRows_port_state_out_0_2_4;
  wire       [2:0]    shiftRows_port_state_out_0_2_5;
  wire       [2:0]    shiftRows_port_state_out_0_2_6;
  wire       [2:0]    shiftRows_port_state_out_0_2_7;
  wire       [2:0]    shiftRows_port_state_out_0_3_0;
  wire       [2:0]    shiftRows_port_state_out_0_3_1;
  wire       [2:0]    shiftRows_port_state_out_0_3_2;
  wire       [2:0]    shiftRows_port_state_out_0_3_3;
  wire       [2:0]    shiftRows_port_state_out_0_3_4;
  wire       [2:0]    shiftRows_port_state_out_0_3_5;
  wire       [2:0]    shiftRows_port_state_out_0_3_6;
  wire       [2:0]    shiftRows_port_state_out_0_3_7;
  wire       [2:0]    shiftRows_port_state_out_1_0_0;
  wire       [2:0]    shiftRows_port_state_out_1_0_1;
  wire       [2:0]    shiftRows_port_state_out_1_0_2;
  wire       [2:0]    shiftRows_port_state_out_1_0_3;
  wire       [2:0]    shiftRows_port_state_out_1_0_4;
  wire       [2:0]    shiftRows_port_state_out_1_0_5;
  wire       [2:0]    shiftRows_port_state_out_1_0_6;
  wire       [2:0]    shiftRows_port_state_out_1_0_7;
  wire       [2:0]    shiftRows_port_state_out_1_1_0;
  wire       [2:0]    shiftRows_port_state_out_1_1_1;
  wire       [2:0]    shiftRows_port_state_out_1_1_2;
  wire       [2:0]    shiftRows_port_state_out_1_1_3;
  wire       [2:0]    shiftRows_port_state_out_1_1_4;
  wire       [2:0]    shiftRows_port_state_out_1_1_5;
  wire       [2:0]    shiftRows_port_state_out_1_1_6;
  wire       [2:0]    shiftRows_port_state_out_1_1_7;
  wire       [2:0]    shiftRows_port_state_out_1_2_0;
  wire       [2:0]    shiftRows_port_state_out_1_2_1;
  wire       [2:0]    shiftRows_port_state_out_1_2_2;
  wire       [2:0]    shiftRows_port_state_out_1_2_3;
  wire       [2:0]    shiftRows_port_state_out_1_2_4;
  wire       [2:0]    shiftRows_port_state_out_1_2_5;
  wire       [2:0]    shiftRows_port_state_out_1_2_6;
  wire       [2:0]    shiftRows_port_state_out_1_2_7;
  wire       [2:0]    shiftRows_port_state_out_1_3_0;
  wire       [2:0]    shiftRows_port_state_out_1_3_1;
  wire       [2:0]    shiftRows_port_state_out_1_3_2;
  wire       [2:0]    shiftRows_port_state_out_1_3_3;
  wire       [2:0]    shiftRows_port_state_out_1_3_4;
  wire       [2:0]    shiftRows_port_state_out_1_3_5;
  wire       [2:0]    shiftRows_port_state_out_1_3_6;
  wire       [2:0]    shiftRows_port_state_out_1_3_7;
  wire       [2:0]    shiftRows_port_state_out_2_0_0;
  wire       [2:0]    shiftRows_port_state_out_2_0_1;
  wire       [2:0]    shiftRows_port_state_out_2_0_2;
  wire       [2:0]    shiftRows_port_state_out_2_0_3;
  wire       [2:0]    shiftRows_port_state_out_2_0_4;
  wire       [2:0]    shiftRows_port_state_out_2_0_5;
  wire       [2:0]    shiftRows_port_state_out_2_0_6;
  wire       [2:0]    shiftRows_port_state_out_2_0_7;
  wire       [2:0]    shiftRows_port_state_out_2_1_0;
  wire       [2:0]    shiftRows_port_state_out_2_1_1;
  wire       [2:0]    shiftRows_port_state_out_2_1_2;
  wire       [2:0]    shiftRows_port_state_out_2_1_3;
  wire       [2:0]    shiftRows_port_state_out_2_1_4;
  wire       [2:0]    shiftRows_port_state_out_2_1_5;
  wire       [2:0]    shiftRows_port_state_out_2_1_6;
  wire       [2:0]    shiftRows_port_state_out_2_1_7;
  wire       [2:0]    shiftRows_port_state_out_2_2_0;
  wire       [2:0]    shiftRows_port_state_out_2_2_1;
  wire       [2:0]    shiftRows_port_state_out_2_2_2;
  wire       [2:0]    shiftRows_port_state_out_2_2_3;
  wire       [2:0]    shiftRows_port_state_out_2_2_4;
  wire       [2:0]    shiftRows_port_state_out_2_2_5;
  wire       [2:0]    shiftRows_port_state_out_2_2_6;
  wire       [2:0]    shiftRows_port_state_out_2_2_7;
  wire       [2:0]    shiftRows_port_state_out_2_3_0;
  wire       [2:0]    shiftRows_port_state_out_2_3_1;
  wire       [2:0]    shiftRows_port_state_out_2_3_2;
  wire       [2:0]    shiftRows_port_state_out_2_3_3;
  wire       [2:0]    shiftRows_port_state_out_2_3_4;
  wire       [2:0]    shiftRows_port_state_out_2_3_5;
  wire       [2:0]    shiftRows_port_state_out_2_3_6;
  wire       [2:0]    shiftRows_port_state_out_2_3_7;
  wire       [2:0]    shiftRows_port_state_out_3_0_0;
  wire       [2:0]    shiftRows_port_state_out_3_0_1;
  wire       [2:0]    shiftRows_port_state_out_3_0_2;
  wire       [2:0]    shiftRows_port_state_out_3_0_3;
  wire       [2:0]    shiftRows_port_state_out_3_0_4;
  wire       [2:0]    shiftRows_port_state_out_3_0_5;
  wire       [2:0]    shiftRows_port_state_out_3_0_6;
  wire       [2:0]    shiftRows_port_state_out_3_0_7;
  wire       [2:0]    shiftRows_port_state_out_3_1_0;
  wire       [2:0]    shiftRows_port_state_out_3_1_1;
  wire       [2:0]    shiftRows_port_state_out_3_1_2;
  wire       [2:0]    shiftRows_port_state_out_3_1_3;
  wire       [2:0]    shiftRows_port_state_out_3_1_4;
  wire       [2:0]    shiftRows_port_state_out_3_1_5;
  wire       [2:0]    shiftRows_port_state_out_3_1_6;
  wire       [2:0]    shiftRows_port_state_out_3_1_7;
  wire       [2:0]    shiftRows_port_state_out_3_2_0;
  wire       [2:0]    shiftRows_port_state_out_3_2_1;
  wire       [2:0]    shiftRows_port_state_out_3_2_2;
  wire       [2:0]    shiftRows_port_state_out_3_2_3;
  wire       [2:0]    shiftRows_port_state_out_3_2_4;
  wire       [2:0]    shiftRows_port_state_out_3_2_5;
  wire       [2:0]    shiftRows_port_state_out_3_2_6;
  wire       [2:0]    shiftRows_port_state_out_3_2_7;
  wire       [2:0]    shiftRows_port_state_out_3_3_0;
  wire       [2:0]    shiftRows_port_state_out_3_3_1;
  wire       [2:0]    shiftRows_port_state_out_3_3_2;
  wire       [2:0]    shiftRows_port_state_out_3_3_3;
  wire       [2:0]    shiftRows_port_state_out_3_3_4;
  wire       [2:0]    shiftRows_port_state_out_3_3_5;
  wire       [2:0]    shiftRows_port_state_out_3_3_6;
  wire       [2:0]    shiftRows_port_state_out_3_3_7;
  wire       [2:0]    shiftRows_port_state_out_4_0_0;
  wire       [2:0]    shiftRows_port_state_out_4_0_1;
  wire       [2:0]    shiftRows_port_state_out_4_0_2;
  wire       [2:0]    shiftRows_port_state_out_4_0_3;
  wire       [2:0]    shiftRows_port_state_out_4_0_4;
  wire       [2:0]    shiftRows_port_state_out_4_0_5;
  wire       [2:0]    shiftRows_port_state_out_4_0_6;
  wire       [2:0]    shiftRows_port_state_out_4_0_7;
  wire       [2:0]    shiftRows_port_state_out_4_1_0;
  wire       [2:0]    shiftRows_port_state_out_4_1_1;
  wire       [2:0]    shiftRows_port_state_out_4_1_2;
  wire       [2:0]    shiftRows_port_state_out_4_1_3;
  wire       [2:0]    shiftRows_port_state_out_4_1_4;
  wire       [2:0]    shiftRows_port_state_out_4_1_5;
  wire       [2:0]    shiftRows_port_state_out_4_1_6;
  wire       [2:0]    shiftRows_port_state_out_4_1_7;
  wire       [2:0]    shiftRows_port_state_out_4_2_0;
  wire       [2:0]    shiftRows_port_state_out_4_2_1;
  wire       [2:0]    shiftRows_port_state_out_4_2_2;
  wire       [2:0]    shiftRows_port_state_out_4_2_3;
  wire       [2:0]    shiftRows_port_state_out_4_2_4;
  wire       [2:0]    shiftRows_port_state_out_4_2_5;
  wire       [2:0]    shiftRows_port_state_out_4_2_6;
  wire       [2:0]    shiftRows_port_state_out_4_2_7;
  wire       [2:0]    shiftRows_port_state_out_4_3_0;
  wire       [2:0]    shiftRows_port_state_out_4_3_1;
  wire       [2:0]    shiftRows_port_state_out_4_3_2;
  wire       [2:0]    shiftRows_port_state_out_4_3_3;
  wire       [2:0]    shiftRows_port_state_out_4_3_4;
  wire       [2:0]    shiftRows_port_state_out_4_3_5;
  wire       [2:0]    shiftRows_port_state_out_4_3_6;
  wire       [2:0]    shiftRows_port_state_out_4_3_7;
  wire       [2:0]    shiftRows_port_state_out_5_0_0;
  wire       [2:0]    shiftRows_port_state_out_5_0_1;
  wire       [2:0]    shiftRows_port_state_out_5_0_2;
  wire       [2:0]    shiftRows_port_state_out_5_0_3;
  wire       [2:0]    shiftRows_port_state_out_5_0_4;
  wire       [2:0]    shiftRows_port_state_out_5_0_5;
  wire       [2:0]    shiftRows_port_state_out_5_0_6;
  wire       [2:0]    shiftRows_port_state_out_5_0_7;
  wire       [2:0]    shiftRows_port_state_out_5_1_0;
  wire       [2:0]    shiftRows_port_state_out_5_1_1;
  wire       [2:0]    shiftRows_port_state_out_5_1_2;
  wire       [2:0]    shiftRows_port_state_out_5_1_3;
  wire       [2:0]    shiftRows_port_state_out_5_1_4;
  wire       [2:0]    shiftRows_port_state_out_5_1_5;
  wire       [2:0]    shiftRows_port_state_out_5_1_6;
  wire       [2:0]    shiftRows_port_state_out_5_1_7;
  wire       [2:0]    shiftRows_port_state_out_5_2_0;
  wire       [2:0]    shiftRows_port_state_out_5_2_1;
  wire       [2:0]    shiftRows_port_state_out_5_2_2;
  wire       [2:0]    shiftRows_port_state_out_5_2_3;
  wire       [2:0]    shiftRows_port_state_out_5_2_4;
  wire       [2:0]    shiftRows_port_state_out_5_2_5;
  wire       [2:0]    shiftRows_port_state_out_5_2_6;
  wire       [2:0]    shiftRows_port_state_out_5_2_7;
  wire       [2:0]    shiftRows_port_state_out_5_3_0;
  wire       [2:0]    shiftRows_port_state_out_5_3_1;
  wire       [2:0]    shiftRows_port_state_out_5_3_2;
  wire       [2:0]    shiftRows_port_state_out_5_3_3;
  wire       [2:0]    shiftRows_port_state_out_5_3_4;
  wire       [2:0]    shiftRows_port_state_out_5_3_5;
  wire       [2:0]    shiftRows_port_state_out_5_3_6;
  wire       [2:0]    shiftRows_port_state_out_5_3_7;
  wire       [2:0]    shiftRows_port_state_out_6_0_0;
  wire       [2:0]    shiftRows_port_state_out_6_0_1;
  wire       [2:0]    shiftRows_port_state_out_6_0_2;
  wire       [2:0]    shiftRows_port_state_out_6_0_3;
  wire       [2:0]    shiftRows_port_state_out_6_0_4;
  wire       [2:0]    shiftRows_port_state_out_6_0_5;
  wire       [2:0]    shiftRows_port_state_out_6_0_6;
  wire       [2:0]    shiftRows_port_state_out_6_0_7;
  wire       [2:0]    shiftRows_port_state_out_6_1_0;
  wire       [2:0]    shiftRows_port_state_out_6_1_1;
  wire       [2:0]    shiftRows_port_state_out_6_1_2;
  wire       [2:0]    shiftRows_port_state_out_6_1_3;
  wire       [2:0]    shiftRows_port_state_out_6_1_4;
  wire       [2:0]    shiftRows_port_state_out_6_1_5;
  wire       [2:0]    shiftRows_port_state_out_6_1_6;
  wire       [2:0]    shiftRows_port_state_out_6_1_7;
  wire       [2:0]    shiftRows_port_state_out_6_2_0;
  wire       [2:0]    shiftRows_port_state_out_6_2_1;
  wire       [2:0]    shiftRows_port_state_out_6_2_2;
  wire       [2:0]    shiftRows_port_state_out_6_2_3;
  wire       [2:0]    shiftRows_port_state_out_6_2_4;
  wire       [2:0]    shiftRows_port_state_out_6_2_5;
  wire       [2:0]    shiftRows_port_state_out_6_2_6;
  wire       [2:0]    shiftRows_port_state_out_6_2_7;
  wire       [2:0]    shiftRows_port_state_out_6_3_0;
  wire       [2:0]    shiftRows_port_state_out_6_3_1;
  wire       [2:0]    shiftRows_port_state_out_6_3_2;
  wire       [2:0]    shiftRows_port_state_out_6_3_3;
  wire       [2:0]    shiftRows_port_state_out_6_3_4;
  wire       [2:0]    shiftRows_port_state_out_6_3_5;
  wire       [2:0]    shiftRows_port_state_out_6_3_6;
  wire       [2:0]    shiftRows_port_state_out_6_3_7;
  wire       [2:0]    shiftRows_port_state_out_7_0_0;
  wire       [2:0]    shiftRows_port_state_out_7_0_1;
  wire       [2:0]    shiftRows_port_state_out_7_0_2;
  wire       [2:0]    shiftRows_port_state_out_7_0_3;
  wire       [2:0]    shiftRows_port_state_out_7_0_4;
  wire       [2:0]    shiftRows_port_state_out_7_0_5;
  wire       [2:0]    shiftRows_port_state_out_7_0_6;
  wire       [2:0]    shiftRows_port_state_out_7_0_7;
  wire       [2:0]    shiftRows_port_state_out_7_1_0;
  wire       [2:0]    shiftRows_port_state_out_7_1_1;
  wire       [2:0]    shiftRows_port_state_out_7_1_2;
  wire       [2:0]    shiftRows_port_state_out_7_1_3;
  wire       [2:0]    shiftRows_port_state_out_7_1_4;
  wire       [2:0]    shiftRows_port_state_out_7_1_5;
  wire       [2:0]    shiftRows_port_state_out_7_1_6;
  wire       [2:0]    shiftRows_port_state_out_7_1_7;
  wire       [2:0]    shiftRows_port_state_out_7_2_0;
  wire       [2:0]    shiftRows_port_state_out_7_2_1;
  wire       [2:0]    shiftRows_port_state_out_7_2_2;
  wire       [2:0]    shiftRows_port_state_out_7_2_3;
  wire       [2:0]    shiftRows_port_state_out_7_2_4;
  wire       [2:0]    shiftRows_port_state_out_7_2_5;
  wire       [2:0]    shiftRows_port_state_out_7_2_6;
  wire       [2:0]    shiftRows_port_state_out_7_2_7;
  wire       [2:0]    shiftRows_port_state_out_7_3_0;
  wire       [2:0]    shiftRows_port_state_out_7_3_1;
  wire       [2:0]    shiftRows_port_state_out_7_3_2;
  wire       [2:0]    shiftRows_port_state_out_7_3_3;
  wire       [2:0]    shiftRows_port_state_out_7_3_4;
  wire       [2:0]    shiftRows_port_state_out_7_3_5;
  wire       [2:0]    shiftRows_port_state_out_7_3_6;
  wire       [2:0]    shiftRows_port_state_out_7_3_7;
  wire       [2:0]    shiftRows_port_state_out_8_0_0;
  wire       [2:0]    shiftRows_port_state_out_8_0_1;
  wire       [2:0]    shiftRows_port_state_out_8_0_2;
  wire       [2:0]    shiftRows_port_state_out_8_0_3;
  wire       [2:0]    shiftRows_port_state_out_8_0_4;
  wire       [2:0]    shiftRows_port_state_out_8_0_5;
  wire       [2:0]    shiftRows_port_state_out_8_0_6;
  wire       [2:0]    shiftRows_port_state_out_8_0_7;
  wire       [2:0]    shiftRows_port_state_out_8_1_0;
  wire       [2:0]    shiftRows_port_state_out_8_1_1;
  wire       [2:0]    shiftRows_port_state_out_8_1_2;
  wire       [2:0]    shiftRows_port_state_out_8_1_3;
  wire       [2:0]    shiftRows_port_state_out_8_1_4;
  wire       [2:0]    shiftRows_port_state_out_8_1_5;
  wire       [2:0]    shiftRows_port_state_out_8_1_6;
  wire       [2:0]    shiftRows_port_state_out_8_1_7;
  wire       [2:0]    shiftRows_port_state_out_8_2_0;
  wire       [2:0]    shiftRows_port_state_out_8_2_1;
  wire       [2:0]    shiftRows_port_state_out_8_2_2;
  wire       [2:0]    shiftRows_port_state_out_8_2_3;
  wire       [2:0]    shiftRows_port_state_out_8_2_4;
  wire       [2:0]    shiftRows_port_state_out_8_2_5;
  wire       [2:0]    shiftRows_port_state_out_8_2_6;
  wire       [2:0]    shiftRows_port_state_out_8_2_7;
  wire       [2:0]    shiftRows_port_state_out_8_3_0;
  wire       [2:0]    shiftRows_port_state_out_8_3_1;
  wire       [2:0]    shiftRows_port_state_out_8_3_2;
  wire       [2:0]    shiftRows_port_state_out_8_3_3;
  wire       [2:0]    shiftRows_port_state_out_8_3_4;
  wire       [2:0]    shiftRows_port_state_out_8_3_5;
  wire       [2:0]    shiftRows_port_state_out_8_3_6;
  wire       [2:0]    shiftRows_port_state_out_8_3_7;
  wire       [2:0]    shiftRows_port_state_out_9_0_0;
  wire       [2:0]    shiftRows_port_state_out_9_0_1;
  wire       [2:0]    shiftRows_port_state_out_9_0_2;
  wire       [2:0]    shiftRows_port_state_out_9_0_3;
  wire       [2:0]    shiftRows_port_state_out_9_0_4;
  wire       [2:0]    shiftRows_port_state_out_9_0_5;
  wire       [2:0]    shiftRows_port_state_out_9_0_6;
  wire       [2:0]    shiftRows_port_state_out_9_0_7;
  wire       [2:0]    shiftRows_port_state_out_9_1_0;
  wire       [2:0]    shiftRows_port_state_out_9_1_1;
  wire       [2:0]    shiftRows_port_state_out_9_1_2;
  wire       [2:0]    shiftRows_port_state_out_9_1_3;
  wire       [2:0]    shiftRows_port_state_out_9_1_4;
  wire       [2:0]    shiftRows_port_state_out_9_1_5;
  wire       [2:0]    shiftRows_port_state_out_9_1_6;
  wire       [2:0]    shiftRows_port_state_out_9_1_7;
  wire       [2:0]    shiftRows_port_state_out_9_2_0;
  wire       [2:0]    shiftRows_port_state_out_9_2_1;
  wire       [2:0]    shiftRows_port_state_out_9_2_2;
  wire       [2:0]    shiftRows_port_state_out_9_2_3;
  wire       [2:0]    shiftRows_port_state_out_9_2_4;
  wire       [2:0]    shiftRows_port_state_out_9_2_5;
  wire       [2:0]    shiftRows_port_state_out_9_2_6;
  wire       [2:0]    shiftRows_port_state_out_9_2_7;
  wire       [2:0]    shiftRows_port_state_out_9_3_0;
  wire       [2:0]    shiftRows_port_state_out_9_3_1;
  wire       [2:0]    shiftRows_port_state_out_9_3_2;
  wire       [2:0]    shiftRows_port_state_out_9_3_3;
  wire       [2:0]    shiftRows_port_state_out_9_3_4;
  wire       [2:0]    shiftRows_port_state_out_9_3_5;
  wire       [2:0]    shiftRows_port_state_out_9_3_6;
  wire       [2:0]    shiftRows_port_state_out_9_3_7;
  wire       [2:0]    shiftRows_port_state_out_10_0_0;
  wire       [2:0]    shiftRows_port_state_out_10_0_1;
  wire       [2:0]    shiftRows_port_state_out_10_0_2;
  wire       [2:0]    shiftRows_port_state_out_10_0_3;
  wire       [2:0]    shiftRows_port_state_out_10_0_4;
  wire       [2:0]    shiftRows_port_state_out_10_0_5;
  wire       [2:0]    shiftRows_port_state_out_10_0_6;
  wire       [2:0]    shiftRows_port_state_out_10_0_7;
  wire       [2:0]    shiftRows_port_state_out_10_1_0;
  wire       [2:0]    shiftRows_port_state_out_10_1_1;
  wire       [2:0]    shiftRows_port_state_out_10_1_2;
  wire       [2:0]    shiftRows_port_state_out_10_1_3;
  wire       [2:0]    shiftRows_port_state_out_10_1_4;
  wire       [2:0]    shiftRows_port_state_out_10_1_5;
  wire       [2:0]    shiftRows_port_state_out_10_1_6;
  wire       [2:0]    shiftRows_port_state_out_10_1_7;
  wire       [2:0]    shiftRows_port_state_out_10_2_0;
  wire       [2:0]    shiftRows_port_state_out_10_2_1;
  wire       [2:0]    shiftRows_port_state_out_10_2_2;
  wire       [2:0]    shiftRows_port_state_out_10_2_3;
  wire       [2:0]    shiftRows_port_state_out_10_2_4;
  wire       [2:0]    shiftRows_port_state_out_10_2_5;
  wire       [2:0]    shiftRows_port_state_out_10_2_6;
  wire       [2:0]    shiftRows_port_state_out_10_2_7;
  wire       [2:0]    shiftRows_port_state_out_10_3_0;
  wire       [2:0]    shiftRows_port_state_out_10_3_1;
  wire       [2:0]    shiftRows_port_state_out_10_3_2;
  wire       [2:0]    shiftRows_port_state_out_10_3_3;
  wire       [2:0]    shiftRows_port_state_out_10_3_4;
  wire       [2:0]    shiftRows_port_state_out_10_3_5;
  wire       [2:0]    shiftRows_port_state_out_10_3_6;
  wire       [2:0]    shiftRows_port_state_out_10_3_7;
  wire       [2:0]    shiftRows_port_state_out_11_0_0;
  wire       [2:0]    shiftRows_port_state_out_11_0_1;
  wire       [2:0]    shiftRows_port_state_out_11_0_2;
  wire       [2:0]    shiftRows_port_state_out_11_0_3;
  wire       [2:0]    shiftRows_port_state_out_11_0_4;
  wire       [2:0]    shiftRows_port_state_out_11_0_5;
  wire       [2:0]    shiftRows_port_state_out_11_0_6;
  wire       [2:0]    shiftRows_port_state_out_11_0_7;
  wire       [2:0]    shiftRows_port_state_out_11_1_0;
  wire       [2:0]    shiftRows_port_state_out_11_1_1;
  wire       [2:0]    shiftRows_port_state_out_11_1_2;
  wire       [2:0]    shiftRows_port_state_out_11_1_3;
  wire       [2:0]    shiftRows_port_state_out_11_1_4;
  wire       [2:0]    shiftRows_port_state_out_11_1_5;
  wire       [2:0]    shiftRows_port_state_out_11_1_6;
  wire       [2:0]    shiftRows_port_state_out_11_1_7;
  wire       [2:0]    shiftRows_port_state_out_11_2_0;
  wire       [2:0]    shiftRows_port_state_out_11_2_1;
  wire       [2:0]    shiftRows_port_state_out_11_2_2;
  wire       [2:0]    shiftRows_port_state_out_11_2_3;
  wire       [2:0]    shiftRows_port_state_out_11_2_4;
  wire       [2:0]    shiftRows_port_state_out_11_2_5;
  wire       [2:0]    shiftRows_port_state_out_11_2_6;
  wire       [2:0]    shiftRows_port_state_out_11_2_7;
  wire       [2:0]    shiftRows_port_state_out_11_3_0;
  wire       [2:0]    shiftRows_port_state_out_11_3_1;
  wire       [2:0]    shiftRows_port_state_out_11_3_2;
  wire       [2:0]    shiftRows_port_state_out_11_3_3;
  wire       [2:0]    shiftRows_port_state_out_11_3_4;
  wire       [2:0]    shiftRows_port_state_out_11_3_5;
  wire       [2:0]    shiftRows_port_state_out_11_3_6;
  wire       [2:0]    shiftRows_port_state_out_11_3_7;
  wire       [2:0]    shiftRows_port_state_out_12_0_0;
  wire       [2:0]    shiftRows_port_state_out_12_0_1;
  wire       [2:0]    shiftRows_port_state_out_12_0_2;
  wire       [2:0]    shiftRows_port_state_out_12_0_3;
  wire       [2:0]    shiftRows_port_state_out_12_0_4;
  wire       [2:0]    shiftRows_port_state_out_12_0_5;
  wire       [2:0]    shiftRows_port_state_out_12_0_6;
  wire       [2:0]    shiftRows_port_state_out_12_0_7;
  wire       [2:0]    shiftRows_port_state_out_12_1_0;
  wire       [2:0]    shiftRows_port_state_out_12_1_1;
  wire       [2:0]    shiftRows_port_state_out_12_1_2;
  wire       [2:0]    shiftRows_port_state_out_12_1_3;
  wire       [2:0]    shiftRows_port_state_out_12_1_4;
  wire       [2:0]    shiftRows_port_state_out_12_1_5;
  wire       [2:0]    shiftRows_port_state_out_12_1_6;
  wire       [2:0]    shiftRows_port_state_out_12_1_7;
  wire       [2:0]    shiftRows_port_state_out_12_2_0;
  wire       [2:0]    shiftRows_port_state_out_12_2_1;
  wire       [2:0]    shiftRows_port_state_out_12_2_2;
  wire       [2:0]    shiftRows_port_state_out_12_2_3;
  wire       [2:0]    shiftRows_port_state_out_12_2_4;
  wire       [2:0]    shiftRows_port_state_out_12_2_5;
  wire       [2:0]    shiftRows_port_state_out_12_2_6;
  wire       [2:0]    shiftRows_port_state_out_12_2_7;
  wire       [2:0]    shiftRows_port_state_out_12_3_0;
  wire       [2:0]    shiftRows_port_state_out_12_3_1;
  wire       [2:0]    shiftRows_port_state_out_12_3_2;
  wire       [2:0]    shiftRows_port_state_out_12_3_3;
  wire       [2:0]    shiftRows_port_state_out_12_3_4;
  wire       [2:0]    shiftRows_port_state_out_12_3_5;
  wire       [2:0]    shiftRows_port_state_out_12_3_6;
  wire       [2:0]    shiftRows_port_state_out_12_3_7;
  wire       [2:0]    shiftRows_port_state_out_13_0_0;
  wire       [2:0]    shiftRows_port_state_out_13_0_1;
  wire       [2:0]    shiftRows_port_state_out_13_0_2;
  wire       [2:0]    shiftRows_port_state_out_13_0_3;
  wire       [2:0]    shiftRows_port_state_out_13_0_4;
  wire       [2:0]    shiftRows_port_state_out_13_0_5;
  wire       [2:0]    shiftRows_port_state_out_13_0_6;
  wire       [2:0]    shiftRows_port_state_out_13_0_7;
  wire       [2:0]    shiftRows_port_state_out_13_1_0;
  wire       [2:0]    shiftRows_port_state_out_13_1_1;
  wire       [2:0]    shiftRows_port_state_out_13_1_2;
  wire       [2:0]    shiftRows_port_state_out_13_1_3;
  wire       [2:0]    shiftRows_port_state_out_13_1_4;
  wire       [2:0]    shiftRows_port_state_out_13_1_5;
  wire       [2:0]    shiftRows_port_state_out_13_1_6;
  wire       [2:0]    shiftRows_port_state_out_13_1_7;
  wire       [2:0]    shiftRows_port_state_out_13_2_0;
  wire       [2:0]    shiftRows_port_state_out_13_2_1;
  wire       [2:0]    shiftRows_port_state_out_13_2_2;
  wire       [2:0]    shiftRows_port_state_out_13_2_3;
  wire       [2:0]    shiftRows_port_state_out_13_2_4;
  wire       [2:0]    shiftRows_port_state_out_13_2_5;
  wire       [2:0]    shiftRows_port_state_out_13_2_6;
  wire       [2:0]    shiftRows_port_state_out_13_2_7;
  wire       [2:0]    shiftRows_port_state_out_13_3_0;
  wire       [2:0]    shiftRows_port_state_out_13_3_1;
  wire       [2:0]    shiftRows_port_state_out_13_3_2;
  wire       [2:0]    shiftRows_port_state_out_13_3_3;
  wire       [2:0]    shiftRows_port_state_out_13_3_4;
  wire       [2:0]    shiftRows_port_state_out_13_3_5;
  wire       [2:0]    shiftRows_port_state_out_13_3_6;
  wire       [2:0]    shiftRows_port_state_out_13_3_7;
  wire       [2:0]    shiftRows_port_state_out_14_0_0;
  wire       [2:0]    shiftRows_port_state_out_14_0_1;
  wire       [2:0]    shiftRows_port_state_out_14_0_2;
  wire       [2:0]    shiftRows_port_state_out_14_0_3;
  wire       [2:0]    shiftRows_port_state_out_14_0_4;
  wire       [2:0]    shiftRows_port_state_out_14_0_5;
  wire       [2:0]    shiftRows_port_state_out_14_0_6;
  wire       [2:0]    shiftRows_port_state_out_14_0_7;
  wire       [2:0]    shiftRows_port_state_out_14_1_0;
  wire       [2:0]    shiftRows_port_state_out_14_1_1;
  wire       [2:0]    shiftRows_port_state_out_14_1_2;
  wire       [2:0]    shiftRows_port_state_out_14_1_3;
  wire       [2:0]    shiftRows_port_state_out_14_1_4;
  wire       [2:0]    shiftRows_port_state_out_14_1_5;
  wire       [2:0]    shiftRows_port_state_out_14_1_6;
  wire       [2:0]    shiftRows_port_state_out_14_1_7;
  wire       [2:0]    shiftRows_port_state_out_14_2_0;
  wire       [2:0]    shiftRows_port_state_out_14_2_1;
  wire       [2:0]    shiftRows_port_state_out_14_2_2;
  wire       [2:0]    shiftRows_port_state_out_14_2_3;
  wire       [2:0]    shiftRows_port_state_out_14_2_4;
  wire       [2:0]    shiftRows_port_state_out_14_2_5;
  wire       [2:0]    shiftRows_port_state_out_14_2_6;
  wire       [2:0]    shiftRows_port_state_out_14_2_7;
  wire       [2:0]    shiftRows_port_state_out_14_3_0;
  wire       [2:0]    shiftRows_port_state_out_14_3_1;
  wire       [2:0]    shiftRows_port_state_out_14_3_2;
  wire       [2:0]    shiftRows_port_state_out_14_3_3;
  wire       [2:0]    shiftRows_port_state_out_14_3_4;
  wire       [2:0]    shiftRows_port_state_out_14_3_5;
  wire       [2:0]    shiftRows_port_state_out_14_3_6;
  wire       [2:0]    shiftRows_port_state_out_14_3_7;
  wire       [2:0]    shiftRows_port_state_out_15_0_0;
  wire       [2:0]    shiftRows_port_state_out_15_0_1;
  wire       [2:0]    shiftRows_port_state_out_15_0_2;
  wire       [2:0]    shiftRows_port_state_out_15_0_3;
  wire       [2:0]    shiftRows_port_state_out_15_0_4;
  wire       [2:0]    shiftRows_port_state_out_15_0_5;
  wire       [2:0]    shiftRows_port_state_out_15_0_6;
  wire       [2:0]    shiftRows_port_state_out_15_0_7;
  wire       [2:0]    shiftRows_port_state_out_15_1_0;
  wire       [2:0]    shiftRows_port_state_out_15_1_1;
  wire       [2:0]    shiftRows_port_state_out_15_1_2;
  wire       [2:0]    shiftRows_port_state_out_15_1_3;
  wire       [2:0]    shiftRows_port_state_out_15_1_4;
  wire       [2:0]    shiftRows_port_state_out_15_1_5;
  wire       [2:0]    shiftRows_port_state_out_15_1_6;
  wire       [2:0]    shiftRows_port_state_out_15_1_7;
  wire       [2:0]    shiftRows_port_state_out_15_2_0;
  wire       [2:0]    shiftRows_port_state_out_15_2_1;
  wire       [2:0]    shiftRows_port_state_out_15_2_2;
  wire       [2:0]    shiftRows_port_state_out_15_2_3;
  wire       [2:0]    shiftRows_port_state_out_15_2_4;
  wire       [2:0]    shiftRows_port_state_out_15_2_5;
  wire       [2:0]    shiftRows_port_state_out_15_2_6;
  wire       [2:0]    shiftRows_port_state_out_15_2_7;
  wire       [2:0]    shiftRows_port_state_out_15_3_0;
  wire       [2:0]    shiftRows_port_state_out_15_3_1;
  wire       [2:0]    shiftRows_port_state_out_15_3_2;
  wire       [2:0]    shiftRows_port_state_out_15_3_3;
  wire       [2:0]    shiftRows_port_state_out_15_3_4;
  wire       [2:0]    shiftRows_port_state_out_15_3_5;
  wire       [2:0]    shiftRows_port_state_out_15_3_6;
  wire       [2:0]    shiftRows_port_state_out_15_3_7;
  wire       [2:0]    mixColumns_port_state_out_0_0_0;
  wire       [2:0]    mixColumns_port_state_out_0_0_1;
  wire       [2:0]    mixColumns_port_state_out_0_0_2;
  wire       [2:0]    mixColumns_port_state_out_0_0_3;
  wire       [2:0]    mixColumns_port_state_out_0_0_4;
  wire       [2:0]    mixColumns_port_state_out_0_0_5;
  wire       [2:0]    mixColumns_port_state_out_0_0_6;
  wire       [2:0]    mixColumns_port_state_out_0_0_7;
  wire       [2:0]    mixColumns_port_state_out_0_1_0;
  wire       [2:0]    mixColumns_port_state_out_0_1_1;
  wire       [2:0]    mixColumns_port_state_out_0_1_2;
  wire       [2:0]    mixColumns_port_state_out_0_1_3;
  wire       [2:0]    mixColumns_port_state_out_0_1_4;
  wire       [2:0]    mixColumns_port_state_out_0_1_5;
  wire       [2:0]    mixColumns_port_state_out_0_1_6;
  wire       [2:0]    mixColumns_port_state_out_0_1_7;
  wire       [2:0]    mixColumns_port_state_out_0_2_0;
  wire       [2:0]    mixColumns_port_state_out_0_2_1;
  wire       [2:0]    mixColumns_port_state_out_0_2_2;
  wire       [2:0]    mixColumns_port_state_out_0_2_3;
  wire       [2:0]    mixColumns_port_state_out_0_2_4;
  wire       [2:0]    mixColumns_port_state_out_0_2_5;
  wire       [2:0]    mixColumns_port_state_out_0_2_6;
  wire       [2:0]    mixColumns_port_state_out_0_2_7;
  wire       [2:0]    mixColumns_port_state_out_0_3_0;
  wire       [2:0]    mixColumns_port_state_out_0_3_1;
  wire       [2:0]    mixColumns_port_state_out_0_3_2;
  wire       [2:0]    mixColumns_port_state_out_0_3_3;
  wire       [2:0]    mixColumns_port_state_out_0_3_4;
  wire       [2:0]    mixColumns_port_state_out_0_3_5;
  wire       [2:0]    mixColumns_port_state_out_0_3_6;
  wire       [2:0]    mixColumns_port_state_out_0_3_7;
  wire       [2:0]    mixColumns_port_state_out_1_0_0;
  wire       [2:0]    mixColumns_port_state_out_1_0_1;
  wire       [2:0]    mixColumns_port_state_out_1_0_2;
  wire       [2:0]    mixColumns_port_state_out_1_0_3;
  wire       [2:0]    mixColumns_port_state_out_1_0_4;
  wire       [2:0]    mixColumns_port_state_out_1_0_5;
  wire       [2:0]    mixColumns_port_state_out_1_0_6;
  wire       [2:0]    mixColumns_port_state_out_1_0_7;
  wire       [2:0]    mixColumns_port_state_out_1_1_0;
  wire       [2:0]    mixColumns_port_state_out_1_1_1;
  wire       [2:0]    mixColumns_port_state_out_1_1_2;
  wire       [2:0]    mixColumns_port_state_out_1_1_3;
  wire       [2:0]    mixColumns_port_state_out_1_1_4;
  wire       [2:0]    mixColumns_port_state_out_1_1_5;
  wire       [2:0]    mixColumns_port_state_out_1_1_6;
  wire       [2:0]    mixColumns_port_state_out_1_1_7;
  wire       [2:0]    mixColumns_port_state_out_1_2_0;
  wire       [2:0]    mixColumns_port_state_out_1_2_1;
  wire       [2:0]    mixColumns_port_state_out_1_2_2;
  wire       [2:0]    mixColumns_port_state_out_1_2_3;
  wire       [2:0]    mixColumns_port_state_out_1_2_4;
  wire       [2:0]    mixColumns_port_state_out_1_2_5;
  wire       [2:0]    mixColumns_port_state_out_1_2_6;
  wire       [2:0]    mixColumns_port_state_out_1_2_7;
  wire       [2:0]    mixColumns_port_state_out_1_3_0;
  wire       [2:0]    mixColumns_port_state_out_1_3_1;
  wire       [2:0]    mixColumns_port_state_out_1_3_2;
  wire       [2:0]    mixColumns_port_state_out_1_3_3;
  wire       [2:0]    mixColumns_port_state_out_1_3_4;
  wire       [2:0]    mixColumns_port_state_out_1_3_5;
  wire       [2:0]    mixColumns_port_state_out_1_3_6;
  wire       [2:0]    mixColumns_port_state_out_1_3_7;
  wire       [2:0]    mixColumns_port_state_out_2_0_0;
  wire       [2:0]    mixColumns_port_state_out_2_0_1;
  wire       [2:0]    mixColumns_port_state_out_2_0_2;
  wire       [2:0]    mixColumns_port_state_out_2_0_3;
  wire       [2:0]    mixColumns_port_state_out_2_0_4;
  wire       [2:0]    mixColumns_port_state_out_2_0_5;
  wire       [2:0]    mixColumns_port_state_out_2_0_6;
  wire       [2:0]    mixColumns_port_state_out_2_0_7;
  wire       [2:0]    mixColumns_port_state_out_2_1_0;
  wire       [2:0]    mixColumns_port_state_out_2_1_1;
  wire       [2:0]    mixColumns_port_state_out_2_1_2;
  wire       [2:0]    mixColumns_port_state_out_2_1_3;
  wire       [2:0]    mixColumns_port_state_out_2_1_4;
  wire       [2:0]    mixColumns_port_state_out_2_1_5;
  wire       [2:0]    mixColumns_port_state_out_2_1_6;
  wire       [2:0]    mixColumns_port_state_out_2_1_7;
  wire       [2:0]    mixColumns_port_state_out_2_2_0;
  wire       [2:0]    mixColumns_port_state_out_2_2_1;
  wire       [2:0]    mixColumns_port_state_out_2_2_2;
  wire       [2:0]    mixColumns_port_state_out_2_2_3;
  wire       [2:0]    mixColumns_port_state_out_2_2_4;
  wire       [2:0]    mixColumns_port_state_out_2_2_5;
  wire       [2:0]    mixColumns_port_state_out_2_2_6;
  wire       [2:0]    mixColumns_port_state_out_2_2_7;
  wire       [2:0]    mixColumns_port_state_out_2_3_0;
  wire       [2:0]    mixColumns_port_state_out_2_3_1;
  wire       [2:0]    mixColumns_port_state_out_2_3_2;
  wire       [2:0]    mixColumns_port_state_out_2_3_3;
  wire       [2:0]    mixColumns_port_state_out_2_3_4;
  wire       [2:0]    mixColumns_port_state_out_2_3_5;
  wire       [2:0]    mixColumns_port_state_out_2_3_6;
  wire       [2:0]    mixColumns_port_state_out_2_3_7;
  wire       [2:0]    mixColumns_port_state_out_3_0_0;
  wire       [2:0]    mixColumns_port_state_out_3_0_1;
  wire       [2:0]    mixColumns_port_state_out_3_0_2;
  wire       [2:0]    mixColumns_port_state_out_3_0_3;
  wire       [2:0]    mixColumns_port_state_out_3_0_4;
  wire       [2:0]    mixColumns_port_state_out_3_0_5;
  wire       [2:0]    mixColumns_port_state_out_3_0_6;
  wire       [2:0]    mixColumns_port_state_out_3_0_7;
  wire       [2:0]    mixColumns_port_state_out_3_1_0;
  wire       [2:0]    mixColumns_port_state_out_3_1_1;
  wire       [2:0]    mixColumns_port_state_out_3_1_2;
  wire       [2:0]    mixColumns_port_state_out_3_1_3;
  wire       [2:0]    mixColumns_port_state_out_3_1_4;
  wire       [2:0]    mixColumns_port_state_out_3_1_5;
  wire       [2:0]    mixColumns_port_state_out_3_1_6;
  wire       [2:0]    mixColumns_port_state_out_3_1_7;
  wire       [2:0]    mixColumns_port_state_out_3_2_0;
  wire       [2:0]    mixColumns_port_state_out_3_2_1;
  wire       [2:0]    mixColumns_port_state_out_3_2_2;
  wire       [2:0]    mixColumns_port_state_out_3_2_3;
  wire       [2:0]    mixColumns_port_state_out_3_2_4;
  wire       [2:0]    mixColumns_port_state_out_3_2_5;
  wire       [2:0]    mixColumns_port_state_out_3_2_6;
  wire       [2:0]    mixColumns_port_state_out_3_2_7;
  wire       [2:0]    mixColumns_port_state_out_3_3_0;
  wire       [2:0]    mixColumns_port_state_out_3_3_1;
  wire       [2:0]    mixColumns_port_state_out_3_3_2;
  wire       [2:0]    mixColumns_port_state_out_3_3_3;
  wire       [2:0]    mixColumns_port_state_out_3_3_4;
  wire       [2:0]    mixColumns_port_state_out_3_3_5;
  wire       [2:0]    mixColumns_port_state_out_3_3_6;
  wire       [2:0]    mixColumns_port_state_out_3_3_7;
  wire       [2:0]    mixColumns_port_state_out_4_0_0;
  wire       [2:0]    mixColumns_port_state_out_4_0_1;
  wire       [2:0]    mixColumns_port_state_out_4_0_2;
  wire       [2:0]    mixColumns_port_state_out_4_0_3;
  wire       [2:0]    mixColumns_port_state_out_4_0_4;
  wire       [2:0]    mixColumns_port_state_out_4_0_5;
  wire       [2:0]    mixColumns_port_state_out_4_0_6;
  wire       [2:0]    mixColumns_port_state_out_4_0_7;
  wire       [2:0]    mixColumns_port_state_out_4_1_0;
  wire       [2:0]    mixColumns_port_state_out_4_1_1;
  wire       [2:0]    mixColumns_port_state_out_4_1_2;
  wire       [2:0]    mixColumns_port_state_out_4_1_3;
  wire       [2:0]    mixColumns_port_state_out_4_1_4;
  wire       [2:0]    mixColumns_port_state_out_4_1_5;
  wire       [2:0]    mixColumns_port_state_out_4_1_6;
  wire       [2:0]    mixColumns_port_state_out_4_1_7;
  wire       [2:0]    mixColumns_port_state_out_4_2_0;
  wire       [2:0]    mixColumns_port_state_out_4_2_1;
  wire       [2:0]    mixColumns_port_state_out_4_2_2;
  wire       [2:0]    mixColumns_port_state_out_4_2_3;
  wire       [2:0]    mixColumns_port_state_out_4_2_4;
  wire       [2:0]    mixColumns_port_state_out_4_2_5;
  wire       [2:0]    mixColumns_port_state_out_4_2_6;
  wire       [2:0]    mixColumns_port_state_out_4_2_7;
  wire       [2:0]    mixColumns_port_state_out_4_3_0;
  wire       [2:0]    mixColumns_port_state_out_4_3_1;
  wire       [2:0]    mixColumns_port_state_out_4_3_2;
  wire       [2:0]    mixColumns_port_state_out_4_3_3;
  wire       [2:0]    mixColumns_port_state_out_4_3_4;
  wire       [2:0]    mixColumns_port_state_out_4_3_5;
  wire       [2:0]    mixColumns_port_state_out_4_3_6;
  wire       [2:0]    mixColumns_port_state_out_4_3_7;
  wire       [2:0]    mixColumns_port_state_out_5_0_0;
  wire       [2:0]    mixColumns_port_state_out_5_0_1;
  wire       [2:0]    mixColumns_port_state_out_5_0_2;
  wire       [2:0]    mixColumns_port_state_out_5_0_3;
  wire       [2:0]    mixColumns_port_state_out_5_0_4;
  wire       [2:0]    mixColumns_port_state_out_5_0_5;
  wire       [2:0]    mixColumns_port_state_out_5_0_6;
  wire       [2:0]    mixColumns_port_state_out_5_0_7;
  wire       [2:0]    mixColumns_port_state_out_5_1_0;
  wire       [2:0]    mixColumns_port_state_out_5_1_1;
  wire       [2:0]    mixColumns_port_state_out_5_1_2;
  wire       [2:0]    mixColumns_port_state_out_5_1_3;
  wire       [2:0]    mixColumns_port_state_out_5_1_4;
  wire       [2:0]    mixColumns_port_state_out_5_1_5;
  wire       [2:0]    mixColumns_port_state_out_5_1_6;
  wire       [2:0]    mixColumns_port_state_out_5_1_7;
  wire       [2:0]    mixColumns_port_state_out_5_2_0;
  wire       [2:0]    mixColumns_port_state_out_5_2_1;
  wire       [2:0]    mixColumns_port_state_out_5_2_2;
  wire       [2:0]    mixColumns_port_state_out_5_2_3;
  wire       [2:0]    mixColumns_port_state_out_5_2_4;
  wire       [2:0]    mixColumns_port_state_out_5_2_5;
  wire       [2:0]    mixColumns_port_state_out_5_2_6;
  wire       [2:0]    mixColumns_port_state_out_5_2_7;
  wire       [2:0]    mixColumns_port_state_out_5_3_0;
  wire       [2:0]    mixColumns_port_state_out_5_3_1;
  wire       [2:0]    mixColumns_port_state_out_5_3_2;
  wire       [2:0]    mixColumns_port_state_out_5_3_3;
  wire       [2:0]    mixColumns_port_state_out_5_3_4;
  wire       [2:0]    mixColumns_port_state_out_5_3_5;
  wire       [2:0]    mixColumns_port_state_out_5_3_6;
  wire       [2:0]    mixColumns_port_state_out_5_3_7;
  wire       [2:0]    mixColumns_port_state_out_6_0_0;
  wire       [2:0]    mixColumns_port_state_out_6_0_1;
  wire       [2:0]    mixColumns_port_state_out_6_0_2;
  wire       [2:0]    mixColumns_port_state_out_6_0_3;
  wire       [2:0]    mixColumns_port_state_out_6_0_4;
  wire       [2:0]    mixColumns_port_state_out_6_0_5;
  wire       [2:0]    mixColumns_port_state_out_6_0_6;
  wire       [2:0]    mixColumns_port_state_out_6_0_7;
  wire       [2:0]    mixColumns_port_state_out_6_1_0;
  wire       [2:0]    mixColumns_port_state_out_6_1_1;
  wire       [2:0]    mixColumns_port_state_out_6_1_2;
  wire       [2:0]    mixColumns_port_state_out_6_1_3;
  wire       [2:0]    mixColumns_port_state_out_6_1_4;
  wire       [2:0]    mixColumns_port_state_out_6_1_5;
  wire       [2:0]    mixColumns_port_state_out_6_1_6;
  wire       [2:0]    mixColumns_port_state_out_6_1_7;
  wire       [2:0]    mixColumns_port_state_out_6_2_0;
  wire       [2:0]    mixColumns_port_state_out_6_2_1;
  wire       [2:0]    mixColumns_port_state_out_6_2_2;
  wire       [2:0]    mixColumns_port_state_out_6_2_3;
  wire       [2:0]    mixColumns_port_state_out_6_2_4;
  wire       [2:0]    mixColumns_port_state_out_6_2_5;
  wire       [2:0]    mixColumns_port_state_out_6_2_6;
  wire       [2:0]    mixColumns_port_state_out_6_2_7;
  wire       [2:0]    mixColumns_port_state_out_6_3_0;
  wire       [2:0]    mixColumns_port_state_out_6_3_1;
  wire       [2:0]    mixColumns_port_state_out_6_3_2;
  wire       [2:0]    mixColumns_port_state_out_6_3_3;
  wire       [2:0]    mixColumns_port_state_out_6_3_4;
  wire       [2:0]    mixColumns_port_state_out_6_3_5;
  wire       [2:0]    mixColumns_port_state_out_6_3_6;
  wire       [2:0]    mixColumns_port_state_out_6_3_7;
  wire       [2:0]    mixColumns_port_state_out_7_0_0;
  wire       [2:0]    mixColumns_port_state_out_7_0_1;
  wire       [2:0]    mixColumns_port_state_out_7_0_2;
  wire       [2:0]    mixColumns_port_state_out_7_0_3;
  wire       [2:0]    mixColumns_port_state_out_7_0_4;
  wire       [2:0]    mixColumns_port_state_out_7_0_5;
  wire       [2:0]    mixColumns_port_state_out_7_0_6;
  wire       [2:0]    mixColumns_port_state_out_7_0_7;
  wire       [2:0]    mixColumns_port_state_out_7_1_0;
  wire       [2:0]    mixColumns_port_state_out_7_1_1;
  wire       [2:0]    mixColumns_port_state_out_7_1_2;
  wire       [2:0]    mixColumns_port_state_out_7_1_3;
  wire       [2:0]    mixColumns_port_state_out_7_1_4;
  wire       [2:0]    mixColumns_port_state_out_7_1_5;
  wire       [2:0]    mixColumns_port_state_out_7_1_6;
  wire       [2:0]    mixColumns_port_state_out_7_1_7;
  wire       [2:0]    mixColumns_port_state_out_7_2_0;
  wire       [2:0]    mixColumns_port_state_out_7_2_1;
  wire       [2:0]    mixColumns_port_state_out_7_2_2;
  wire       [2:0]    mixColumns_port_state_out_7_2_3;
  wire       [2:0]    mixColumns_port_state_out_7_2_4;
  wire       [2:0]    mixColumns_port_state_out_7_2_5;
  wire       [2:0]    mixColumns_port_state_out_7_2_6;
  wire       [2:0]    mixColumns_port_state_out_7_2_7;
  wire       [2:0]    mixColumns_port_state_out_7_3_0;
  wire       [2:0]    mixColumns_port_state_out_7_3_1;
  wire       [2:0]    mixColumns_port_state_out_7_3_2;
  wire       [2:0]    mixColumns_port_state_out_7_3_3;
  wire       [2:0]    mixColumns_port_state_out_7_3_4;
  wire       [2:0]    mixColumns_port_state_out_7_3_5;
  wire       [2:0]    mixColumns_port_state_out_7_3_6;
  wire       [2:0]    mixColumns_port_state_out_7_3_7;
  wire       [2:0]    mixColumns_port_state_out_8_0_0;
  wire       [2:0]    mixColumns_port_state_out_8_0_1;
  wire       [2:0]    mixColumns_port_state_out_8_0_2;
  wire       [2:0]    mixColumns_port_state_out_8_0_3;
  wire       [2:0]    mixColumns_port_state_out_8_0_4;
  wire       [2:0]    mixColumns_port_state_out_8_0_5;
  wire       [2:0]    mixColumns_port_state_out_8_0_6;
  wire       [2:0]    mixColumns_port_state_out_8_0_7;
  wire       [2:0]    mixColumns_port_state_out_8_1_0;
  wire       [2:0]    mixColumns_port_state_out_8_1_1;
  wire       [2:0]    mixColumns_port_state_out_8_1_2;
  wire       [2:0]    mixColumns_port_state_out_8_1_3;
  wire       [2:0]    mixColumns_port_state_out_8_1_4;
  wire       [2:0]    mixColumns_port_state_out_8_1_5;
  wire       [2:0]    mixColumns_port_state_out_8_1_6;
  wire       [2:0]    mixColumns_port_state_out_8_1_7;
  wire       [2:0]    mixColumns_port_state_out_8_2_0;
  wire       [2:0]    mixColumns_port_state_out_8_2_1;
  wire       [2:0]    mixColumns_port_state_out_8_2_2;
  wire       [2:0]    mixColumns_port_state_out_8_2_3;
  wire       [2:0]    mixColumns_port_state_out_8_2_4;
  wire       [2:0]    mixColumns_port_state_out_8_2_5;
  wire       [2:0]    mixColumns_port_state_out_8_2_6;
  wire       [2:0]    mixColumns_port_state_out_8_2_7;
  wire       [2:0]    mixColumns_port_state_out_8_3_0;
  wire       [2:0]    mixColumns_port_state_out_8_3_1;
  wire       [2:0]    mixColumns_port_state_out_8_3_2;
  wire       [2:0]    mixColumns_port_state_out_8_3_3;
  wire       [2:0]    mixColumns_port_state_out_8_3_4;
  wire       [2:0]    mixColumns_port_state_out_8_3_5;
  wire       [2:0]    mixColumns_port_state_out_8_3_6;
  wire       [2:0]    mixColumns_port_state_out_8_3_7;
  wire       [2:0]    mixColumns_port_state_out_9_0_0;
  wire       [2:0]    mixColumns_port_state_out_9_0_1;
  wire       [2:0]    mixColumns_port_state_out_9_0_2;
  wire       [2:0]    mixColumns_port_state_out_9_0_3;
  wire       [2:0]    mixColumns_port_state_out_9_0_4;
  wire       [2:0]    mixColumns_port_state_out_9_0_5;
  wire       [2:0]    mixColumns_port_state_out_9_0_6;
  wire       [2:0]    mixColumns_port_state_out_9_0_7;
  wire       [2:0]    mixColumns_port_state_out_9_1_0;
  wire       [2:0]    mixColumns_port_state_out_9_1_1;
  wire       [2:0]    mixColumns_port_state_out_9_1_2;
  wire       [2:0]    mixColumns_port_state_out_9_1_3;
  wire       [2:0]    mixColumns_port_state_out_9_1_4;
  wire       [2:0]    mixColumns_port_state_out_9_1_5;
  wire       [2:0]    mixColumns_port_state_out_9_1_6;
  wire       [2:0]    mixColumns_port_state_out_9_1_7;
  wire       [2:0]    mixColumns_port_state_out_9_2_0;
  wire       [2:0]    mixColumns_port_state_out_9_2_1;
  wire       [2:0]    mixColumns_port_state_out_9_2_2;
  wire       [2:0]    mixColumns_port_state_out_9_2_3;
  wire       [2:0]    mixColumns_port_state_out_9_2_4;
  wire       [2:0]    mixColumns_port_state_out_9_2_5;
  wire       [2:0]    mixColumns_port_state_out_9_2_6;
  wire       [2:0]    mixColumns_port_state_out_9_2_7;
  wire       [2:0]    mixColumns_port_state_out_9_3_0;
  wire       [2:0]    mixColumns_port_state_out_9_3_1;
  wire       [2:0]    mixColumns_port_state_out_9_3_2;
  wire       [2:0]    mixColumns_port_state_out_9_3_3;
  wire       [2:0]    mixColumns_port_state_out_9_3_4;
  wire       [2:0]    mixColumns_port_state_out_9_3_5;
  wire       [2:0]    mixColumns_port_state_out_9_3_6;
  wire       [2:0]    mixColumns_port_state_out_9_3_7;
  wire       [2:0]    mixColumns_port_state_out_10_0_0;
  wire       [2:0]    mixColumns_port_state_out_10_0_1;
  wire       [2:0]    mixColumns_port_state_out_10_0_2;
  wire       [2:0]    mixColumns_port_state_out_10_0_3;
  wire       [2:0]    mixColumns_port_state_out_10_0_4;
  wire       [2:0]    mixColumns_port_state_out_10_0_5;
  wire       [2:0]    mixColumns_port_state_out_10_0_6;
  wire       [2:0]    mixColumns_port_state_out_10_0_7;
  wire       [2:0]    mixColumns_port_state_out_10_1_0;
  wire       [2:0]    mixColumns_port_state_out_10_1_1;
  wire       [2:0]    mixColumns_port_state_out_10_1_2;
  wire       [2:0]    mixColumns_port_state_out_10_1_3;
  wire       [2:0]    mixColumns_port_state_out_10_1_4;
  wire       [2:0]    mixColumns_port_state_out_10_1_5;
  wire       [2:0]    mixColumns_port_state_out_10_1_6;
  wire       [2:0]    mixColumns_port_state_out_10_1_7;
  wire       [2:0]    mixColumns_port_state_out_10_2_0;
  wire       [2:0]    mixColumns_port_state_out_10_2_1;
  wire       [2:0]    mixColumns_port_state_out_10_2_2;
  wire       [2:0]    mixColumns_port_state_out_10_2_3;
  wire       [2:0]    mixColumns_port_state_out_10_2_4;
  wire       [2:0]    mixColumns_port_state_out_10_2_5;
  wire       [2:0]    mixColumns_port_state_out_10_2_6;
  wire       [2:0]    mixColumns_port_state_out_10_2_7;
  wire       [2:0]    mixColumns_port_state_out_10_3_0;
  wire       [2:0]    mixColumns_port_state_out_10_3_1;
  wire       [2:0]    mixColumns_port_state_out_10_3_2;
  wire       [2:0]    mixColumns_port_state_out_10_3_3;
  wire       [2:0]    mixColumns_port_state_out_10_3_4;
  wire       [2:0]    mixColumns_port_state_out_10_3_5;
  wire       [2:0]    mixColumns_port_state_out_10_3_6;
  wire       [2:0]    mixColumns_port_state_out_10_3_7;
  wire       [2:0]    mixColumns_port_state_out_11_0_0;
  wire       [2:0]    mixColumns_port_state_out_11_0_1;
  wire       [2:0]    mixColumns_port_state_out_11_0_2;
  wire       [2:0]    mixColumns_port_state_out_11_0_3;
  wire       [2:0]    mixColumns_port_state_out_11_0_4;
  wire       [2:0]    mixColumns_port_state_out_11_0_5;
  wire       [2:0]    mixColumns_port_state_out_11_0_6;
  wire       [2:0]    mixColumns_port_state_out_11_0_7;
  wire       [2:0]    mixColumns_port_state_out_11_1_0;
  wire       [2:0]    mixColumns_port_state_out_11_1_1;
  wire       [2:0]    mixColumns_port_state_out_11_1_2;
  wire       [2:0]    mixColumns_port_state_out_11_1_3;
  wire       [2:0]    mixColumns_port_state_out_11_1_4;
  wire       [2:0]    mixColumns_port_state_out_11_1_5;
  wire       [2:0]    mixColumns_port_state_out_11_1_6;
  wire       [2:0]    mixColumns_port_state_out_11_1_7;
  wire       [2:0]    mixColumns_port_state_out_11_2_0;
  wire       [2:0]    mixColumns_port_state_out_11_2_1;
  wire       [2:0]    mixColumns_port_state_out_11_2_2;
  wire       [2:0]    mixColumns_port_state_out_11_2_3;
  wire       [2:0]    mixColumns_port_state_out_11_2_4;
  wire       [2:0]    mixColumns_port_state_out_11_2_5;
  wire       [2:0]    mixColumns_port_state_out_11_2_6;
  wire       [2:0]    mixColumns_port_state_out_11_2_7;
  wire       [2:0]    mixColumns_port_state_out_11_3_0;
  wire       [2:0]    mixColumns_port_state_out_11_3_1;
  wire       [2:0]    mixColumns_port_state_out_11_3_2;
  wire       [2:0]    mixColumns_port_state_out_11_3_3;
  wire       [2:0]    mixColumns_port_state_out_11_3_4;
  wire       [2:0]    mixColumns_port_state_out_11_3_5;
  wire       [2:0]    mixColumns_port_state_out_11_3_6;
  wire       [2:0]    mixColumns_port_state_out_11_3_7;
  wire       [2:0]    mixColumns_port_state_out_12_0_0;
  wire       [2:0]    mixColumns_port_state_out_12_0_1;
  wire       [2:0]    mixColumns_port_state_out_12_0_2;
  wire       [2:0]    mixColumns_port_state_out_12_0_3;
  wire       [2:0]    mixColumns_port_state_out_12_0_4;
  wire       [2:0]    mixColumns_port_state_out_12_0_5;
  wire       [2:0]    mixColumns_port_state_out_12_0_6;
  wire       [2:0]    mixColumns_port_state_out_12_0_7;
  wire       [2:0]    mixColumns_port_state_out_12_1_0;
  wire       [2:0]    mixColumns_port_state_out_12_1_1;
  wire       [2:0]    mixColumns_port_state_out_12_1_2;
  wire       [2:0]    mixColumns_port_state_out_12_1_3;
  wire       [2:0]    mixColumns_port_state_out_12_1_4;
  wire       [2:0]    mixColumns_port_state_out_12_1_5;
  wire       [2:0]    mixColumns_port_state_out_12_1_6;
  wire       [2:0]    mixColumns_port_state_out_12_1_7;
  wire       [2:0]    mixColumns_port_state_out_12_2_0;
  wire       [2:0]    mixColumns_port_state_out_12_2_1;
  wire       [2:0]    mixColumns_port_state_out_12_2_2;
  wire       [2:0]    mixColumns_port_state_out_12_2_3;
  wire       [2:0]    mixColumns_port_state_out_12_2_4;
  wire       [2:0]    mixColumns_port_state_out_12_2_5;
  wire       [2:0]    mixColumns_port_state_out_12_2_6;
  wire       [2:0]    mixColumns_port_state_out_12_2_7;
  wire       [2:0]    mixColumns_port_state_out_12_3_0;
  wire       [2:0]    mixColumns_port_state_out_12_3_1;
  wire       [2:0]    mixColumns_port_state_out_12_3_2;
  wire       [2:0]    mixColumns_port_state_out_12_3_3;
  wire       [2:0]    mixColumns_port_state_out_12_3_4;
  wire       [2:0]    mixColumns_port_state_out_12_3_5;
  wire       [2:0]    mixColumns_port_state_out_12_3_6;
  wire       [2:0]    mixColumns_port_state_out_12_3_7;
  wire       [2:0]    mixColumns_port_state_out_13_0_0;
  wire       [2:0]    mixColumns_port_state_out_13_0_1;
  wire       [2:0]    mixColumns_port_state_out_13_0_2;
  wire       [2:0]    mixColumns_port_state_out_13_0_3;
  wire       [2:0]    mixColumns_port_state_out_13_0_4;
  wire       [2:0]    mixColumns_port_state_out_13_0_5;
  wire       [2:0]    mixColumns_port_state_out_13_0_6;
  wire       [2:0]    mixColumns_port_state_out_13_0_7;
  wire       [2:0]    mixColumns_port_state_out_13_1_0;
  wire       [2:0]    mixColumns_port_state_out_13_1_1;
  wire       [2:0]    mixColumns_port_state_out_13_1_2;
  wire       [2:0]    mixColumns_port_state_out_13_1_3;
  wire       [2:0]    mixColumns_port_state_out_13_1_4;
  wire       [2:0]    mixColumns_port_state_out_13_1_5;
  wire       [2:0]    mixColumns_port_state_out_13_1_6;
  wire       [2:0]    mixColumns_port_state_out_13_1_7;
  wire       [2:0]    mixColumns_port_state_out_13_2_0;
  wire       [2:0]    mixColumns_port_state_out_13_2_1;
  wire       [2:0]    mixColumns_port_state_out_13_2_2;
  wire       [2:0]    mixColumns_port_state_out_13_2_3;
  wire       [2:0]    mixColumns_port_state_out_13_2_4;
  wire       [2:0]    mixColumns_port_state_out_13_2_5;
  wire       [2:0]    mixColumns_port_state_out_13_2_6;
  wire       [2:0]    mixColumns_port_state_out_13_2_7;
  wire       [2:0]    mixColumns_port_state_out_13_3_0;
  wire       [2:0]    mixColumns_port_state_out_13_3_1;
  wire       [2:0]    mixColumns_port_state_out_13_3_2;
  wire       [2:0]    mixColumns_port_state_out_13_3_3;
  wire       [2:0]    mixColumns_port_state_out_13_3_4;
  wire       [2:0]    mixColumns_port_state_out_13_3_5;
  wire       [2:0]    mixColumns_port_state_out_13_3_6;
  wire       [2:0]    mixColumns_port_state_out_13_3_7;
  wire       [2:0]    mixColumns_port_state_out_14_0_0;
  wire       [2:0]    mixColumns_port_state_out_14_0_1;
  wire       [2:0]    mixColumns_port_state_out_14_0_2;
  wire       [2:0]    mixColumns_port_state_out_14_0_3;
  wire       [2:0]    mixColumns_port_state_out_14_0_4;
  wire       [2:0]    mixColumns_port_state_out_14_0_5;
  wire       [2:0]    mixColumns_port_state_out_14_0_6;
  wire       [2:0]    mixColumns_port_state_out_14_0_7;
  wire       [2:0]    mixColumns_port_state_out_14_1_0;
  wire       [2:0]    mixColumns_port_state_out_14_1_1;
  wire       [2:0]    mixColumns_port_state_out_14_1_2;
  wire       [2:0]    mixColumns_port_state_out_14_1_3;
  wire       [2:0]    mixColumns_port_state_out_14_1_4;
  wire       [2:0]    mixColumns_port_state_out_14_1_5;
  wire       [2:0]    mixColumns_port_state_out_14_1_6;
  wire       [2:0]    mixColumns_port_state_out_14_1_7;
  wire       [2:0]    mixColumns_port_state_out_14_2_0;
  wire       [2:0]    mixColumns_port_state_out_14_2_1;
  wire       [2:0]    mixColumns_port_state_out_14_2_2;
  wire       [2:0]    mixColumns_port_state_out_14_2_3;
  wire       [2:0]    mixColumns_port_state_out_14_2_4;
  wire       [2:0]    mixColumns_port_state_out_14_2_5;
  wire       [2:0]    mixColumns_port_state_out_14_2_6;
  wire       [2:0]    mixColumns_port_state_out_14_2_7;
  wire       [2:0]    mixColumns_port_state_out_14_3_0;
  wire       [2:0]    mixColumns_port_state_out_14_3_1;
  wire       [2:0]    mixColumns_port_state_out_14_3_2;
  wire       [2:0]    mixColumns_port_state_out_14_3_3;
  wire       [2:0]    mixColumns_port_state_out_14_3_4;
  wire       [2:0]    mixColumns_port_state_out_14_3_5;
  wire       [2:0]    mixColumns_port_state_out_14_3_6;
  wire       [2:0]    mixColumns_port_state_out_14_3_7;
  wire       [2:0]    mixColumns_port_state_out_15_0_0;
  wire       [2:0]    mixColumns_port_state_out_15_0_1;
  wire       [2:0]    mixColumns_port_state_out_15_0_2;
  wire       [2:0]    mixColumns_port_state_out_15_0_3;
  wire       [2:0]    mixColumns_port_state_out_15_0_4;
  wire       [2:0]    mixColumns_port_state_out_15_0_5;
  wire       [2:0]    mixColumns_port_state_out_15_0_6;
  wire       [2:0]    mixColumns_port_state_out_15_0_7;
  wire       [2:0]    mixColumns_port_state_out_15_1_0;
  wire       [2:0]    mixColumns_port_state_out_15_1_1;
  wire       [2:0]    mixColumns_port_state_out_15_1_2;
  wire       [2:0]    mixColumns_port_state_out_15_1_3;
  wire       [2:0]    mixColumns_port_state_out_15_1_4;
  wire       [2:0]    mixColumns_port_state_out_15_1_5;
  wire       [2:0]    mixColumns_port_state_out_15_1_6;
  wire       [2:0]    mixColumns_port_state_out_15_1_7;
  wire       [2:0]    mixColumns_port_state_out_15_2_0;
  wire       [2:0]    mixColumns_port_state_out_15_2_1;
  wire       [2:0]    mixColumns_port_state_out_15_2_2;
  wire       [2:0]    mixColumns_port_state_out_15_2_3;
  wire       [2:0]    mixColumns_port_state_out_15_2_4;
  wire       [2:0]    mixColumns_port_state_out_15_2_5;
  wire       [2:0]    mixColumns_port_state_out_15_2_6;
  wire       [2:0]    mixColumns_port_state_out_15_2_7;
  wire       [2:0]    mixColumns_port_state_out_15_3_0;
  wire       [2:0]    mixColumns_port_state_out_15_3_1;
  wire       [2:0]    mixColumns_port_state_out_15_3_2;
  wire       [2:0]    mixColumns_port_state_out_15_3_3;
  wire       [2:0]    mixColumns_port_state_out_15_3_4;
  wire       [2:0]    mixColumns_port_state_out_15_3_5;
  wire       [2:0]    mixColumns_port_state_out_15_3_6;
  wire       [2:0]    mixColumns_port_state_out_15_3_7;
  wire                majority_4608_port_o;
  wire                majority_4609_port_o;
  wire                majority_4610_port_o;
  wire                majority_4611_port_o;
  wire                majority_4612_port_o;
  wire                majority_4613_port_o;
  wire                majority_4614_port_o;
  wire                majority_4615_port_o;
  wire                majority_4616_port_o;
  wire                majority_4617_port_o;
  wire                majority_4618_port_o;
  wire                majority_4619_port_o;
  wire                majority_4620_port_o;
  wire                majority_4621_port_o;
  wire                majority_4622_port_o;
  wire                majority_4623_port_o;
  wire                majority_4624_port_o;
  wire                majority_4625_port_o;
  wire                majority_4626_port_o;
  wire                majority_4627_port_o;
  wire                majority_4628_port_o;
  wire                majority_4629_port_o;
  wire                majority_4630_port_o;
  wire                majority_4631_port_o;
  wire                majority_4632_port_o;
  wire                majority_4633_port_o;
  wire                majority_4634_port_o;
  wire                majority_4635_port_o;
  wire                majority_4636_port_o;
  wire                majority_4637_port_o;
  wire                majority_4638_port_o;
  wire                majority_4639_port_o;
  wire                majority_4640_port_o;
  wire                majority_4641_port_o;
  wire                majority_4642_port_o;
  wire                majority_4643_port_o;
  wire                majority_4644_port_o;
  wire                majority_4645_port_o;
  wire                majority_4646_port_o;
  wire                majority_4647_port_o;
  wire                majority_4648_port_o;
  wire                majority_4649_port_o;
  wire                majority_4650_port_o;
  wire                majority_4651_port_o;
  wire                majority_4652_port_o;
  wire                majority_4653_port_o;
  wire                majority_4654_port_o;
  wire                majority_4655_port_o;
  wire                majority_4656_port_o;
  wire                majority_4657_port_o;
  wire                majority_4658_port_o;
  wire                majority_4659_port_o;
  wire                majority_4660_port_o;
  wire                majority_4661_port_o;
  wire                majority_4662_port_o;
  wire                majority_4663_port_o;
  wire                majority_4664_port_o;
  wire                majority_4665_port_o;
  wire                majority_4666_port_o;
  wire                majority_4667_port_o;
  wire                majority_4668_port_o;
  wire                majority_4669_port_o;
  wire                majority_4670_port_o;
  wire                majority_4671_port_o;
  wire                majority_4672_port_o;
  wire                majority_4673_port_o;
  wire                majority_4674_port_o;
  wire                majority_4675_port_o;
  wire                majority_4676_port_o;
  wire                majority_4677_port_o;
  wire                majority_4678_port_o;
  wire                majority_4679_port_o;
  wire                majority_4680_port_o;
  wire                majority_4681_port_o;
  wire                majority_4682_port_o;
  wire                majority_4683_port_o;
  wire                majority_4684_port_o;
  wire                majority_4685_port_o;
  wire                majority_4686_port_o;
  wire                majority_4687_port_o;
  wire                majority_4688_port_o;
  wire                majority_4689_port_o;
  wire                majority_4690_port_o;
  wire                majority_4691_port_o;
  wire                majority_4692_port_o;
  wire                majority_4693_port_o;
  wire                majority_4694_port_o;
  wire                majority_4695_port_o;
  wire                majority_4696_port_o;
  wire                majority_4697_port_o;
  wire                majority_4698_port_o;
  wire                majority_4699_port_o;
  wire                majority_4700_port_o;
  wire                majority_4701_port_o;
  wire                majority_4702_port_o;
  wire                majority_4703_port_o;
  wire                majority_4704_port_o;
  wire                majority_4705_port_o;
  wire                majority_4706_port_o;
  wire                majority_4707_port_o;
  wire                majority_4708_port_o;
  wire                majority_4709_port_o;
  wire                majority_4710_port_o;
  wire                majority_4711_port_o;
  wire                majority_4712_port_o;
  wire                majority_4713_port_o;
  wire                majority_4714_port_o;
  wire                majority_4715_port_o;
  wire                majority_4716_port_o;
  wire                majority_4717_port_o;
  wire                majority_4718_port_o;
  wire                majority_4719_port_o;
  wire                majority_4720_port_o;
  wire                majority_4721_port_o;
  wire                majority_4722_port_o;
  wire                majority_4723_port_o;
  wire                majority_4724_port_o;
  wire                majority_4725_port_o;
  wire                majority_4726_port_o;
  wire                majority_4727_port_o;
  wire                majority_4728_port_o;
  wire                majority_4729_port_o;
  wire                majority_4730_port_o;
  wire                majority_4731_port_o;
  wire                majority_4732_port_o;
  wire                majority_4733_port_o;
  wire                majority_4734_port_o;
  wire                majority_4735_port_o;
  wire                majority_4736_port_o;
  wire                majority_4737_port_o;
  wire                majority_4738_port_o;
  wire                majority_4739_port_o;
  wire                majority_4740_port_o;
  wire                majority_4741_port_o;
  wire                majority_4742_port_o;
  wire                majority_4743_port_o;
  wire                majority_4744_port_o;
  wire                majority_4745_port_o;
  wire                majority_4746_port_o;
  wire                majority_4747_port_o;
  wire                majority_4748_port_o;
  wire                majority_4749_port_o;
  wire                majority_4750_port_o;
  wire                majority_4751_port_o;
  wire                majority_4752_port_o;
  wire                majority_4753_port_o;
  wire                majority_4754_port_o;
  wire                majority_4755_port_o;
  wire                majority_4756_port_o;
  wire                majority_4757_port_o;
  wire                majority_4758_port_o;
  wire                majority_4759_port_o;
  wire                majority_4760_port_o;
  wire                majority_4761_port_o;
  wire                majority_4762_port_o;
  wire                majority_4763_port_o;
  wire                majority_4764_port_o;
  wire                majority_4765_port_o;
  wire                majority_4766_port_o;
  wire                majority_4767_port_o;
  wire                majority_4768_port_o;
  wire                majority_4769_port_o;
  wire                majority_4770_port_o;
  wire                majority_4771_port_o;
  wire                majority_4772_port_o;
  wire                majority_4773_port_o;
  wire                majority_4774_port_o;
  wire                majority_4775_port_o;
  wire                majority_4776_port_o;
  wire                majority_4777_port_o;
  wire                majority_4778_port_o;
  wire                majority_4779_port_o;
  wire                majority_4780_port_o;
  wire                majority_4781_port_o;
  wire                majority_4782_port_o;
  wire                majority_4783_port_o;
  wire                majority_4784_port_o;
  wire                majority_4785_port_o;
  wire                majority_4786_port_o;
  wire                majority_4787_port_o;
  wire                majority_4788_port_o;
  wire                majority_4789_port_o;
  wire                majority_4790_port_o;
  wire                majority_4791_port_o;
  wire                majority_4792_port_o;
  wire                majority_4793_port_o;
  wire                majority_4794_port_o;
  wire                majority_4795_port_o;
  wire                majority_4796_port_o;
  wire                majority_4797_port_o;
  wire                majority_4798_port_o;
  wire                majority_4799_port_o;
  wire                majority_4800_port_o;
  wire                majority_4801_port_o;
  wire                majority_4802_port_o;
  wire                majority_4803_port_o;
  wire                majority_4804_port_o;
  wire                majority_4805_port_o;
  wire                majority_4806_port_o;
  wire                majority_4807_port_o;
  wire                majority_4808_port_o;
  wire                majority_4809_port_o;
  wire                majority_4810_port_o;
  wire                majority_4811_port_o;
  wire                majority_4812_port_o;
  wire                majority_4813_port_o;
  wire                majority_4814_port_o;
  wire                majority_4815_port_o;
  wire                majority_4816_port_o;
  wire                majority_4817_port_o;
  wire                majority_4818_port_o;
  wire                majority_4819_port_o;
  wire                majority_4820_port_o;
  wire                majority_4821_port_o;
  wire                majority_4822_port_o;
  wire                majority_4823_port_o;
  wire                majority_4824_port_o;
  wire                majority_4825_port_o;
  wire                majority_4826_port_o;
  wire                majority_4827_port_o;
  wire                majority_4828_port_o;
  wire                majority_4829_port_o;
  wire                majority_4830_port_o;
  wire                majority_4831_port_o;
  wire                majority_4832_port_o;
  wire                majority_4833_port_o;
  wire                majority_4834_port_o;
  wire                majority_4835_port_o;
  wire                majority_4836_port_o;
  wire                majority_4837_port_o;
  wire                majority_4838_port_o;
  wire                majority_4839_port_o;
  wire                majority_4840_port_o;
  wire                majority_4841_port_o;
  wire                majority_4842_port_o;
  wire                majority_4843_port_o;
  wire                majority_4844_port_o;
  wire                majority_4845_port_o;
  wire                majority_4846_port_o;
  wire                majority_4847_port_o;
  wire                majority_4848_port_o;
  wire                majority_4849_port_o;
  wire                majority_4850_port_o;
  wire                majority_4851_port_o;
  wire                majority_4852_port_o;
  wire                majority_4853_port_o;
  wire                majority_4854_port_o;
  wire                majority_4855_port_o;
  wire                majority_4856_port_o;
  wire                majority_4857_port_o;
  wire                majority_4858_port_o;
  wire                majority_4859_port_o;
  wire                majority_4860_port_o;
  wire                majority_4861_port_o;
  wire                majority_4862_port_o;
  wire                majority_4863_port_o;
  wire                majority_4864_port_o;
  wire                majority_4865_port_o;
  wire                majority_4866_port_o;
  wire                majority_4867_port_o;
  wire                majority_4868_port_o;
  wire                majority_4869_port_o;
  wire                majority_4870_port_o;
  wire                majority_4871_port_o;
  wire                majority_4872_port_o;
  wire                majority_4873_port_o;
  wire                majority_4874_port_o;
  wire                majority_4875_port_o;
  wire                majority_4876_port_o;
  wire                majority_4877_port_o;
  wire                majority_4878_port_o;
  wire                majority_4879_port_o;
  wire                majority_4880_port_o;
  wire                majority_4881_port_o;
  wire                majority_4882_port_o;
  wire                majority_4883_port_o;
  wire                majority_4884_port_o;
  wire                majority_4885_port_o;
  wire                majority_4886_port_o;
  wire                majority_4887_port_o;
  wire                majority_4888_port_o;
  wire                majority_4889_port_o;
  wire                majority_4890_port_o;
  wire                majority_4891_port_o;
  wire                majority_4892_port_o;
  wire                majority_4893_port_o;
  wire                majority_4894_port_o;
  wire                majority_4895_port_o;
  wire                majority_4896_port_o;
  wire                majority_4897_port_o;
  wire                majority_4898_port_o;
  wire                majority_4899_port_o;
  wire                majority_4900_port_o;
  wire                majority_4901_port_o;
  wire                majority_4902_port_o;
  wire                majority_4903_port_o;
  wire                majority_4904_port_o;
  wire                majority_4905_port_o;
  wire                majority_4906_port_o;
  wire                majority_4907_port_o;
  wire                majority_4908_port_o;
  wire                majority_4909_port_o;
  wire                majority_4910_port_o;
  wire                majority_4911_port_o;
  wire                majority_4912_port_o;
  wire                majority_4913_port_o;
  wire                majority_4914_port_o;
  wire                majority_4915_port_o;
  wire                majority_4916_port_o;
  wire                majority_4917_port_o;
  wire                majority_4918_port_o;
  wire                majority_4919_port_o;
  wire                majority_4920_port_o;
  wire                majority_4921_port_o;
  wire                majority_4922_port_o;
  wire                majority_4923_port_o;
  wire                majority_4924_port_o;
  wire                majority_4925_port_o;
  wire                majority_4926_port_o;
  wire                majority_4927_port_o;
  wire                majority_4928_port_o;
  wire                majority_4929_port_o;
  wire                majority_4930_port_o;
  wire                majority_4931_port_o;
  wire                majority_4932_port_o;
  wire                majority_4933_port_o;
  wire                majority_4934_port_o;
  wire                majority_4935_port_o;
  wire                majority_4936_port_o;
  wire                majority_4937_port_o;
  wire                majority_4938_port_o;
  wire                majority_4939_port_o;
  wire                majority_4940_port_o;
  wire                majority_4941_port_o;
  wire                majority_4942_port_o;
  wire                majority_4943_port_o;
  wire                majority_4944_port_o;
  wire                majority_4945_port_o;
  wire                majority_4946_port_o;
  wire                majority_4947_port_o;
  wire                majority_4948_port_o;
  wire                majority_4949_port_o;
  wire                majority_4950_port_o;
  wire                majority_4951_port_o;
  wire                majority_4952_port_o;
  wire                majority_4953_port_o;
  wire                majority_4954_port_o;
  wire                majority_4955_port_o;
  wire                majority_4956_port_o;
  wire                majority_4957_port_o;
  wire                majority_4958_port_o;
  wire                majority_4959_port_o;
  wire                majority_4960_port_o;
  wire                majority_4961_port_o;
  wire                majority_4962_port_o;
  wire                majority_4963_port_o;
  wire                majority_4964_port_o;
  wire                majority_4965_port_o;
  wire                majority_4966_port_o;
  wire                majority_4967_port_o;
  wire                majority_4968_port_o;
  wire                majority_4969_port_o;
  wire                majority_4970_port_o;
  wire                majority_4971_port_o;
  wire                majority_4972_port_o;
  wire                majority_4973_port_o;
  wire                majority_4974_port_o;
  wire                majority_4975_port_o;
  wire                majority_4976_port_o;
  wire                majority_4977_port_o;
  wire                majority_4978_port_o;
  wire                majority_4979_port_o;
  wire                majority_4980_port_o;
  wire                majority_4981_port_o;
  wire                majority_4982_port_o;
  wire                majority_4983_port_o;
  wire                majority_4984_port_o;
  wire                majority_4985_port_o;
  wire                majority_4986_port_o;
  wire                majority_4987_port_o;
  wire                majority_4988_port_o;
  wire                majority_4989_port_o;
  wire                majority_4990_port_o;
  wire                majority_4991_port_o;
  wire                majority_4992_port_o;
  wire                majority_4993_port_o;
  wire                majority_4994_port_o;
  wire                majority_4995_port_o;
  wire                majority_4996_port_o;
  wire                majority_4997_port_o;
  wire                majority_4998_port_o;
  wire                majority_4999_port_o;
  wire                majority_5000_port_o;
  wire                majority_5001_port_o;
  wire                majority_5002_port_o;
  wire                majority_5003_port_o;
  wire                majority_5004_port_o;
  wire                majority_5005_port_o;
  wire                majority_5006_port_o;
  wire                majority_5007_port_o;
  wire                majority_5008_port_o;
  wire                majority_5009_port_o;
  wire                majority_5010_port_o;
  wire                majority_5011_port_o;
  wire                majority_5012_port_o;
  wire                majority_5013_port_o;
  wire                majority_5014_port_o;
  wire                majority_5015_port_o;
  wire                majority_5016_port_o;
  wire                majority_5017_port_o;
  wire                majority_5018_port_o;
  wire                majority_5019_port_o;
  wire                majority_5020_port_o;
  wire                majority_5021_port_o;
  wire                majority_5022_port_o;
  wire                majority_5023_port_o;
  wire                majority_5024_port_o;
  wire                majority_5025_port_o;
  wire                majority_5026_port_o;
  wire                majority_5027_port_o;
  wire                majority_5028_port_o;
  wire                majority_5029_port_o;
  wire                majority_5030_port_o;
  wire                majority_5031_port_o;
  wire                majority_5032_port_o;
  wire                majority_5033_port_o;
  wire                majority_5034_port_o;
  wire                majority_5035_port_o;
  wire                majority_5036_port_o;
  wire                majority_5037_port_o;
  wire                majority_5038_port_o;
  wire                majority_5039_port_o;
  wire                majority_5040_port_o;
  wire                majority_5041_port_o;
  wire                majority_5042_port_o;
  wire                majority_5043_port_o;
  wire                majority_5044_port_o;
  wire                majority_5045_port_o;
  wire                majority_5046_port_o;
  wire                majority_5047_port_o;
  wire                majority_5048_port_o;
  wire                majority_5049_port_o;
  wire                majority_5050_port_o;
  wire                majority_5051_port_o;
  wire                majority_5052_port_o;
  wire                majority_5053_port_o;
  wire                majority_5054_port_o;
  wire                majority_5055_port_o;
  wire                majority_5056_port_o;
  wire                majority_5057_port_o;
  wire                majority_5058_port_o;
  wire                majority_5059_port_o;
  wire                majority_5060_port_o;
  wire                majority_5061_port_o;
  wire                majority_5062_port_o;
  wire                majority_5063_port_o;
  wire                majority_5064_port_o;
  wire                majority_5065_port_o;
  wire                majority_5066_port_o;
  wire                majority_5067_port_o;
  wire                majority_5068_port_o;
  wire                majority_5069_port_o;
  wire                majority_5070_port_o;
  wire                majority_5071_port_o;
  wire                majority_5072_port_o;
  wire                majority_5073_port_o;
  wire                majority_5074_port_o;
  wire                majority_5075_port_o;
  wire                majority_5076_port_o;
  wire                majority_5077_port_o;
  wire                majority_5078_port_o;
  wire                majority_5079_port_o;
  wire                majority_5080_port_o;
  wire                majority_5081_port_o;
  wire                majority_5082_port_o;
  wire                majority_5083_port_o;
  wire                majority_5084_port_o;
  wire                majority_5085_port_o;
  wire                majority_5086_port_o;
  wire                majority_5087_port_o;
  wire                majority_5088_port_o;
  wire                majority_5089_port_o;
  wire                majority_5090_port_o;
  wire                majority_5091_port_o;
  wire                majority_5092_port_o;
  wire                majority_5093_port_o;
  wire                majority_5094_port_o;
  wire                majority_5095_port_o;
  wire                majority_5096_port_o;
  wire                majority_5097_port_o;
  wire                majority_5098_port_o;
  wire                majority_5099_port_o;
  wire                majority_5100_port_o;
  wire                majority_5101_port_o;
  wire                majority_5102_port_o;
  wire                majority_5103_port_o;
  wire                majority_5104_port_o;
  wire                majority_5105_port_o;
  wire                majority_5106_port_o;
  wire                majority_5107_port_o;
  wire                majority_5108_port_o;
  wire                majority_5109_port_o;
  wire                majority_5110_port_o;
  wire                majority_5111_port_o;
  wire                majority_5112_port_o;
  wire                majority_5113_port_o;
  wire                majority_5114_port_o;
  wire                majority_5115_port_o;
  wire                majority_5116_port_o;
  wire                majority_5117_port_o;
  wire                majority_5118_port_o;
  wire                majority_5119_port_o;
  wire                majority_5120_port_o;
  wire                majority_5121_port_o;
  wire                majority_5122_port_o;
  wire                majority_5123_port_o;
  wire                majority_5124_port_o;
  wire                majority_5125_port_o;
  wire                majority_5126_port_o;
  wire                majority_5127_port_o;
  wire                majority_5128_port_o;
  wire                majority_5129_port_o;
  wire                majority_5130_port_o;
  wire                majority_5131_port_o;
  wire                majority_5132_port_o;
  wire                majority_5133_port_o;
  wire                majority_5134_port_o;
  wire                majority_5135_port_o;
  wire                majority_5136_port_o;
  wire                majority_5137_port_o;
  wire                majority_5138_port_o;
  wire                majority_5139_port_o;
  wire                majority_5140_port_o;
  wire                majority_5141_port_o;
  wire                majority_5142_port_o;
  wire                majority_5143_port_o;
  wire                majority_5144_port_o;
  wire                majority_5145_port_o;
  wire                majority_5146_port_o;
  wire                majority_5147_port_o;
  wire                majority_5148_port_o;
  wire                majority_5149_port_o;
  wire                majority_5150_port_o;
  wire                majority_5151_port_o;
  wire                majority_5152_port_o;
  wire                majority_5153_port_o;
  wire                majority_5154_port_o;
  wire                majority_5155_port_o;
  wire                majority_5156_port_o;
  wire                majority_5157_port_o;
  wire                majority_5158_port_o;
  wire                majority_5159_port_o;
  wire                majority_5160_port_o;
  wire                majority_5161_port_o;
  wire                majority_5162_port_o;
  wire                majority_5163_port_o;
  wire                majority_5164_port_o;
  wire                majority_5165_port_o;
  wire                majority_5166_port_o;
  wire                majority_5167_port_o;
  wire                majority_5168_port_o;
  wire                majority_5169_port_o;
  wire                majority_5170_port_o;
  wire                majority_5171_port_o;
  wire                majority_5172_port_o;
  wire                majority_5173_port_o;
  wire                majority_5174_port_o;
  wire                majority_5175_port_o;
  wire                majority_5176_port_o;
  wire                majority_5177_port_o;
  wire                majority_5178_port_o;
  wire                majority_5179_port_o;
  wire                majority_5180_port_o;
  wire                majority_5181_port_o;
  wire                majority_5182_port_o;
  wire                majority_5183_port_o;
  wire                majority_5184_port_o;
  wire                majority_5185_port_o;
  wire                majority_5186_port_o;
  wire                majority_5187_port_o;
  wire                majority_5188_port_o;
  wire                majority_5189_port_o;
  wire                majority_5190_port_o;
  wire                majority_5191_port_o;
  wire                majority_5192_port_o;
  wire                majority_5193_port_o;
  wire                majority_5194_port_o;
  wire                majority_5195_port_o;
  wire                majority_5196_port_o;
  wire                majority_5197_port_o;
  wire                majority_5198_port_o;
  wire                majority_5199_port_o;
  wire                majority_5200_port_o;
  wire                majority_5201_port_o;
  wire                majority_5202_port_o;
  wire                majority_5203_port_o;
  wire                majority_5204_port_o;
  wire                majority_5205_port_o;
  wire                majority_5206_port_o;
  wire                majority_5207_port_o;
  wire                majority_5208_port_o;
  wire                majority_5209_port_o;
  wire                majority_5210_port_o;
  wire                majority_5211_port_o;
  wire                majority_5212_port_o;
  wire                majority_5213_port_o;
  wire                majority_5214_port_o;
  wire                majority_5215_port_o;
  wire                majority_5216_port_o;
  wire                majority_5217_port_o;
  wire                majority_5218_port_o;
  wire                majority_5219_port_o;
  wire                majority_5220_port_o;
  wire                majority_5221_port_o;
  wire                majority_5222_port_o;
  wire                majority_5223_port_o;
  wire                majority_5224_port_o;
  wire                majority_5225_port_o;
  wire                majority_5226_port_o;
  wire                majority_5227_port_o;
  wire                majority_5228_port_o;
  wire                majority_5229_port_o;
  wire                majority_5230_port_o;
  wire                majority_5231_port_o;
  wire                majority_5232_port_o;
  wire                majority_5233_port_o;
  wire                majority_5234_port_o;
  wire                majority_5235_port_o;
  wire                majority_5236_port_o;
  wire                majority_5237_port_o;
  wire                majority_5238_port_o;
  wire                majority_5239_port_o;
  wire                majority_5240_port_o;
  wire                majority_5241_port_o;
  wire                majority_5242_port_o;
  wire                majority_5243_port_o;
  wire                majority_5244_port_o;
  wire                majority_5245_port_o;
  wire                majority_5246_port_o;
  wire                majority_5247_port_o;
  wire                majority_5248_port_o;
  wire                majority_5249_port_o;
  wire                majority_5250_port_o;
  wire                majority_5251_port_o;
  wire                majority_5252_port_o;
  wire                majority_5253_port_o;
  wire                majority_5254_port_o;
  wire                majority_5255_port_o;
  wire                majority_5256_port_o;
  wire                majority_5257_port_o;
  wire                majority_5258_port_o;
  wire                majority_5259_port_o;
  wire                majority_5260_port_o;
  wire                majority_5261_port_o;
  wire                majority_5262_port_o;
  wire                majority_5263_port_o;
  wire                majority_5264_port_o;
  wire                majority_5265_port_o;
  wire                majority_5266_port_o;
  wire                majority_5267_port_o;
  wire                majority_5268_port_o;
  wire                majority_5269_port_o;
  wire                majority_5270_port_o;
  wire                majority_5271_port_o;
  wire                majority_5272_port_o;
  wire                majority_5273_port_o;
  wire                majority_5274_port_o;
  wire                majority_5275_port_o;
  wire                majority_5276_port_o;
  wire                majority_5277_port_o;
  wire                majority_5278_port_o;
  wire                majority_5279_port_o;
  wire                majority_5280_port_o;
  wire                majority_5281_port_o;
  wire                majority_5282_port_o;
  wire                majority_5283_port_o;
  wire                majority_5284_port_o;
  wire                majority_5285_port_o;
  wire                majority_5286_port_o;
  wire                majority_5287_port_o;
  wire                majority_5288_port_o;
  wire                majority_5289_port_o;
  wire                majority_5290_port_o;
  wire                majority_5291_port_o;
  wire                majority_5292_port_o;
  wire                majority_5293_port_o;
  wire                majority_5294_port_o;
  wire                majority_5295_port_o;
  wire                majority_5296_port_o;
  wire                majority_5297_port_o;
  wire                majority_5298_port_o;
  wire                majority_5299_port_o;
  wire                majority_5300_port_o;
  wire                majority_5301_port_o;
  wire                majority_5302_port_o;
  wire                majority_5303_port_o;
  wire                majority_5304_port_o;
  wire                majority_5305_port_o;
  wire                majority_5306_port_o;
  wire                majority_5307_port_o;
  wire                majority_5308_port_o;
  wire                majority_5309_port_o;
  wire                majority_5310_port_o;
  wire                majority_5311_port_o;
  wire                majority_5312_port_o;
  wire                majority_5313_port_o;
  wire                majority_5314_port_o;
  wire                majority_5315_port_o;
  wire                majority_5316_port_o;
  wire                majority_5317_port_o;
  wire                majority_5318_port_o;
  wire                majority_5319_port_o;
  wire                majority_5320_port_o;
  wire                majority_5321_port_o;
  wire                majority_5322_port_o;
  wire                majority_5323_port_o;
  wire                majority_5324_port_o;
  wire                majority_5325_port_o;
  wire                majority_5326_port_o;
  wire                majority_5327_port_o;
  wire                majority_5328_port_o;
  wire                majority_5329_port_o;
  wire                majority_5330_port_o;
  wire                majority_5331_port_o;
  wire                majority_5332_port_o;
  wire                majority_5333_port_o;
  wire                majority_5334_port_o;
  wire                majority_5335_port_o;
  wire                majority_5336_port_o;
  wire                majority_5337_port_o;
  wire                majority_5338_port_o;
  wire                majority_5339_port_o;
  wire                majority_5340_port_o;
  wire                majority_5341_port_o;
  wire                majority_5342_port_o;
  wire                majority_5343_port_o;
  wire                majority_5344_port_o;
  wire                majority_5345_port_o;
  wire                majority_5346_port_o;
  wire                majority_5347_port_o;
  wire                majority_5348_port_o;
  wire                majority_5349_port_o;
  wire                majority_5350_port_o;
  wire                majority_5351_port_o;
  wire                majority_5352_port_o;
  wire                majority_5353_port_o;
  wire                majority_5354_port_o;
  wire                majority_5355_port_o;
  wire                majority_5356_port_o;
  wire                majority_5357_port_o;
  wire                majority_5358_port_o;
  wire                majority_5359_port_o;
  wire                majority_5360_port_o;
  wire                majority_5361_port_o;
  wire                majority_5362_port_o;
  wire                majority_5363_port_o;
  wire                majority_5364_port_o;
  wire                majority_5365_port_o;
  wire                majority_5366_port_o;
  wire                majority_5367_port_o;
  wire                majority_5368_port_o;
  wire                majority_5369_port_o;
  wire                majority_5370_port_o;
  wire                majority_5371_port_o;
  wire                majority_5372_port_o;
  wire                majority_5373_port_o;
  wire                majority_5374_port_o;
  wire                majority_5375_port_o;
  wire                majority_5376_port_o;
  wire                majority_5377_port_o;
  wire                majority_5378_port_o;
  wire                majority_5379_port_o;
  wire                majority_5380_port_o;
  wire                majority_5381_port_o;
  wire                majority_5382_port_o;
  wire                majority_5383_port_o;
  wire                majority_5384_port_o;
  wire                majority_5385_port_o;
  wire                majority_5386_port_o;
  wire                majority_5387_port_o;
  wire                majority_5388_port_o;
  wire                majority_5389_port_o;
  wire                majority_5390_port_o;
  wire                majority_5391_port_o;
  wire                majority_5392_port_o;
  wire                majority_5393_port_o;
  wire                majority_5394_port_o;
  wire                majority_5395_port_o;
  wire                majority_5396_port_o;
  wire                majority_5397_port_o;
  wire                majority_5398_port_o;
  wire                majority_5399_port_o;
  wire                majority_5400_port_o;
  wire                majority_5401_port_o;
  wire                majority_5402_port_o;
  wire                majority_5403_port_o;
  wire                majority_5404_port_o;
  wire                majority_5405_port_o;
  wire                majority_5406_port_o;
  wire                majority_5407_port_o;
  wire                majority_5408_port_o;
  wire                majority_5409_port_o;
  wire                majority_5410_port_o;
  wire                majority_5411_port_o;
  wire                majority_5412_port_o;
  wire                majority_5413_port_o;
  wire                majority_5414_port_o;
  wire                majority_5415_port_o;
  wire                majority_5416_port_o;
  wire                majority_5417_port_o;
  wire                majority_5418_port_o;
  wire                majority_5419_port_o;
  wire                majority_5420_port_o;
  wire                majority_5421_port_o;
  wire                majority_5422_port_o;
  wire                majority_5423_port_o;
  wire                majority_5424_port_o;
  wire                majority_5425_port_o;
  wire                majority_5426_port_o;
  wire                majority_5427_port_o;
  wire                majority_5428_port_o;
  wire                majority_5429_port_o;
  wire                majority_5430_port_o;
  wire                majority_5431_port_o;
  wire                majority_5432_port_o;
  wire                majority_5433_port_o;
  wire                majority_5434_port_o;
  wire                majority_5435_port_o;
  wire                majority_5436_port_o;
  wire                majority_5437_port_o;
  wire                majority_5438_port_o;
  wire                majority_5439_port_o;
  wire                majority_5440_port_o;
  wire                majority_5441_port_o;
  wire                majority_5442_port_o;
  wire                majority_5443_port_o;
  wire                majority_5444_port_o;
  wire                majority_5445_port_o;
  wire                majority_5446_port_o;
  wire                majority_5447_port_o;
  wire                majority_5448_port_o;
  wire                majority_5449_port_o;
  wire                majority_5450_port_o;
  wire                majority_5451_port_o;
  wire                majority_5452_port_o;
  wire                majority_5453_port_o;
  wire                majority_5454_port_o;
  wire                majority_5455_port_o;
  wire                majority_5456_port_o;
  wire                majority_5457_port_o;
  wire                majority_5458_port_o;
  wire                majority_5459_port_o;
  wire                majority_5460_port_o;
  wire                majority_5461_port_o;
  wire                majority_5462_port_o;
  wire                majority_5463_port_o;
  wire                majority_5464_port_o;
  wire                majority_5465_port_o;
  wire                majority_5466_port_o;
  wire                majority_5467_port_o;
  wire                majority_5468_port_o;
  wire                majority_5469_port_o;
  wire                majority_5470_port_o;
  wire                majority_5471_port_o;
  wire                majority_5472_port_o;
  wire                majority_5473_port_o;
  wire                majority_5474_port_o;
  wire                majority_5475_port_o;
  wire                majority_5476_port_o;
  wire                majority_5477_port_o;
  wire                majority_5478_port_o;
  wire                majority_5479_port_o;
  wire                majority_5480_port_o;
  wire                majority_5481_port_o;
  wire                majority_5482_port_o;
  wire                majority_5483_port_o;
  wire                majority_5484_port_o;
  wire                majority_5485_port_o;
  wire                majority_5486_port_o;
  wire                majority_5487_port_o;
  wire                majority_5488_port_o;
  wire                majority_5489_port_o;
  wire                majority_5490_port_o;
  wire                majority_5491_port_o;
  wire                majority_5492_port_o;
  wire                majority_5493_port_o;
  wire                majority_5494_port_o;
  wire                majority_5495_port_o;
  wire                majority_5496_port_o;
  wire                majority_5497_port_o;
  wire                majority_5498_port_o;
  wire                majority_5499_port_o;
  wire                majority_5500_port_o;
  wire                majority_5501_port_o;
  wire                majority_5502_port_o;
  wire                majority_5503_port_o;
  wire                majority_5504_port_o;
  wire                majority_5505_port_o;
  wire                majority_5506_port_o;
  wire                majority_5507_port_o;
  wire                majority_5508_port_o;
  wire                majority_5509_port_o;
  wire                majority_5510_port_o;
  wire                majority_5511_port_o;
  wire                majority_5512_port_o;
  wire                majority_5513_port_o;
  wire                majority_5514_port_o;
  wire                majority_5515_port_o;
  wire                majority_5516_port_o;
  wire                majority_5517_port_o;
  wire                majority_5518_port_o;
  wire                majority_5519_port_o;
  wire                majority_5520_port_o;
  wire                majority_5521_port_o;
  wire                majority_5522_port_o;
  wire                majority_5523_port_o;
  wire                majority_5524_port_o;
  wire                majority_5525_port_o;
  wire                majority_5526_port_o;
  wire                majority_5527_port_o;
  wire                majority_5528_port_o;
  wire                majority_5529_port_o;
  wire                majority_5530_port_o;
  wire                majority_5531_port_o;
  wire                majority_5532_port_o;
  wire                majority_5533_port_o;
  wire                majority_5534_port_o;
  wire                majority_5535_port_o;
  wire                majority_5536_port_o;
  wire                majority_5537_port_o;
  wire                majority_5538_port_o;
  wire                majority_5539_port_o;
  wire                majority_5540_port_o;
  wire                majority_5541_port_o;
  wire                majority_5542_port_o;
  wire                majority_5543_port_o;
  wire                majority_5544_port_o;
  wire                majority_5545_port_o;
  wire                majority_5546_port_o;
  wire                majority_5547_port_o;
  wire                majority_5548_port_o;
  wire                majority_5549_port_o;
  wire                majority_5550_port_o;
  wire                majority_5551_port_o;
  wire                majority_5552_port_o;
  wire                majority_5553_port_o;
  wire                majority_5554_port_o;
  wire                majority_5555_port_o;
  wire                majority_5556_port_o;
  wire                majority_5557_port_o;
  wire                majority_5558_port_o;
  wire                majority_5559_port_o;
  wire                majority_5560_port_o;
  wire                majority_5561_port_o;
  wire                majority_5562_port_o;
  wire                majority_5563_port_o;
  wire                majority_5564_port_o;
  wire                majority_5565_port_o;
  wire                majority_5566_port_o;
  wire                majority_5567_port_o;
  wire                majority_5568_port_o;
  wire                majority_5569_port_o;
  wire                majority_5570_port_o;
  wire                majority_5571_port_o;
  wire                majority_5572_port_o;
  wire                majority_5573_port_o;
  wire                majority_5574_port_o;
  wire                majority_5575_port_o;
  wire                majority_5576_port_o;
  wire                majority_5577_port_o;
  wire                majority_5578_port_o;
  wire                majority_5579_port_o;
  wire                majority_5580_port_o;
  wire                majority_5581_port_o;
  wire                majority_5582_port_o;
  wire                majority_5583_port_o;
  wire                majority_5584_port_o;
  wire                majority_5585_port_o;
  wire                majority_5586_port_o;
  wire                majority_5587_port_o;
  wire                majority_5588_port_o;
  wire                majority_5589_port_o;
  wire                majority_5590_port_o;
  wire                majority_5591_port_o;
  wire                majority_5592_port_o;
  wire                majority_5593_port_o;
  wire                majority_5594_port_o;
  wire                majority_5595_port_o;
  wire                majority_5596_port_o;
  wire                majority_5597_port_o;
  wire                majority_5598_port_o;
  wire                majority_5599_port_o;
  wire                majority_5600_port_o;
  wire                majority_5601_port_o;
  wire                majority_5602_port_o;
  wire                majority_5603_port_o;
  wire                majority_5604_port_o;
  wire                majority_5605_port_o;
  wire                majority_5606_port_o;
  wire                majority_5607_port_o;
  wire                majority_5608_port_o;
  wire                majority_5609_port_o;
  wire                majority_5610_port_o;
  wire                majority_5611_port_o;
  wire                majority_5612_port_o;
  wire                majority_5613_port_o;
  wire                majority_5614_port_o;
  wire                majority_5615_port_o;
  wire                majority_5616_port_o;
  wire                majority_5617_port_o;
  wire                majority_5618_port_o;
  wire                majority_5619_port_o;
  wire                majority_5620_port_o;
  wire                majority_5621_port_o;
  wire                majority_5622_port_o;
  wire                majority_5623_port_o;
  wire                majority_5624_port_o;
  wire                majority_5625_port_o;
  wire                majority_5626_port_o;
  wire                majority_5627_port_o;
  wire                majority_5628_port_o;
  wire                majority_5629_port_o;
  wire                majority_5630_port_o;
  wire                majority_5631_port_o;
  wire                majority_5632_port_o;
  wire                majority_5633_port_o;
  wire                majority_5634_port_o;
  wire                majority_5635_port_o;
  wire                majority_5636_port_o;
  wire                majority_5637_port_o;
  wire                majority_5638_port_o;
  wire                majority_5639_port_o;
  wire                majority_5640_port_o;
  wire                majority_5641_port_o;
  wire                majority_5642_port_o;
  wire                majority_5643_port_o;
  wire                majority_5644_port_o;
  wire                majority_5645_port_o;
  wire                majority_5646_port_o;
  wire                majority_5647_port_o;
  wire                majority_5648_port_o;
  wire                majority_5649_port_o;
  wire                majority_5650_port_o;
  wire                majority_5651_port_o;
  wire                majority_5652_port_o;
  wire                majority_5653_port_o;
  wire                majority_5654_port_o;
  wire                majority_5655_port_o;
  wire                majority_5656_port_o;
  wire                majority_5657_port_o;
  wire                majority_5658_port_o;
  wire                majority_5659_port_o;
  wire                majority_5660_port_o;
  wire                majority_5661_port_o;
  wire                majority_5662_port_o;
  wire                majority_5663_port_o;
  wire                majority_5664_port_o;
  wire                majority_5665_port_o;
  wire                majority_5666_port_o;
  wire                majority_5667_port_o;
  wire                majority_5668_port_o;
  wire                majority_5669_port_o;
  wire                majority_5670_port_o;
  wire                majority_5671_port_o;
  wire                majority_5672_port_o;
  wire                majority_5673_port_o;
  wire                majority_5674_port_o;
  wire                majority_5675_port_o;
  wire                majority_5676_port_o;
  wire                majority_5677_port_o;
  wire                majority_5678_port_o;
  wire                majority_5679_port_o;
  wire                majority_5680_port_o;
  wire                majority_5681_port_o;
  wire                majority_5682_port_o;
  wire                majority_5683_port_o;
  wire                majority_5684_port_o;
  wire                majority_5685_port_o;
  wire                majority_5686_port_o;
  wire                majority_5687_port_o;
  wire                majority_5688_port_o;
  wire                majority_5689_port_o;
  wire                majority_5690_port_o;
  wire                majority_5691_port_o;
  wire                majority_5692_port_o;
  wire                majority_5693_port_o;
  wire                majority_5694_port_o;
  wire                majority_5695_port_o;
  wire                majority_5696_port_o;
  wire                majority_5697_port_o;
  wire                majority_5698_port_o;
  wire                majority_5699_port_o;
  wire                majority_5700_port_o;
  wire                majority_5701_port_o;
  wire                majority_5702_port_o;
  wire                majority_5703_port_o;
  wire                majority_5704_port_o;
  wire                majority_5705_port_o;
  wire                majority_5706_port_o;
  wire                majority_5707_port_o;
  wire                majority_5708_port_o;
  wire                majority_5709_port_o;
  wire                majority_5710_port_o;
  wire                majority_5711_port_o;
  wire                majority_5712_port_o;
  wire                majority_5713_port_o;
  wire                majority_5714_port_o;
  wire                majority_5715_port_o;
  wire                majority_5716_port_o;
  wire                majority_5717_port_o;
  wire                majority_5718_port_o;
  wire                majority_5719_port_o;
  wire                majority_5720_port_o;
  wire                majority_5721_port_o;
  wire                majority_5722_port_o;
  wire                majority_5723_port_o;
  wire                majority_5724_port_o;
  wire                majority_5725_port_o;
  wire                majority_5726_port_o;
  wire                majority_5727_port_o;
  wire                majority_5728_port_o;
  wire                majority_5729_port_o;
  wire                majority_5730_port_o;
  wire                majority_5731_port_o;
  wire                majority_5732_port_o;
  wire                majority_5733_port_o;
  wire                majority_5734_port_o;
  wire                majority_5735_port_o;
  wire                majority_5736_port_o;
  wire                majority_5737_port_o;
  wire                majority_5738_port_o;
  wire                majority_5739_port_o;
  wire                majority_5740_port_o;
  wire                majority_5741_port_o;
  wire                majority_5742_port_o;
  wire                majority_5743_port_o;
  wire                majority_5744_port_o;
  wire                majority_5745_port_o;
  wire                majority_5746_port_o;
  wire                majority_5747_port_o;
  wire                majority_5748_port_o;
  wire                majority_5749_port_o;
  wire                majority_5750_port_o;
  wire                majority_5751_port_o;
  wire                majority_5752_port_o;
  wire                majority_5753_port_o;
  wire                majority_5754_port_o;
  wire                majority_5755_port_o;
  wire                majority_5756_port_o;
  wire                majority_5757_port_o;
  wire                majority_5758_port_o;
  wire                majority_5759_port_o;
  wire                majority_5760_port_o;
  wire                majority_5761_port_o;
  wire                majority_5762_port_o;
  wire                majority_5763_port_o;
  wire                majority_5764_port_o;
  wire                majority_5765_port_o;
  wire                majority_5766_port_o;
  wire                majority_5767_port_o;
  wire                majority_5768_port_o;
  wire                majority_5769_port_o;
  wire                majority_5770_port_o;
  wire                majority_5771_port_o;
  wire                majority_5772_port_o;
  wire                majority_5773_port_o;
  wire                majority_5774_port_o;
  wire                majority_5775_port_o;
  wire                majority_5776_port_o;
  wire                majority_5777_port_o;
  wire                majority_5778_port_o;
  wire                majority_5779_port_o;
  wire                majority_5780_port_o;
  wire                majority_5781_port_o;
  wire                majority_5782_port_o;
  wire                majority_5783_port_o;
  wire                majority_5784_port_o;
  wire                majority_5785_port_o;
  wire                majority_5786_port_o;
  wire                majority_5787_port_o;
  wire                majority_5788_port_o;
  wire                majority_5789_port_o;
  wire                majority_5790_port_o;
  wire                majority_5791_port_o;
  wire                majority_5792_port_o;
  wire                majority_5793_port_o;
  wire                majority_5794_port_o;
  wire                majority_5795_port_o;
  wire                majority_5796_port_o;
  wire                majority_5797_port_o;
  wire                majority_5798_port_o;
  wire                majority_5799_port_o;
  wire                majority_5800_port_o;
  wire                majority_5801_port_o;
  wire                majority_5802_port_o;
  wire                majority_5803_port_o;
  wire                majority_5804_port_o;
  wire                majority_5805_port_o;
  wire                majority_5806_port_o;
  wire                majority_5807_port_o;
  wire                majority_5808_port_o;
  wire                majority_5809_port_o;
  wire                majority_5810_port_o;
  wire                majority_5811_port_o;
  wire                majority_5812_port_o;
  wire                majority_5813_port_o;
  wire                majority_5814_port_o;
  wire                majority_5815_port_o;
  wire                majority_5816_port_o;
  wire                majority_5817_port_o;
  wire                majority_5818_port_o;
  wire                majority_5819_port_o;
  wire                majority_5820_port_o;
  wire                majority_5821_port_o;
  wire                majority_5822_port_o;
  wire                majority_5823_port_o;
  wire                majority_5824_port_o;
  wire                majority_5825_port_o;
  wire                majority_5826_port_o;
  wire                majority_5827_port_o;
  wire                majority_5828_port_o;
  wire                majority_5829_port_o;
  wire                majority_5830_port_o;
  wire                majority_5831_port_o;
  wire                majority_5832_port_o;
  wire                majority_5833_port_o;
  wire                majority_5834_port_o;
  wire                majority_5835_port_o;
  wire                majority_5836_port_o;
  wire                majority_5837_port_o;
  wire                majority_5838_port_o;
  wire                majority_5839_port_o;
  wire                majority_5840_port_o;
  wire                majority_5841_port_o;
  wire                majority_5842_port_o;
  wire                majority_5843_port_o;
  wire                majority_5844_port_o;
  wire                majority_5845_port_o;
  wire                majority_5846_port_o;
  wire                majority_5847_port_o;
  wire                majority_5848_port_o;
  wire                majority_5849_port_o;
  wire                majority_5850_port_o;
  wire                majority_5851_port_o;
  wire                majority_5852_port_o;
  wire                majority_5853_port_o;
  wire                majority_5854_port_o;
  wire                majority_5855_port_o;
  wire                majority_5856_port_o;
  wire                majority_5857_port_o;
  wire                majority_5858_port_o;
  wire                majority_5859_port_o;
  wire                majority_5860_port_o;
  wire                majority_5861_port_o;
  wire                majority_5862_port_o;
  wire                majority_5863_port_o;
  wire                majority_5864_port_o;
  wire                majority_5865_port_o;
  wire                majority_5866_port_o;
  wire                majority_5867_port_o;
  wire                majority_5868_port_o;
  wire                majority_5869_port_o;
  wire                majority_5870_port_o;
  wire                majority_5871_port_o;
  wire                majority_5872_port_o;
  wire                majority_5873_port_o;
  wire                majority_5874_port_o;
  wire                majority_5875_port_o;
  wire                majority_5876_port_o;
  wire                majority_5877_port_o;
  wire                majority_5878_port_o;
  wire                majority_5879_port_o;
  wire                majority_5880_port_o;
  wire                majority_5881_port_o;
  wire                majority_5882_port_o;
  wire                majority_5883_port_o;
  wire                majority_5884_port_o;
  wire                majority_5885_port_o;
  wire                majority_5886_port_o;
  wire                majority_5887_port_o;
  wire                majority_5888_port_o;
  wire                majority_5889_port_o;
  wire                majority_5890_port_o;
  wire                majority_5891_port_o;
  wire                majority_5892_port_o;
  wire                majority_5893_port_o;
  wire                majority_5894_port_o;
  wire                majority_5895_port_o;
  wire                majority_5896_port_o;
  wire                majority_5897_port_o;
  wire                majority_5898_port_o;
  wire                majority_5899_port_o;
  wire                majority_5900_port_o;
  wire                majority_5901_port_o;
  wire                majority_5902_port_o;
  wire                majority_5903_port_o;
  wire                majority_5904_port_o;
  wire                majority_5905_port_o;
  wire                majority_5906_port_o;
  wire                majority_5907_port_o;
  wire                majority_5908_port_o;
  wire                majority_5909_port_o;
  wire                majority_5910_port_o;
  wire                majority_5911_port_o;
  wire                majority_5912_port_o;
  wire                majority_5913_port_o;
  wire                majority_5914_port_o;
  wire                majority_5915_port_o;
  wire                majority_5916_port_o;
  wire                majority_5917_port_o;
  wire                majority_5918_port_o;
  wire                majority_5919_port_o;
  wire                majority_5920_port_o;
  wire                majority_5921_port_o;
  wire                majority_5922_port_o;
  wire                majority_5923_port_o;
  wire                majority_5924_port_o;
  wire                majority_5925_port_o;
  wire                majority_5926_port_o;
  wire                majority_5927_port_o;
  wire                majority_5928_port_o;
  wire                majority_5929_port_o;
  wire                majority_5930_port_o;
  wire                majority_5931_port_o;
  wire                majority_5932_port_o;
  wire                majority_5933_port_o;
  wire                majority_5934_port_o;
  wire                majority_5935_port_o;
  wire                majority_5936_port_o;
  wire                majority_5937_port_o;
  wire                majority_5938_port_o;
  wire                majority_5939_port_o;
  wire                majority_5940_port_o;
  wire                majority_5941_port_o;
  wire                majority_5942_port_o;
  wire                majority_5943_port_o;
  wire                majority_5944_port_o;
  wire                majority_5945_port_o;
  wire                majority_5946_port_o;
  wire                majority_5947_port_o;
  wire                majority_5948_port_o;
  wire                majority_5949_port_o;
  wire                majority_5950_port_o;
  wire                majority_5951_port_o;
  wire                majority_5952_port_o;
  wire                majority_5953_port_o;
  wire                majority_5954_port_o;
  wire                majority_5955_port_o;
  wire                majority_5956_port_o;
  wire                majority_5957_port_o;
  wire                majority_5958_port_o;
  wire                majority_5959_port_o;
  wire                majority_5960_port_o;
  wire                majority_5961_port_o;
  wire                majority_5962_port_o;
  wire                majority_5963_port_o;
  wire                majority_5964_port_o;
  wire                majority_5965_port_o;
  wire                majority_5966_port_o;
  wire                majority_5967_port_o;
  wire                majority_5968_port_o;
  wire                majority_5969_port_o;
  wire                majority_5970_port_o;
  wire                majority_5971_port_o;
  wire                majority_5972_port_o;
  wire                majority_5973_port_o;
  wire                majority_5974_port_o;
  wire                majority_5975_port_o;
  wire                majority_5976_port_o;
  wire                majority_5977_port_o;
  wire                majority_5978_port_o;
  wire                majority_5979_port_o;
  wire                majority_5980_port_o;
  wire                majority_5981_port_o;
  wire                majority_5982_port_o;
  wire                majority_5983_port_o;
  wire                majority_5984_port_o;
  wire                majority_5985_port_o;
  wire                majority_5986_port_o;
  wire                majority_5987_port_o;
  wire                majority_5988_port_o;
  wire                majority_5989_port_o;
  wire                majority_5990_port_o;
  wire                majority_5991_port_o;
  wire                majority_5992_port_o;
  wire                majority_5993_port_o;
  wire                majority_5994_port_o;
  wire                majority_5995_port_o;
  wire                majority_5996_port_o;
  wire                majority_5997_port_o;
  wire                majority_5998_port_o;
  wire                majority_5999_port_o;
  wire                majority_6000_port_o;
  wire                majority_6001_port_o;
  wire                majority_6002_port_o;
  wire                majority_6003_port_o;
  wire                majority_6004_port_o;
  wire                majority_6005_port_o;
  wire                majority_6006_port_o;
  wire                majority_6007_port_o;
  wire                majority_6008_port_o;
  wire                majority_6009_port_o;
  wire                majority_6010_port_o;
  wire                majority_6011_port_o;
  wire                majority_6012_port_o;
  wire                majority_6013_port_o;
  wire                majority_6014_port_o;
  wire                majority_6015_port_o;
  wire                majority_6016_port_o;
  wire                majority_6017_port_o;
  wire                majority_6018_port_o;
  wire                majority_6019_port_o;
  wire                majority_6020_port_o;
  wire                majority_6021_port_o;
  wire                majority_6022_port_o;
  wire                majority_6023_port_o;
  wire                majority_6024_port_o;
  wire                majority_6025_port_o;
  wire                majority_6026_port_o;
  wire                majority_6027_port_o;
  wire                majority_6028_port_o;
  wire                majority_6029_port_o;
  wire                majority_6030_port_o;
  wire                majority_6031_port_o;
  wire                majority_6032_port_o;
  wire                majority_6033_port_o;
  wire                majority_6034_port_o;
  wire                majority_6035_port_o;
  wire                majority_6036_port_o;
  wire                majority_6037_port_o;
  wire                majority_6038_port_o;
  wire                majority_6039_port_o;
  wire                majority_6040_port_o;
  wire                majority_6041_port_o;
  wire                majority_6042_port_o;
  wire                majority_6043_port_o;
  wire                majority_6044_port_o;
  wire                majority_6045_port_o;
  wire                majority_6046_port_o;
  wire                majority_6047_port_o;
  wire                majority_6048_port_o;
  wire                majority_6049_port_o;
  wire                majority_6050_port_o;
  wire                majority_6051_port_o;
  wire                majority_6052_port_o;
  wire                majority_6053_port_o;
  wire                majority_6054_port_o;
  wire                majority_6055_port_o;
  wire                majority_6056_port_o;
  wire                majority_6057_port_o;
  wire                majority_6058_port_o;
  wire                majority_6059_port_o;
  wire                majority_6060_port_o;
  wire                majority_6061_port_o;
  wire                majority_6062_port_o;
  wire                majority_6063_port_o;
  wire                majority_6064_port_o;
  wire                majority_6065_port_o;
  wire                majority_6066_port_o;
  wire                majority_6067_port_o;
  wire                majority_6068_port_o;
  wire                majority_6069_port_o;
  wire                majority_6070_port_o;
  wire                majority_6071_port_o;
  wire                majority_6072_port_o;
  wire                majority_6073_port_o;
  wire                majority_6074_port_o;
  wire                majority_6075_port_o;
  wire                majority_6076_port_o;
  wire                majority_6077_port_o;
  wire                majority_6078_port_o;
  wire                majority_6079_port_o;
  wire                majority_6080_port_o;
  wire                majority_6081_port_o;
  wire                majority_6082_port_o;
  wire                majority_6083_port_o;
  wire                majority_6084_port_o;
  wire                majority_6085_port_o;
  wire                majority_6086_port_o;
  wire                majority_6087_port_o;
  wire                majority_6088_port_o;
  wire                majority_6089_port_o;
  wire                majority_6090_port_o;
  wire                majority_6091_port_o;
  wire                majority_6092_port_o;
  wire                majority_6093_port_o;
  wire                majority_6094_port_o;
  wire                majority_6095_port_o;
  wire                majority_6096_port_o;
  wire                majority_6097_port_o;
  wire                majority_6098_port_o;
  wire                majority_6099_port_o;
  wire                majority_6100_port_o;
  wire                majority_6101_port_o;
  wire                majority_6102_port_o;
  wire                majority_6103_port_o;
  wire                majority_6104_port_o;
  wire                majority_6105_port_o;
  wire                majority_6106_port_o;
  wire                majority_6107_port_o;
  wire                majority_6108_port_o;
  wire                majority_6109_port_o;
  wire                majority_6110_port_o;
  wire                majority_6111_port_o;
  wire                majority_6112_port_o;
  wire                majority_6113_port_o;
  wire                majority_6114_port_o;
  wire                majority_6115_port_o;
  wire                majority_6116_port_o;
  wire                majority_6117_port_o;
  wire                majority_6118_port_o;
  wire                majority_6119_port_o;
  wire                majority_6120_port_o;
  wire                majority_6121_port_o;
  wire                majority_6122_port_o;
  wire                majority_6123_port_o;
  wire                majority_6124_port_o;
  wire                majority_6125_port_o;
  wire                majority_6126_port_o;
  wire                majority_6127_port_o;
  wire                majority_6128_port_o;
  wire                majority_6129_port_o;
  wire                majority_6130_port_o;
  wire                majority_6131_port_o;
  wire                majority_6132_port_o;
  wire                majority_6133_port_o;
  wire                majority_6134_port_o;
  wire                majority_6135_port_o;
  wire                majority_6136_port_o;
  wire                majority_6137_port_o;
  wire                majority_6138_port_o;
  wire                majority_6139_port_o;
  wire                majority_6140_port_o;
  wire                majority_6141_port_o;
  wire                majority_6142_port_o;
  wire                majority_6143_port_o;
  wire       [2:0]    subBytes_out_0_0_0;
  wire       [2:0]    subBytes_out_0_0_1;
  wire       [2:0]    subBytes_out_0_0_2;
  wire       [2:0]    subBytes_out_0_0_3;
  wire       [2:0]    subBytes_out_0_0_4;
  wire       [2:0]    subBytes_out_0_0_5;
  wire       [2:0]    subBytes_out_0_0_6;
  wire       [2:0]    subBytes_out_0_0_7;
  wire       [2:0]    subBytes_out_0_1_0;
  wire       [2:0]    subBytes_out_0_1_1;
  wire       [2:0]    subBytes_out_0_1_2;
  wire       [2:0]    subBytes_out_0_1_3;
  wire       [2:0]    subBytes_out_0_1_4;
  wire       [2:0]    subBytes_out_0_1_5;
  wire       [2:0]    subBytes_out_0_1_6;
  wire       [2:0]    subBytes_out_0_1_7;
  wire       [2:0]    subBytes_out_0_2_0;
  wire       [2:0]    subBytes_out_0_2_1;
  wire       [2:0]    subBytes_out_0_2_2;
  wire       [2:0]    subBytes_out_0_2_3;
  wire       [2:0]    subBytes_out_0_2_4;
  wire       [2:0]    subBytes_out_0_2_5;
  wire       [2:0]    subBytes_out_0_2_6;
  wire       [2:0]    subBytes_out_0_2_7;
  wire       [2:0]    subBytes_out_0_3_0;
  wire       [2:0]    subBytes_out_0_3_1;
  wire       [2:0]    subBytes_out_0_3_2;
  wire       [2:0]    subBytes_out_0_3_3;
  wire       [2:0]    subBytes_out_0_3_4;
  wire       [2:0]    subBytes_out_0_3_5;
  wire       [2:0]    subBytes_out_0_3_6;
  wire       [2:0]    subBytes_out_0_3_7;
  wire       [2:0]    subBytes_out_1_0_0;
  wire       [2:0]    subBytes_out_1_0_1;
  wire       [2:0]    subBytes_out_1_0_2;
  wire       [2:0]    subBytes_out_1_0_3;
  wire       [2:0]    subBytes_out_1_0_4;
  wire       [2:0]    subBytes_out_1_0_5;
  wire       [2:0]    subBytes_out_1_0_6;
  wire       [2:0]    subBytes_out_1_0_7;
  wire       [2:0]    subBytes_out_1_1_0;
  wire       [2:0]    subBytes_out_1_1_1;
  wire       [2:0]    subBytes_out_1_1_2;
  wire       [2:0]    subBytes_out_1_1_3;
  wire       [2:0]    subBytes_out_1_1_4;
  wire       [2:0]    subBytes_out_1_1_5;
  wire       [2:0]    subBytes_out_1_1_6;
  wire       [2:0]    subBytes_out_1_1_7;
  wire       [2:0]    subBytes_out_1_2_0;
  wire       [2:0]    subBytes_out_1_2_1;
  wire       [2:0]    subBytes_out_1_2_2;
  wire       [2:0]    subBytes_out_1_2_3;
  wire       [2:0]    subBytes_out_1_2_4;
  wire       [2:0]    subBytes_out_1_2_5;
  wire       [2:0]    subBytes_out_1_2_6;
  wire       [2:0]    subBytes_out_1_2_7;
  wire       [2:0]    subBytes_out_1_3_0;
  wire       [2:0]    subBytes_out_1_3_1;
  wire       [2:0]    subBytes_out_1_3_2;
  wire       [2:0]    subBytes_out_1_3_3;
  wire       [2:0]    subBytes_out_1_3_4;
  wire       [2:0]    subBytes_out_1_3_5;
  wire       [2:0]    subBytes_out_1_3_6;
  wire       [2:0]    subBytes_out_1_3_7;
  wire       [2:0]    subBytes_out_2_0_0;
  wire       [2:0]    subBytes_out_2_0_1;
  wire       [2:0]    subBytes_out_2_0_2;
  wire       [2:0]    subBytes_out_2_0_3;
  wire       [2:0]    subBytes_out_2_0_4;
  wire       [2:0]    subBytes_out_2_0_5;
  wire       [2:0]    subBytes_out_2_0_6;
  wire       [2:0]    subBytes_out_2_0_7;
  wire       [2:0]    subBytes_out_2_1_0;
  wire       [2:0]    subBytes_out_2_1_1;
  wire       [2:0]    subBytes_out_2_1_2;
  wire       [2:0]    subBytes_out_2_1_3;
  wire       [2:0]    subBytes_out_2_1_4;
  wire       [2:0]    subBytes_out_2_1_5;
  wire       [2:0]    subBytes_out_2_1_6;
  wire       [2:0]    subBytes_out_2_1_7;
  wire       [2:0]    subBytes_out_2_2_0;
  wire       [2:0]    subBytes_out_2_2_1;
  wire       [2:0]    subBytes_out_2_2_2;
  wire       [2:0]    subBytes_out_2_2_3;
  wire       [2:0]    subBytes_out_2_2_4;
  wire       [2:0]    subBytes_out_2_2_5;
  wire       [2:0]    subBytes_out_2_2_6;
  wire       [2:0]    subBytes_out_2_2_7;
  wire       [2:0]    subBytes_out_2_3_0;
  wire       [2:0]    subBytes_out_2_3_1;
  wire       [2:0]    subBytes_out_2_3_2;
  wire       [2:0]    subBytes_out_2_3_3;
  wire       [2:0]    subBytes_out_2_3_4;
  wire       [2:0]    subBytes_out_2_3_5;
  wire       [2:0]    subBytes_out_2_3_6;
  wire       [2:0]    subBytes_out_2_3_7;
  wire       [2:0]    subBytes_out_3_0_0;
  wire       [2:0]    subBytes_out_3_0_1;
  wire       [2:0]    subBytes_out_3_0_2;
  wire       [2:0]    subBytes_out_3_0_3;
  wire       [2:0]    subBytes_out_3_0_4;
  wire       [2:0]    subBytes_out_3_0_5;
  wire       [2:0]    subBytes_out_3_0_6;
  wire       [2:0]    subBytes_out_3_0_7;
  wire       [2:0]    subBytes_out_3_1_0;
  wire       [2:0]    subBytes_out_3_1_1;
  wire       [2:0]    subBytes_out_3_1_2;
  wire       [2:0]    subBytes_out_3_1_3;
  wire       [2:0]    subBytes_out_3_1_4;
  wire       [2:0]    subBytes_out_3_1_5;
  wire       [2:0]    subBytes_out_3_1_6;
  wire       [2:0]    subBytes_out_3_1_7;
  wire       [2:0]    subBytes_out_3_2_0;
  wire       [2:0]    subBytes_out_3_2_1;
  wire       [2:0]    subBytes_out_3_2_2;
  wire       [2:0]    subBytes_out_3_2_3;
  wire       [2:0]    subBytes_out_3_2_4;
  wire       [2:0]    subBytes_out_3_2_5;
  wire       [2:0]    subBytes_out_3_2_6;
  wire       [2:0]    subBytes_out_3_2_7;
  wire       [2:0]    subBytes_out_3_3_0;
  wire       [2:0]    subBytes_out_3_3_1;
  wire       [2:0]    subBytes_out_3_3_2;
  wire       [2:0]    subBytes_out_3_3_3;
  wire       [2:0]    subBytes_out_3_3_4;
  wire       [2:0]    subBytes_out_3_3_5;
  wire       [2:0]    subBytes_out_3_3_6;
  wire       [2:0]    subBytes_out_3_3_7;
  wire       [2:0]    subBytes_out_4_0_0;
  wire       [2:0]    subBytes_out_4_0_1;
  wire       [2:0]    subBytes_out_4_0_2;
  wire       [2:0]    subBytes_out_4_0_3;
  wire       [2:0]    subBytes_out_4_0_4;
  wire       [2:0]    subBytes_out_4_0_5;
  wire       [2:0]    subBytes_out_4_0_6;
  wire       [2:0]    subBytes_out_4_0_7;
  wire       [2:0]    subBytes_out_4_1_0;
  wire       [2:0]    subBytes_out_4_1_1;
  wire       [2:0]    subBytes_out_4_1_2;
  wire       [2:0]    subBytes_out_4_1_3;
  wire       [2:0]    subBytes_out_4_1_4;
  wire       [2:0]    subBytes_out_4_1_5;
  wire       [2:0]    subBytes_out_4_1_6;
  wire       [2:0]    subBytes_out_4_1_7;
  wire       [2:0]    subBytes_out_4_2_0;
  wire       [2:0]    subBytes_out_4_2_1;
  wire       [2:0]    subBytes_out_4_2_2;
  wire       [2:0]    subBytes_out_4_2_3;
  wire       [2:0]    subBytes_out_4_2_4;
  wire       [2:0]    subBytes_out_4_2_5;
  wire       [2:0]    subBytes_out_4_2_6;
  wire       [2:0]    subBytes_out_4_2_7;
  wire       [2:0]    subBytes_out_4_3_0;
  wire       [2:0]    subBytes_out_4_3_1;
  wire       [2:0]    subBytes_out_4_3_2;
  wire       [2:0]    subBytes_out_4_3_3;
  wire       [2:0]    subBytes_out_4_3_4;
  wire       [2:0]    subBytes_out_4_3_5;
  wire       [2:0]    subBytes_out_4_3_6;
  wire       [2:0]    subBytes_out_4_3_7;
  wire       [2:0]    subBytes_out_5_0_0;
  wire       [2:0]    subBytes_out_5_0_1;
  wire       [2:0]    subBytes_out_5_0_2;
  wire       [2:0]    subBytes_out_5_0_3;
  wire       [2:0]    subBytes_out_5_0_4;
  wire       [2:0]    subBytes_out_5_0_5;
  wire       [2:0]    subBytes_out_5_0_6;
  wire       [2:0]    subBytes_out_5_0_7;
  wire       [2:0]    subBytes_out_5_1_0;
  wire       [2:0]    subBytes_out_5_1_1;
  wire       [2:0]    subBytes_out_5_1_2;
  wire       [2:0]    subBytes_out_5_1_3;
  wire       [2:0]    subBytes_out_5_1_4;
  wire       [2:0]    subBytes_out_5_1_5;
  wire       [2:0]    subBytes_out_5_1_6;
  wire       [2:0]    subBytes_out_5_1_7;
  wire       [2:0]    subBytes_out_5_2_0;
  wire       [2:0]    subBytes_out_5_2_1;
  wire       [2:0]    subBytes_out_5_2_2;
  wire       [2:0]    subBytes_out_5_2_3;
  wire       [2:0]    subBytes_out_5_2_4;
  wire       [2:0]    subBytes_out_5_2_5;
  wire       [2:0]    subBytes_out_5_2_6;
  wire       [2:0]    subBytes_out_5_2_7;
  wire       [2:0]    subBytes_out_5_3_0;
  wire       [2:0]    subBytes_out_5_3_1;
  wire       [2:0]    subBytes_out_5_3_2;
  wire       [2:0]    subBytes_out_5_3_3;
  wire       [2:0]    subBytes_out_5_3_4;
  wire       [2:0]    subBytes_out_5_3_5;
  wire       [2:0]    subBytes_out_5_3_6;
  wire       [2:0]    subBytes_out_5_3_7;
  wire       [2:0]    subBytes_out_6_0_0;
  wire       [2:0]    subBytes_out_6_0_1;
  wire       [2:0]    subBytes_out_6_0_2;
  wire       [2:0]    subBytes_out_6_0_3;
  wire       [2:0]    subBytes_out_6_0_4;
  wire       [2:0]    subBytes_out_6_0_5;
  wire       [2:0]    subBytes_out_6_0_6;
  wire       [2:0]    subBytes_out_6_0_7;
  wire       [2:0]    subBytes_out_6_1_0;
  wire       [2:0]    subBytes_out_6_1_1;
  wire       [2:0]    subBytes_out_6_1_2;
  wire       [2:0]    subBytes_out_6_1_3;
  wire       [2:0]    subBytes_out_6_1_4;
  wire       [2:0]    subBytes_out_6_1_5;
  wire       [2:0]    subBytes_out_6_1_6;
  wire       [2:0]    subBytes_out_6_1_7;
  wire       [2:0]    subBytes_out_6_2_0;
  wire       [2:0]    subBytes_out_6_2_1;
  wire       [2:0]    subBytes_out_6_2_2;
  wire       [2:0]    subBytes_out_6_2_3;
  wire       [2:0]    subBytes_out_6_2_4;
  wire       [2:0]    subBytes_out_6_2_5;
  wire       [2:0]    subBytes_out_6_2_6;
  wire       [2:0]    subBytes_out_6_2_7;
  wire       [2:0]    subBytes_out_6_3_0;
  wire       [2:0]    subBytes_out_6_3_1;
  wire       [2:0]    subBytes_out_6_3_2;
  wire       [2:0]    subBytes_out_6_3_3;
  wire       [2:0]    subBytes_out_6_3_4;
  wire       [2:0]    subBytes_out_6_3_5;
  wire       [2:0]    subBytes_out_6_3_6;
  wire       [2:0]    subBytes_out_6_3_7;
  wire       [2:0]    subBytes_out_7_0_0;
  wire       [2:0]    subBytes_out_7_0_1;
  wire       [2:0]    subBytes_out_7_0_2;
  wire       [2:0]    subBytes_out_7_0_3;
  wire       [2:0]    subBytes_out_7_0_4;
  wire       [2:0]    subBytes_out_7_0_5;
  wire       [2:0]    subBytes_out_7_0_6;
  wire       [2:0]    subBytes_out_7_0_7;
  wire       [2:0]    subBytes_out_7_1_0;
  wire       [2:0]    subBytes_out_7_1_1;
  wire       [2:0]    subBytes_out_7_1_2;
  wire       [2:0]    subBytes_out_7_1_3;
  wire       [2:0]    subBytes_out_7_1_4;
  wire       [2:0]    subBytes_out_7_1_5;
  wire       [2:0]    subBytes_out_7_1_6;
  wire       [2:0]    subBytes_out_7_1_7;
  wire       [2:0]    subBytes_out_7_2_0;
  wire       [2:0]    subBytes_out_7_2_1;
  wire       [2:0]    subBytes_out_7_2_2;
  wire       [2:0]    subBytes_out_7_2_3;
  wire       [2:0]    subBytes_out_7_2_4;
  wire       [2:0]    subBytes_out_7_2_5;
  wire       [2:0]    subBytes_out_7_2_6;
  wire       [2:0]    subBytes_out_7_2_7;
  wire       [2:0]    subBytes_out_7_3_0;
  wire       [2:0]    subBytes_out_7_3_1;
  wire       [2:0]    subBytes_out_7_3_2;
  wire       [2:0]    subBytes_out_7_3_3;
  wire       [2:0]    subBytes_out_7_3_4;
  wire       [2:0]    subBytes_out_7_3_5;
  wire       [2:0]    subBytes_out_7_3_6;
  wire       [2:0]    subBytes_out_7_3_7;
  wire       [2:0]    subBytes_out_8_0_0;
  wire       [2:0]    subBytes_out_8_0_1;
  wire       [2:0]    subBytes_out_8_0_2;
  wire       [2:0]    subBytes_out_8_0_3;
  wire       [2:0]    subBytes_out_8_0_4;
  wire       [2:0]    subBytes_out_8_0_5;
  wire       [2:0]    subBytes_out_8_0_6;
  wire       [2:0]    subBytes_out_8_0_7;
  wire       [2:0]    subBytes_out_8_1_0;
  wire       [2:0]    subBytes_out_8_1_1;
  wire       [2:0]    subBytes_out_8_1_2;
  wire       [2:0]    subBytes_out_8_1_3;
  wire       [2:0]    subBytes_out_8_1_4;
  wire       [2:0]    subBytes_out_8_1_5;
  wire       [2:0]    subBytes_out_8_1_6;
  wire       [2:0]    subBytes_out_8_1_7;
  wire       [2:0]    subBytes_out_8_2_0;
  wire       [2:0]    subBytes_out_8_2_1;
  wire       [2:0]    subBytes_out_8_2_2;
  wire       [2:0]    subBytes_out_8_2_3;
  wire       [2:0]    subBytes_out_8_2_4;
  wire       [2:0]    subBytes_out_8_2_5;
  wire       [2:0]    subBytes_out_8_2_6;
  wire       [2:0]    subBytes_out_8_2_7;
  wire       [2:0]    subBytes_out_8_3_0;
  wire       [2:0]    subBytes_out_8_3_1;
  wire       [2:0]    subBytes_out_8_3_2;
  wire       [2:0]    subBytes_out_8_3_3;
  wire       [2:0]    subBytes_out_8_3_4;
  wire       [2:0]    subBytes_out_8_3_5;
  wire       [2:0]    subBytes_out_8_3_6;
  wire       [2:0]    subBytes_out_8_3_7;
  wire       [2:0]    subBytes_out_9_0_0;
  wire       [2:0]    subBytes_out_9_0_1;
  wire       [2:0]    subBytes_out_9_0_2;
  wire       [2:0]    subBytes_out_9_0_3;
  wire       [2:0]    subBytes_out_9_0_4;
  wire       [2:0]    subBytes_out_9_0_5;
  wire       [2:0]    subBytes_out_9_0_6;
  wire       [2:0]    subBytes_out_9_0_7;
  wire       [2:0]    subBytes_out_9_1_0;
  wire       [2:0]    subBytes_out_9_1_1;
  wire       [2:0]    subBytes_out_9_1_2;
  wire       [2:0]    subBytes_out_9_1_3;
  wire       [2:0]    subBytes_out_9_1_4;
  wire       [2:0]    subBytes_out_9_1_5;
  wire       [2:0]    subBytes_out_9_1_6;
  wire       [2:0]    subBytes_out_9_1_7;
  wire       [2:0]    subBytes_out_9_2_0;
  wire       [2:0]    subBytes_out_9_2_1;
  wire       [2:0]    subBytes_out_9_2_2;
  wire       [2:0]    subBytes_out_9_2_3;
  wire       [2:0]    subBytes_out_9_2_4;
  wire       [2:0]    subBytes_out_9_2_5;
  wire       [2:0]    subBytes_out_9_2_6;
  wire       [2:0]    subBytes_out_9_2_7;
  wire       [2:0]    subBytes_out_9_3_0;
  wire       [2:0]    subBytes_out_9_3_1;
  wire       [2:0]    subBytes_out_9_3_2;
  wire       [2:0]    subBytes_out_9_3_3;
  wire       [2:0]    subBytes_out_9_3_4;
  wire       [2:0]    subBytes_out_9_3_5;
  wire       [2:0]    subBytes_out_9_3_6;
  wire       [2:0]    subBytes_out_9_3_7;
  wire       [2:0]    subBytes_out_10_0_0;
  wire       [2:0]    subBytes_out_10_0_1;
  wire       [2:0]    subBytes_out_10_0_2;
  wire       [2:0]    subBytes_out_10_0_3;
  wire       [2:0]    subBytes_out_10_0_4;
  wire       [2:0]    subBytes_out_10_0_5;
  wire       [2:0]    subBytes_out_10_0_6;
  wire       [2:0]    subBytes_out_10_0_7;
  wire       [2:0]    subBytes_out_10_1_0;
  wire       [2:0]    subBytes_out_10_1_1;
  wire       [2:0]    subBytes_out_10_1_2;
  wire       [2:0]    subBytes_out_10_1_3;
  wire       [2:0]    subBytes_out_10_1_4;
  wire       [2:0]    subBytes_out_10_1_5;
  wire       [2:0]    subBytes_out_10_1_6;
  wire       [2:0]    subBytes_out_10_1_7;
  wire       [2:0]    subBytes_out_10_2_0;
  wire       [2:0]    subBytes_out_10_2_1;
  wire       [2:0]    subBytes_out_10_2_2;
  wire       [2:0]    subBytes_out_10_2_3;
  wire       [2:0]    subBytes_out_10_2_4;
  wire       [2:0]    subBytes_out_10_2_5;
  wire       [2:0]    subBytes_out_10_2_6;
  wire       [2:0]    subBytes_out_10_2_7;
  wire       [2:0]    subBytes_out_10_3_0;
  wire       [2:0]    subBytes_out_10_3_1;
  wire       [2:0]    subBytes_out_10_3_2;
  wire       [2:0]    subBytes_out_10_3_3;
  wire       [2:0]    subBytes_out_10_3_4;
  wire       [2:0]    subBytes_out_10_3_5;
  wire       [2:0]    subBytes_out_10_3_6;
  wire       [2:0]    subBytes_out_10_3_7;
  wire       [2:0]    subBytes_out_11_0_0;
  wire       [2:0]    subBytes_out_11_0_1;
  wire       [2:0]    subBytes_out_11_0_2;
  wire       [2:0]    subBytes_out_11_0_3;
  wire       [2:0]    subBytes_out_11_0_4;
  wire       [2:0]    subBytes_out_11_0_5;
  wire       [2:0]    subBytes_out_11_0_6;
  wire       [2:0]    subBytes_out_11_0_7;
  wire       [2:0]    subBytes_out_11_1_0;
  wire       [2:0]    subBytes_out_11_1_1;
  wire       [2:0]    subBytes_out_11_1_2;
  wire       [2:0]    subBytes_out_11_1_3;
  wire       [2:0]    subBytes_out_11_1_4;
  wire       [2:0]    subBytes_out_11_1_5;
  wire       [2:0]    subBytes_out_11_1_6;
  wire       [2:0]    subBytes_out_11_1_7;
  wire       [2:0]    subBytes_out_11_2_0;
  wire       [2:0]    subBytes_out_11_2_1;
  wire       [2:0]    subBytes_out_11_2_2;
  wire       [2:0]    subBytes_out_11_2_3;
  wire       [2:0]    subBytes_out_11_2_4;
  wire       [2:0]    subBytes_out_11_2_5;
  wire       [2:0]    subBytes_out_11_2_6;
  wire       [2:0]    subBytes_out_11_2_7;
  wire       [2:0]    subBytes_out_11_3_0;
  wire       [2:0]    subBytes_out_11_3_1;
  wire       [2:0]    subBytes_out_11_3_2;
  wire       [2:0]    subBytes_out_11_3_3;
  wire       [2:0]    subBytes_out_11_3_4;
  wire       [2:0]    subBytes_out_11_3_5;
  wire       [2:0]    subBytes_out_11_3_6;
  wire       [2:0]    subBytes_out_11_3_7;
  wire       [2:0]    subBytes_out_12_0_0;
  wire       [2:0]    subBytes_out_12_0_1;
  wire       [2:0]    subBytes_out_12_0_2;
  wire       [2:0]    subBytes_out_12_0_3;
  wire       [2:0]    subBytes_out_12_0_4;
  wire       [2:0]    subBytes_out_12_0_5;
  wire       [2:0]    subBytes_out_12_0_6;
  wire       [2:0]    subBytes_out_12_0_7;
  wire       [2:0]    subBytes_out_12_1_0;
  wire       [2:0]    subBytes_out_12_1_1;
  wire       [2:0]    subBytes_out_12_1_2;
  wire       [2:0]    subBytes_out_12_1_3;
  wire       [2:0]    subBytes_out_12_1_4;
  wire       [2:0]    subBytes_out_12_1_5;
  wire       [2:0]    subBytes_out_12_1_6;
  wire       [2:0]    subBytes_out_12_1_7;
  wire       [2:0]    subBytes_out_12_2_0;
  wire       [2:0]    subBytes_out_12_2_1;
  wire       [2:0]    subBytes_out_12_2_2;
  wire       [2:0]    subBytes_out_12_2_3;
  wire       [2:0]    subBytes_out_12_2_4;
  wire       [2:0]    subBytes_out_12_2_5;
  wire       [2:0]    subBytes_out_12_2_6;
  wire       [2:0]    subBytes_out_12_2_7;
  wire       [2:0]    subBytes_out_12_3_0;
  wire       [2:0]    subBytes_out_12_3_1;
  wire       [2:0]    subBytes_out_12_3_2;
  wire       [2:0]    subBytes_out_12_3_3;
  wire       [2:0]    subBytes_out_12_3_4;
  wire       [2:0]    subBytes_out_12_3_5;
  wire       [2:0]    subBytes_out_12_3_6;
  wire       [2:0]    subBytes_out_12_3_7;
  wire       [2:0]    subBytes_out_13_0_0;
  wire       [2:0]    subBytes_out_13_0_1;
  wire       [2:0]    subBytes_out_13_0_2;
  wire       [2:0]    subBytes_out_13_0_3;
  wire       [2:0]    subBytes_out_13_0_4;
  wire       [2:0]    subBytes_out_13_0_5;
  wire       [2:0]    subBytes_out_13_0_6;
  wire       [2:0]    subBytes_out_13_0_7;
  wire       [2:0]    subBytes_out_13_1_0;
  wire       [2:0]    subBytes_out_13_1_1;
  wire       [2:0]    subBytes_out_13_1_2;
  wire       [2:0]    subBytes_out_13_1_3;
  wire       [2:0]    subBytes_out_13_1_4;
  wire       [2:0]    subBytes_out_13_1_5;
  wire       [2:0]    subBytes_out_13_1_6;
  wire       [2:0]    subBytes_out_13_1_7;
  wire       [2:0]    subBytes_out_13_2_0;
  wire       [2:0]    subBytes_out_13_2_1;
  wire       [2:0]    subBytes_out_13_2_2;
  wire       [2:0]    subBytes_out_13_2_3;
  wire       [2:0]    subBytes_out_13_2_4;
  wire       [2:0]    subBytes_out_13_2_5;
  wire       [2:0]    subBytes_out_13_2_6;
  wire       [2:0]    subBytes_out_13_2_7;
  wire       [2:0]    subBytes_out_13_3_0;
  wire       [2:0]    subBytes_out_13_3_1;
  wire       [2:0]    subBytes_out_13_3_2;
  wire       [2:0]    subBytes_out_13_3_3;
  wire       [2:0]    subBytes_out_13_3_4;
  wire       [2:0]    subBytes_out_13_3_5;
  wire       [2:0]    subBytes_out_13_3_6;
  wire       [2:0]    subBytes_out_13_3_7;
  wire       [2:0]    subBytes_out_14_0_0;
  wire       [2:0]    subBytes_out_14_0_1;
  wire       [2:0]    subBytes_out_14_0_2;
  wire       [2:0]    subBytes_out_14_0_3;
  wire       [2:0]    subBytes_out_14_0_4;
  wire       [2:0]    subBytes_out_14_0_5;
  wire       [2:0]    subBytes_out_14_0_6;
  wire       [2:0]    subBytes_out_14_0_7;
  wire       [2:0]    subBytes_out_14_1_0;
  wire       [2:0]    subBytes_out_14_1_1;
  wire       [2:0]    subBytes_out_14_1_2;
  wire       [2:0]    subBytes_out_14_1_3;
  wire       [2:0]    subBytes_out_14_1_4;
  wire       [2:0]    subBytes_out_14_1_5;
  wire       [2:0]    subBytes_out_14_1_6;
  wire       [2:0]    subBytes_out_14_1_7;
  wire       [2:0]    subBytes_out_14_2_0;
  wire       [2:0]    subBytes_out_14_2_1;
  wire       [2:0]    subBytes_out_14_2_2;
  wire       [2:0]    subBytes_out_14_2_3;
  wire       [2:0]    subBytes_out_14_2_4;
  wire       [2:0]    subBytes_out_14_2_5;
  wire       [2:0]    subBytes_out_14_2_6;
  wire       [2:0]    subBytes_out_14_2_7;
  wire       [2:0]    subBytes_out_14_3_0;
  wire       [2:0]    subBytes_out_14_3_1;
  wire       [2:0]    subBytes_out_14_3_2;
  wire       [2:0]    subBytes_out_14_3_3;
  wire       [2:0]    subBytes_out_14_3_4;
  wire       [2:0]    subBytes_out_14_3_5;
  wire       [2:0]    subBytes_out_14_3_6;
  wire       [2:0]    subBytes_out_14_3_7;
  wire       [2:0]    subBytes_out_15_0_0;
  wire       [2:0]    subBytes_out_15_0_1;
  wire       [2:0]    subBytes_out_15_0_2;
  wire       [2:0]    subBytes_out_15_0_3;
  wire       [2:0]    subBytes_out_15_0_4;
  wire       [2:0]    subBytes_out_15_0_5;
  wire       [2:0]    subBytes_out_15_0_6;
  wire       [2:0]    subBytes_out_15_0_7;
  wire       [2:0]    subBytes_out_15_1_0;
  wire       [2:0]    subBytes_out_15_1_1;
  wire       [2:0]    subBytes_out_15_1_2;
  wire       [2:0]    subBytes_out_15_1_3;
  wire       [2:0]    subBytes_out_15_1_4;
  wire       [2:0]    subBytes_out_15_1_5;
  wire       [2:0]    subBytes_out_15_1_6;
  wire       [2:0]    subBytes_out_15_1_7;
  wire       [2:0]    subBytes_out_15_2_0;
  wire       [2:0]    subBytes_out_15_2_1;
  wire       [2:0]    subBytes_out_15_2_2;
  wire       [2:0]    subBytes_out_15_2_3;
  wire       [2:0]    subBytes_out_15_2_4;
  wire       [2:0]    subBytes_out_15_2_5;
  wire       [2:0]    subBytes_out_15_2_6;
  wire       [2:0]    subBytes_out_15_2_7;
  wire       [2:0]    subBytes_out_15_3_0;
  wire       [2:0]    subBytes_out_15_3_1;
  wire       [2:0]    subBytes_out_15_3_2;
  wire       [2:0]    subBytes_out_15_3_3;
  wire       [2:0]    subBytes_out_15_3_4;
  wire       [2:0]    subBytes_out_15_3_5;
  wire       [2:0]    subBytes_out_15_3_6;
  wire       [2:0]    subBytes_out_15_3_7;
  reg        [2:0]    roundReg_0_0_0;
  reg        [2:0]    roundReg_0_0_1;
  reg        [2:0]    roundReg_0_0_2;
  reg        [2:0]    roundReg_0_0_3;
  reg        [2:0]    roundReg_0_0_4;
  reg        [2:0]    roundReg_0_0_5;
  reg        [2:0]    roundReg_0_0_6;
  reg        [2:0]    roundReg_0_0_7;
  reg        [2:0]    roundReg_0_1_0;
  reg        [2:0]    roundReg_0_1_1;
  reg        [2:0]    roundReg_0_1_2;
  reg        [2:0]    roundReg_0_1_3;
  reg        [2:0]    roundReg_0_1_4;
  reg        [2:0]    roundReg_0_1_5;
  reg        [2:0]    roundReg_0_1_6;
  reg        [2:0]    roundReg_0_1_7;
  reg        [2:0]    roundReg_0_2_0;
  reg        [2:0]    roundReg_0_2_1;
  reg        [2:0]    roundReg_0_2_2;
  reg        [2:0]    roundReg_0_2_3;
  reg        [2:0]    roundReg_0_2_4;
  reg        [2:0]    roundReg_0_2_5;
  reg        [2:0]    roundReg_0_2_6;
  reg        [2:0]    roundReg_0_2_7;
  reg        [2:0]    roundReg_0_3_0;
  reg        [2:0]    roundReg_0_3_1;
  reg        [2:0]    roundReg_0_3_2;
  reg        [2:0]    roundReg_0_3_3;
  reg        [2:0]    roundReg_0_3_4;
  reg        [2:0]    roundReg_0_3_5;
  reg        [2:0]    roundReg_0_3_6;
  reg        [2:0]    roundReg_0_3_7;
  reg        [2:0]    roundReg_1_0_0;
  reg        [2:0]    roundReg_1_0_1;
  reg        [2:0]    roundReg_1_0_2;
  reg        [2:0]    roundReg_1_0_3;
  reg        [2:0]    roundReg_1_0_4;
  reg        [2:0]    roundReg_1_0_5;
  reg        [2:0]    roundReg_1_0_6;
  reg        [2:0]    roundReg_1_0_7;
  reg        [2:0]    roundReg_1_1_0;
  reg        [2:0]    roundReg_1_1_1;
  reg        [2:0]    roundReg_1_1_2;
  reg        [2:0]    roundReg_1_1_3;
  reg        [2:0]    roundReg_1_1_4;
  reg        [2:0]    roundReg_1_1_5;
  reg        [2:0]    roundReg_1_1_6;
  reg        [2:0]    roundReg_1_1_7;
  reg        [2:0]    roundReg_1_2_0;
  reg        [2:0]    roundReg_1_2_1;
  reg        [2:0]    roundReg_1_2_2;
  reg        [2:0]    roundReg_1_2_3;
  reg        [2:0]    roundReg_1_2_4;
  reg        [2:0]    roundReg_1_2_5;
  reg        [2:0]    roundReg_1_2_6;
  reg        [2:0]    roundReg_1_2_7;
  reg        [2:0]    roundReg_1_3_0;
  reg        [2:0]    roundReg_1_3_1;
  reg        [2:0]    roundReg_1_3_2;
  reg        [2:0]    roundReg_1_3_3;
  reg        [2:0]    roundReg_1_3_4;
  reg        [2:0]    roundReg_1_3_5;
  reg        [2:0]    roundReg_1_3_6;
  reg        [2:0]    roundReg_1_3_7;
  reg        [2:0]    roundReg_2_0_0;
  reg        [2:0]    roundReg_2_0_1;
  reg        [2:0]    roundReg_2_0_2;
  reg        [2:0]    roundReg_2_0_3;
  reg        [2:0]    roundReg_2_0_4;
  reg        [2:0]    roundReg_2_0_5;
  reg        [2:0]    roundReg_2_0_6;
  reg        [2:0]    roundReg_2_0_7;
  reg        [2:0]    roundReg_2_1_0;
  reg        [2:0]    roundReg_2_1_1;
  reg        [2:0]    roundReg_2_1_2;
  reg        [2:0]    roundReg_2_1_3;
  reg        [2:0]    roundReg_2_1_4;
  reg        [2:0]    roundReg_2_1_5;
  reg        [2:0]    roundReg_2_1_6;
  reg        [2:0]    roundReg_2_1_7;
  reg        [2:0]    roundReg_2_2_0;
  reg        [2:0]    roundReg_2_2_1;
  reg        [2:0]    roundReg_2_2_2;
  reg        [2:0]    roundReg_2_2_3;
  reg        [2:0]    roundReg_2_2_4;
  reg        [2:0]    roundReg_2_2_5;
  reg        [2:0]    roundReg_2_2_6;
  reg        [2:0]    roundReg_2_2_7;
  reg        [2:0]    roundReg_2_3_0;
  reg        [2:0]    roundReg_2_3_1;
  reg        [2:0]    roundReg_2_3_2;
  reg        [2:0]    roundReg_2_3_3;
  reg        [2:0]    roundReg_2_3_4;
  reg        [2:0]    roundReg_2_3_5;
  reg        [2:0]    roundReg_2_3_6;
  reg        [2:0]    roundReg_2_3_7;
  reg        [2:0]    roundReg_3_0_0;
  reg        [2:0]    roundReg_3_0_1;
  reg        [2:0]    roundReg_3_0_2;
  reg        [2:0]    roundReg_3_0_3;
  reg        [2:0]    roundReg_3_0_4;
  reg        [2:0]    roundReg_3_0_5;
  reg        [2:0]    roundReg_3_0_6;
  reg        [2:0]    roundReg_3_0_7;
  reg        [2:0]    roundReg_3_1_0;
  reg        [2:0]    roundReg_3_1_1;
  reg        [2:0]    roundReg_3_1_2;
  reg        [2:0]    roundReg_3_1_3;
  reg        [2:0]    roundReg_3_1_4;
  reg        [2:0]    roundReg_3_1_5;
  reg        [2:0]    roundReg_3_1_6;
  reg        [2:0]    roundReg_3_1_7;
  reg        [2:0]    roundReg_3_2_0;
  reg        [2:0]    roundReg_3_2_1;
  reg        [2:0]    roundReg_3_2_2;
  reg        [2:0]    roundReg_3_2_3;
  reg        [2:0]    roundReg_3_2_4;
  reg        [2:0]    roundReg_3_2_5;
  reg        [2:0]    roundReg_3_2_6;
  reg        [2:0]    roundReg_3_2_7;
  reg        [2:0]    roundReg_3_3_0;
  reg        [2:0]    roundReg_3_3_1;
  reg        [2:0]    roundReg_3_3_2;
  reg        [2:0]    roundReg_3_3_3;
  reg        [2:0]    roundReg_3_3_4;
  reg        [2:0]    roundReg_3_3_5;
  reg        [2:0]    roundReg_3_3_6;
  reg        [2:0]    roundReg_3_3_7;
  reg        [2:0]    roundReg_4_0_0;
  reg        [2:0]    roundReg_4_0_1;
  reg        [2:0]    roundReg_4_0_2;
  reg        [2:0]    roundReg_4_0_3;
  reg        [2:0]    roundReg_4_0_4;
  reg        [2:0]    roundReg_4_0_5;
  reg        [2:0]    roundReg_4_0_6;
  reg        [2:0]    roundReg_4_0_7;
  reg        [2:0]    roundReg_4_1_0;
  reg        [2:0]    roundReg_4_1_1;
  reg        [2:0]    roundReg_4_1_2;
  reg        [2:0]    roundReg_4_1_3;
  reg        [2:0]    roundReg_4_1_4;
  reg        [2:0]    roundReg_4_1_5;
  reg        [2:0]    roundReg_4_1_6;
  reg        [2:0]    roundReg_4_1_7;
  reg        [2:0]    roundReg_4_2_0;
  reg        [2:0]    roundReg_4_2_1;
  reg        [2:0]    roundReg_4_2_2;
  reg        [2:0]    roundReg_4_2_3;
  reg        [2:0]    roundReg_4_2_4;
  reg        [2:0]    roundReg_4_2_5;
  reg        [2:0]    roundReg_4_2_6;
  reg        [2:0]    roundReg_4_2_7;
  reg        [2:0]    roundReg_4_3_0;
  reg        [2:0]    roundReg_4_3_1;
  reg        [2:0]    roundReg_4_3_2;
  reg        [2:0]    roundReg_4_3_3;
  reg        [2:0]    roundReg_4_3_4;
  reg        [2:0]    roundReg_4_3_5;
  reg        [2:0]    roundReg_4_3_6;
  reg        [2:0]    roundReg_4_3_7;
  reg        [2:0]    roundReg_5_0_0;
  reg        [2:0]    roundReg_5_0_1;
  reg        [2:0]    roundReg_5_0_2;
  reg        [2:0]    roundReg_5_0_3;
  reg        [2:0]    roundReg_5_0_4;
  reg        [2:0]    roundReg_5_0_5;
  reg        [2:0]    roundReg_5_0_6;
  reg        [2:0]    roundReg_5_0_7;
  reg        [2:0]    roundReg_5_1_0;
  reg        [2:0]    roundReg_5_1_1;
  reg        [2:0]    roundReg_5_1_2;
  reg        [2:0]    roundReg_5_1_3;
  reg        [2:0]    roundReg_5_1_4;
  reg        [2:0]    roundReg_5_1_5;
  reg        [2:0]    roundReg_5_1_6;
  reg        [2:0]    roundReg_5_1_7;
  reg        [2:0]    roundReg_5_2_0;
  reg        [2:0]    roundReg_5_2_1;
  reg        [2:0]    roundReg_5_2_2;
  reg        [2:0]    roundReg_5_2_3;
  reg        [2:0]    roundReg_5_2_4;
  reg        [2:0]    roundReg_5_2_5;
  reg        [2:0]    roundReg_5_2_6;
  reg        [2:0]    roundReg_5_2_7;
  reg        [2:0]    roundReg_5_3_0;
  reg        [2:0]    roundReg_5_3_1;
  reg        [2:0]    roundReg_5_3_2;
  reg        [2:0]    roundReg_5_3_3;
  reg        [2:0]    roundReg_5_3_4;
  reg        [2:0]    roundReg_5_3_5;
  reg        [2:0]    roundReg_5_3_6;
  reg        [2:0]    roundReg_5_3_7;
  reg        [2:0]    roundReg_6_0_0;
  reg        [2:0]    roundReg_6_0_1;
  reg        [2:0]    roundReg_6_0_2;
  reg        [2:0]    roundReg_6_0_3;
  reg        [2:0]    roundReg_6_0_4;
  reg        [2:0]    roundReg_6_0_5;
  reg        [2:0]    roundReg_6_0_6;
  reg        [2:0]    roundReg_6_0_7;
  reg        [2:0]    roundReg_6_1_0;
  reg        [2:0]    roundReg_6_1_1;
  reg        [2:0]    roundReg_6_1_2;
  reg        [2:0]    roundReg_6_1_3;
  reg        [2:0]    roundReg_6_1_4;
  reg        [2:0]    roundReg_6_1_5;
  reg        [2:0]    roundReg_6_1_6;
  reg        [2:0]    roundReg_6_1_7;
  reg        [2:0]    roundReg_6_2_0;
  reg        [2:0]    roundReg_6_2_1;
  reg        [2:0]    roundReg_6_2_2;
  reg        [2:0]    roundReg_6_2_3;
  reg        [2:0]    roundReg_6_2_4;
  reg        [2:0]    roundReg_6_2_5;
  reg        [2:0]    roundReg_6_2_6;
  reg        [2:0]    roundReg_6_2_7;
  reg        [2:0]    roundReg_6_3_0;
  reg        [2:0]    roundReg_6_3_1;
  reg        [2:0]    roundReg_6_3_2;
  reg        [2:0]    roundReg_6_3_3;
  reg        [2:0]    roundReg_6_3_4;
  reg        [2:0]    roundReg_6_3_5;
  reg        [2:0]    roundReg_6_3_6;
  reg        [2:0]    roundReg_6_3_7;
  reg        [2:0]    roundReg_7_0_0;
  reg        [2:0]    roundReg_7_0_1;
  reg        [2:0]    roundReg_7_0_2;
  reg        [2:0]    roundReg_7_0_3;
  reg        [2:0]    roundReg_7_0_4;
  reg        [2:0]    roundReg_7_0_5;
  reg        [2:0]    roundReg_7_0_6;
  reg        [2:0]    roundReg_7_0_7;
  reg        [2:0]    roundReg_7_1_0;
  reg        [2:0]    roundReg_7_1_1;
  reg        [2:0]    roundReg_7_1_2;
  reg        [2:0]    roundReg_7_1_3;
  reg        [2:0]    roundReg_7_1_4;
  reg        [2:0]    roundReg_7_1_5;
  reg        [2:0]    roundReg_7_1_6;
  reg        [2:0]    roundReg_7_1_7;
  reg        [2:0]    roundReg_7_2_0;
  reg        [2:0]    roundReg_7_2_1;
  reg        [2:0]    roundReg_7_2_2;
  reg        [2:0]    roundReg_7_2_3;
  reg        [2:0]    roundReg_7_2_4;
  reg        [2:0]    roundReg_7_2_5;
  reg        [2:0]    roundReg_7_2_6;
  reg        [2:0]    roundReg_7_2_7;
  reg        [2:0]    roundReg_7_3_0;
  reg        [2:0]    roundReg_7_3_1;
  reg        [2:0]    roundReg_7_3_2;
  reg        [2:0]    roundReg_7_3_3;
  reg        [2:0]    roundReg_7_3_4;
  reg        [2:0]    roundReg_7_3_5;
  reg        [2:0]    roundReg_7_3_6;
  reg        [2:0]    roundReg_7_3_7;
  reg        [2:0]    roundReg_8_0_0;
  reg        [2:0]    roundReg_8_0_1;
  reg        [2:0]    roundReg_8_0_2;
  reg        [2:0]    roundReg_8_0_3;
  reg        [2:0]    roundReg_8_0_4;
  reg        [2:0]    roundReg_8_0_5;
  reg        [2:0]    roundReg_8_0_6;
  reg        [2:0]    roundReg_8_0_7;
  reg        [2:0]    roundReg_8_1_0;
  reg        [2:0]    roundReg_8_1_1;
  reg        [2:0]    roundReg_8_1_2;
  reg        [2:0]    roundReg_8_1_3;
  reg        [2:0]    roundReg_8_1_4;
  reg        [2:0]    roundReg_8_1_5;
  reg        [2:0]    roundReg_8_1_6;
  reg        [2:0]    roundReg_8_1_7;
  reg        [2:0]    roundReg_8_2_0;
  reg        [2:0]    roundReg_8_2_1;
  reg        [2:0]    roundReg_8_2_2;
  reg        [2:0]    roundReg_8_2_3;
  reg        [2:0]    roundReg_8_2_4;
  reg        [2:0]    roundReg_8_2_5;
  reg        [2:0]    roundReg_8_2_6;
  reg        [2:0]    roundReg_8_2_7;
  reg        [2:0]    roundReg_8_3_0;
  reg        [2:0]    roundReg_8_3_1;
  reg        [2:0]    roundReg_8_3_2;
  reg        [2:0]    roundReg_8_3_3;
  reg        [2:0]    roundReg_8_3_4;
  reg        [2:0]    roundReg_8_3_5;
  reg        [2:0]    roundReg_8_3_6;
  reg        [2:0]    roundReg_8_3_7;
  reg        [2:0]    roundReg_9_0_0;
  reg        [2:0]    roundReg_9_0_1;
  reg        [2:0]    roundReg_9_0_2;
  reg        [2:0]    roundReg_9_0_3;
  reg        [2:0]    roundReg_9_0_4;
  reg        [2:0]    roundReg_9_0_5;
  reg        [2:0]    roundReg_9_0_6;
  reg        [2:0]    roundReg_9_0_7;
  reg        [2:0]    roundReg_9_1_0;
  reg        [2:0]    roundReg_9_1_1;
  reg        [2:0]    roundReg_9_1_2;
  reg        [2:0]    roundReg_9_1_3;
  reg        [2:0]    roundReg_9_1_4;
  reg        [2:0]    roundReg_9_1_5;
  reg        [2:0]    roundReg_9_1_6;
  reg        [2:0]    roundReg_9_1_7;
  reg        [2:0]    roundReg_9_2_0;
  reg        [2:0]    roundReg_9_2_1;
  reg        [2:0]    roundReg_9_2_2;
  reg        [2:0]    roundReg_9_2_3;
  reg        [2:0]    roundReg_9_2_4;
  reg        [2:0]    roundReg_9_2_5;
  reg        [2:0]    roundReg_9_2_6;
  reg        [2:0]    roundReg_9_2_7;
  reg        [2:0]    roundReg_9_3_0;
  reg        [2:0]    roundReg_9_3_1;
  reg        [2:0]    roundReg_9_3_2;
  reg        [2:0]    roundReg_9_3_3;
  reg        [2:0]    roundReg_9_3_4;
  reg        [2:0]    roundReg_9_3_5;
  reg        [2:0]    roundReg_9_3_6;
  reg        [2:0]    roundReg_9_3_7;
  reg        [2:0]    roundReg_10_0_0;
  reg        [2:0]    roundReg_10_0_1;
  reg        [2:0]    roundReg_10_0_2;
  reg        [2:0]    roundReg_10_0_3;
  reg        [2:0]    roundReg_10_0_4;
  reg        [2:0]    roundReg_10_0_5;
  reg        [2:0]    roundReg_10_0_6;
  reg        [2:0]    roundReg_10_0_7;
  reg        [2:0]    roundReg_10_1_0;
  reg        [2:0]    roundReg_10_1_1;
  reg        [2:0]    roundReg_10_1_2;
  reg        [2:0]    roundReg_10_1_3;
  reg        [2:0]    roundReg_10_1_4;
  reg        [2:0]    roundReg_10_1_5;
  reg        [2:0]    roundReg_10_1_6;
  reg        [2:0]    roundReg_10_1_7;
  reg        [2:0]    roundReg_10_2_0;
  reg        [2:0]    roundReg_10_2_1;
  reg        [2:0]    roundReg_10_2_2;
  reg        [2:0]    roundReg_10_2_3;
  reg        [2:0]    roundReg_10_2_4;
  reg        [2:0]    roundReg_10_2_5;
  reg        [2:0]    roundReg_10_2_6;
  reg        [2:0]    roundReg_10_2_7;
  reg        [2:0]    roundReg_10_3_0;
  reg        [2:0]    roundReg_10_3_1;
  reg        [2:0]    roundReg_10_3_2;
  reg        [2:0]    roundReg_10_3_3;
  reg        [2:0]    roundReg_10_3_4;
  reg        [2:0]    roundReg_10_3_5;
  reg        [2:0]    roundReg_10_3_6;
  reg        [2:0]    roundReg_10_3_7;
  reg        [2:0]    roundReg_11_0_0;
  reg        [2:0]    roundReg_11_0_1;
  reg        [2:0]    roundReg_11_0_2;
  reg        [2:0]    roundReg_11_0_3;
  reg        [2:0]    roundReg_11_0_4;
  reg        [2:0]    roundReg_11_0_5;
  reg        [2:0]    roundReg_11_0_6;
  reg        [2:0]    roundReg_11_0_7;
  reg        [2:0]    roundReg_11_1_0;
  reg        [2:0]    roundReg_11_1_1;
  reg        [2:0]    roundReg_11_1_2;
  reg        [2:0]    roundReg_11_1_3;
  reg        [2:0]    roundReg_11_1_4;
  reg        [2:0]    roundReg_11_1_5;
  reg        [2:0]    roundReg_11_1_6;
  reg        [2:0]    roundReg_11_1_7;
  reg        [2:0]    roundReg_11_2_0;
  reg        [2:0]    roundReg_11_2_1;
  reg        [2:0]    roundReg_11_2_2;
  reg        [2:0]    roundReg_11_2_3;
  reg        [2:0]    roundReg_11_2_4;
  reg        [2:0]    roundReg_11_2_5;
  reg        [2:0]    roundReg_11_2_6;
  reg        [2:0]    roundReg_11_2_7;
  reg        [2:0]    roundReg_11_3_0;
  reg        [2:0]    roundReg_11_3_1;
  reg        [2:0]    roundReg_11_3_2;
  reg        [2:0]    roundReg_11_3_3;
  reg        [2:0]    roundReg_11_3_4;
  reg        [2:0]    roundReg_11_3_5;
  reg        [2:0]    roundReg_11_3_6;
  reg        [2:0]    roundReg_11_3_7;
  reg        [2:0]    roundReg_12_0_0;
  reg        [2:0]    roundReg_12_0_1;
  reg        [2:0]    roundReg_12_0_2;
  reg        [2:0]    roundReg_12_0_3;
  reg        [2:0]    roundReg_12_0_4;
  reg        [2:0]    roundReg_12_0_5;
  reg        [2:0]    roundReg_12_0_6;
  reg        [2:0]    roundReg_12_0_7;
  reg        [2:0]    roundReg_12_1_0;
  reg        [2:0]    roundReg_12_1_1;
  reg        [2:0]    roundReg_12_1_2;
  reg        [2:0]    roundReg_12_1_3;
  reg        [2:0]    roundReg_12_1_4;
  reg        [2:0]    roundReg_12_1_5;
  reg        [2:0]    roundReg_12_1_6;
  reg        [2:0]    roundReg_12_1_7;
  reg        [2:0]    roundReg_12_2_0;
  reg        [2:0]    roundReg_12_2_1;
  reg        [2:0]    roundReg_12_2_2;
  reg        [2:0]    roundReg_12_2_3;
  reg        [2:0]    roundReg_12_2_4;
  reg        [2:0]    roundReg_12_2_5;
  reg        [2:0]    roundReg_12_2_6;
  reg        [2:0]    roundReg_12_2_7;
  reg        [2:0]    roundReg_12_3_0;
  reg        [2:0]    roundReg_12_3_1;
  reg        [2:0]    roundReg_12_3_2;
  reg        [2:0]    roundReg_12_3_3;
  reg        [2:0]    roundReg_12_3_4;
  reg        [2:0]    roundReg_12_3_5;
  reg        [2:0]    roundReg_12_3_6;
  reg        [2:0]    roundReg_12_3_7;
  reg        [2:0]    roundReg_13_0_0;
  reg        [2:0]    roundReg_13_0_1;
  reg        [2:0]    roundReg_13_0_2;
  reg        [2:0]    roundReg_13_0_3;
  reg        [2:0]    roundReg_13_0_4;
  reg        [2:0]    roundReg_13_0_5;
  reg        [2:0]    roundReg_13_0_6;
  reg        [2:0]    roundReg_13_0_7;
  reg        [2:0]    roundReg_13_1_0;
  reg        [2:0]    roundReg_13_1_1;
  reg        [2:0]    roundReg_13_1_2;
  reg        [2:0]    roundReg_13_1_3;
  reg        [2:0]    roundReg_13_1_4;
  reg        [2:0]    roundReg_13_1_5;
  reg        [2:0]    roundReg_13_1_6;
  reg        [2:0]    roundReg_13_1_7;
  reg        [2:0]    roundReg_13_2_0;
  reg        [2:0]    roundReg_13_2_1;
  reg        [2:0]    roundReg_13_2_2;
  reg        [2:0]    roundReg_13_2_3;
  reg        [2:0]    roundReg_13_2_4;
  reg        [2:0]    roundReg_13_2_5;
  reg        [2:0]    roundReg_13_2_6;
  reg        [2:0]    roundReg_13_2_7;
  reg        [2:0]    roundReg_13_3_0;
  reg        [2:0]    roundReg_13_3_1;
  reg        [2:0]    roundReg_13_3_2;
  reg        [2:0]    roundReg_13_3_3;
  reg        [2:0]    roundReg_13_3_4;
  reg        [2:0]    roundReg_13_3_5;
  reg        [2:0]    roundReg_13_3_6;
  reg        [2:0]    roundReg_13_3_7;
  reg        [2:0]    roundReg_14_0_0;
  reg        [2:0]    roundReg_14_0_1;
  reg        [2:0]    roundReg_14_0_2;
  reg        [2:0]    roundReg_14_0_3;
  reg        [2:0]    roundReg_14_0_4;
  reg        [2:0]    roundReg_14_0_5;
  reg        [2:0]    roundReg_14_0_6;
  reg        [2:0]    roundReg_14_0_7;
  reg        [2:0]    roundReg_14_1_0;
  reg        [2:0]    roundReg_14_1_1;
  reg        [2:0]    roundReg_14_1_2;
  reg        [2:0]    roundReg_14_1_3;
  reg        [2:0]    roundReg_14_1_4;
  reg        [2:0]    roundReg_14_1_5;
  reg        [2:0]    roundReg_14_1_6;
  reg        [2:0]    roundReg_14_1_7;
  reg        [2:0]    roundReg_14_2_0;
  reg        [2:0]    roundReg_14_2_1;
  reg        [2:0]    roundReg_14_2_2;
  reg        [2:0]    roundReg_14_2_3;
  reg        [2:0]    roundReg_14_2_4;
  reg        [2:0]    roundReg_14_2_5;
  reg        [2:0]    roundReg_14_2_6;
  reg        [2:0]    roundReg_14_2_7;
  reg        [2:0]    roundReg_14_3_0;
  reg        [2:0]    roundReg_14_3_1;
  reg        [2:0]    roundReg_14_3_2;
  reg        [2:0]    roundReg_14_3_3;
  reg        [2:0]    roundReg_14_3_4;
  reg        [2:0]    roundReg_14_3_5;
  reg        [2:0]    roundReg_14_3_6;
  reg        [2:0]    roundReg_14_3_7;
  reg        [2:0]    roundReg_15_0_0;
  reg        [2:0]    roundReg_15_0_1;
  reg        [2:0]    roundReg_15_0_2;
  reg        [2:0]    roundReg_15_0_3;
  reg        [2:0]    roundReg_15_0_4;
  reg        [2:0]    roundReg_15_0_5;
  reg        [2:0]    roundReg_15_0_6;
  reg        [2:0]    roundReg_15_0_7;
  reg        [2:0]    roundReg_15_1_0;
  reg        [2:0]    roundReg_15_1_1;
  reg        [2:0]    roundReg_15_1_2;
  reg        [2:0]    roundReg_15_1_3;
  reg        [2:0]    roundReg_15_1_4;
  reg        [2:0]    roundReg_15_1_5;
  reg        [2:0]    roundReg_15_1_6;
  reg        [2:0]    roundReg_15_1_7;
  reg        [2:0]    roundReg_15_2_0;
  reg        [2:0]    roundReg_15_2_1;
  reg        [2:0]    roundReg_15_2_2;
  reg        [2:0]    roundReg_15_2_3;
  reg        [2:0]    roundReg_15_2_4;
  reg        [2:0]    roundReg_15_2_5;
  reg        [2:0]    roundReg_15_2_6;
  reg        [2:0]    roundReg_15_2_7;
  reg        [2:0]    roundReg_15_3_0;
  reg        [2:0]    roundReg_15_3_1;
  reg        [2:0]    roundReg_15_3_2;
  reg        [2:0]    roundReg_15_3_3;
  reg        [2:0]    roundReg_15_3_4;
  reg        [2:0]    roundReg_15_3_5;
  reg        [2:0]    roundReg_15_3_6;
  reg        [2:0]    roundReg_15_3_7;

  AES_KeyAddition keyAdd (
    .port_state_in_0_0_0   (port_state_in_0_0_0[2:0]         ), //i
    .port_state_in_0_0_1   (port_state_in_0_0_1[2:0]         ), //i
    .port_state_in_0_0_2   (port_state_in_0_0_2[2:0]         ), //i
    .port_state_in_0_0_3   (port_state_in_0_0_3[2:0]         ), //i
    .port_state_in_0_0_4   (port_state_in_0_0_4[2:0]         ), //i
    .port_state_in_0_0_5   (port_state_in_0_0_5[2:0]         ), //i
    .port_state_in_0_0_6   (port_state_in_0_0_6[2:0]         ), //i
    .port_state_in_0_0_7   (port_state_in_0_0_7[2:0]         ), //i
    .port_state_in_0_1_0   (port_state_in_0_1_0[2:0]         ), //i
    .port_state_in_0_1_1   (port_state_in_0_1_1[2:0]         ), //i
    .port_state_in_0_1_2   (port_state_in_0_1_2[2:0]         ), //i
    .port_state_in_0_1_3   (port_state_in_0_1_3[2:0]         ), //i
    .port_state_in_0_1_4   (port_state_in_0_1_4[2:0]         ), //i
    .port_state_in_0_1_5   (port_state_in_0_1_5[2:0]         ), //i
    .port_state_in_0_1_6   (port_state_in_0_1_6[2:0]         ), //i
    .port_state_in_0_1_7   (port_state_in_0_1_7[2:0]         ), //i
    .port_state_in_0_2_0   (port_state_in_0_2_0[2:0]         ), //i
    .port_state_in_0_2_1   (port_state_in_0_2_1[2:0]         ), //i
    .port_state_in_0_2_2   (port_state_in_0_2_2[2:0]         ), //i
    .port_state_in_0_2_3   (port_state_in_0_2_3[2:0]         ), //i
    .port_state_in_0_2_4   (port_state_in_0_2_4[2:0]         ), //i
    .port_state_in_0_2_5   (port_state_in_0_2_5[2:0]         ), //i
    .port_state_in_0_2_6   (port_state_in_0_2_6[2:0]         ), //i
    .port_state_in_0_2_7   (port_state_in_0_2_7[2:0]         ), //i
    .port_state_in_0_3_0   (port_state_in_0_3_0[2:0]         ), //i
    .port_state_in_0_3_1   (port_state_in_0_3_1[2:0]         ), //i
    .port_state_in_0_3_2   (port_state_in_0_3_2[2:0]         ), //i
    .port_state_in_0_3_3   (port_state_in_0_3_3[2:0]         ), //i
    .port_state_in_0_3_4   (port_state_in_0_3_4[2:0]         ), //i
    .port_state_in_0_3_5   (port_state_in_0_3_5[2:0]         ), //i
    .port_state_in_0_3_6   (port_state_in_0_3_6[2:0]         ), //i
    .port_state_in_0_3_7   (port_state_in_0_3_7[2:0]         ), //i
    .port_state_in_1_0_0   (port_state_in_1_0_0[2:0]         ), //i
    .port_state_in_1_0_1   (port_state_in_1_0_1[2:0]         ), //i
    .port_state_in_1_0_2   (port_state_in_1_0_2[2:0]         ), //i
    .port_state_in_1_0_3   (port_state_in_1_0_3[2:0]         ), //i
    .port_state_in_1_0_4   (port_state_in_1_0_4[2:0]         ), //i
    .port_state_in_1_0_5   (port_state_in_1_0_5[2:0]         ), //i
    .port_state_in_1_0_6   (port_state_in_1_0_6[2:0]         ), //i
    .port_state_in_1_0_7   (port_state_in_1_0_7[2:0]         ), //i
    .port_state_in_1_1_0   (port_state_in_1_1_0[2:0]         ), //i
    .port_state_in_1_1_1   (port_state_in_1_1_1[2:0]         ), //i
    .port_state_in_1_1_2   (port_state_in_1_1_2[2:0]         ), //i
    .port_state_in_1_1_3   (port_state_in_1_1_3[2:0]         ), //i
    .port_state_in_1_1_4   (port_state_in_1_1_4[2:0]         ), //i
    .port_state_in_1_1_5   (port_state_in_1_1_5[2:0]         ), //i
    .port_state_in_1_1_6   (port_state_in_1_1_6[2:0]         ), //i
    .port_state_in_1_1_7   (port_state_in_1_1_7[2:0]         ), //i
    .port_state_in_1_2_0   (port_state_in_1_2_0[2:0]         ), //i
    .port_state_in_1_2_1   (port_state_in_1_2_1[2:0]         ), //i
    .port_state_in_1_2_2   (port_state_in_1_2_2[2:0]         ), //i
    .port_state_in_1_2_3   (port_state_in_1_2_3[2:0]         ), //i
    .port_state_in_1_2_4   (port_state_in_1_2_4[2:0]         ), //i
    .port_state_in_1_2_5   (port_state_in_1_2_5[2:0]         ), //i
    .port_state_in_1_2_6   (port_state_in_1_2_6[2:0]         ), //i
    .port_state_in_1_2_7   (port_state_in_1_2_7[2:0]         ), //i
    .port_state_in_1_3_0   (port_state_in_1_3_0[2:0]         ), //i
    .port_state_in_1_3_1   (port_state_in_1_3_1[2:0]         ), //i
    .port_state_in_1_3_2   (port_state_in_1_3_2[2:0]         ), //i
    .port_state_in_1_3_3   (port_state_in_1_3_3[2:0]         ), //i
    .port_state_in_1_3_4   (port_state_in_1_3_4[2:0]         ), //i
    .port_state_in_1_3_5   (port_state_in_1_3_5[2:0]         ), //i
    .port_state_in_1_3_6   (port_state_in_1_3_6[2:0]         ), //i
    .port_state_in_1_3_7   (port_state_in_1_3_7[2:0]         ), //i
    .port_state_in_2_0_0   (port_state_in_2_0_0[2:0]         ), //i
    .port_state_in_2_0_1   (port_state_in_2_0_1[2:0]         ), //i
    .port_state_in_2_0_2   (port_state_in_2_0_2[2:0]         ), //i
    .port_state_in_2_0_3   (port_state_in_2_0_3[2:0]         ), //i
    .port_state_in_2_0_4   (port_state_in_2_0_4[2:0]         ), //i
    .port_state_in_2_0_5   (port_state_in_2_0_5[2:0]         ), //i
    .port_state_in_2_0_6   (port_state_in_2_0_6[2:0]         ), //i
    .port_state_in_2_0_7   (port_state_in_2_0_7[2:0]         ), //i
    .port_state_in_2_1_0   (port_state_in_2_1_0[2:0]         ), //i
    .port_state_in_2_1_1   (port_state_in_2_1_1[2:0]         ), //i
    .port_state_in_2_1_2   (port_state_in_2_1_2[2:0]         ), //i
    .port_state_in_2_1_3   (port_state_in_2_1_3[2:0]         ), //i
    .port_state_in_2_1_4   (port_state_in_2_1_4[2:0]         ), //i
    .port_state_in_2_1_5   (port_state_in_2_1_5[2:0]         ), //i
    .port_state_in_2_1_6   (port_state_in_2_1_6[2:0]         ), //i
    .port_state_in_2_1_7   (port_state_in_2_1_7[2:0]         ), //i
    .port_state_in_2_2_0   (port_state_in_2_2_0[2:0]         ), //i
    .port_state_in_2_2_1   (port_state_in_2_2_1[2:0]         ), //i
    .port_state_in_2_2_2   (port_state_in_2_2_2[2:0]         ), //i
    .port_state_in_2_2_3   (port_state_in_2_2_3[2:0]         ), //i
    .port_state_in_2_2_4   (port_state_in_2_2_4[2:0]         ), //i
    .port_state_in_2_2_5   (port_state_in_2_2_5[2:0]         ), //i
    .port_state_in_2_2_6   (port_state_in_2_2_6[2:0]         ), //i
    .port_state_in_2_2_7   (port_state_in_2_2_7[2:0]         ), //i
    .port_state_in_2_3_0   (port_state_in_2_3_0[2:0]         ), //i
    .port_state_in_2_3_1   (port_state_in_2_3_1[2:0]         ), //i
    .port_state_in_2_3_2   (port_state_in_2_3_2[2:0]         ), //i
    .port_state_in_2_3_3   (port_state_in_2_3_3[2:0]         ), //i
    .port_state_in_2_3_4   (port_state_in_2_3_4[2:0]         ), //i
    .port_state_in_2_3_5   (port_state_in_2_3_5[2:0]         ), //i
    .port_state_in_2_3_6   (port_state_in_2_3_6[2:0]         ), //i
    .port_state_in_2_3_7   (port_state_in_2_3_7[2:0]         ), //i
    .port_state_in_3_0_0   (port_state_in_3_0_0[2:0]         ), //i
    .port_state_in_3_0_1   (port_state_in_3_0_1[2:0]         ), //i
    .port_state_in_3_0_2   (port_state_in_3_0_2[2:0]         ), //i
    .port_state_in_3_0_3   (port_state_in_3_0_3[2:0]         ), //i
    .port_state_in_3_0_4   (port_state_in_3_0_4[2:0]         ), //i
    .port_state_in_3_0_5   (port_state_in_3_0_5[2:0]         ), //i
    .port_state_in_3_0_6   (port_state_in_3_0_6[2:0]         ), //i
    .port_state_in_3_0_7   (port_state_in_3_0_7[2:0]         ), //i
    .port_state_in_3_1_0   (port_state_in_3_1_0[2:0]         ), //i
    .port_state_in_3_1_1   (port_state_in_3_1_1[2:0]         ), //i
    .port_state_in_3_1_2   (port_state_in_3_1_2[2:0]         ), //i
    .port_state_in_3_1_3   (port_state_in_3_1_3[2:0]         ), //i
    .port_state_in_3_1_4   (port_state_in_3_1_4[2:0]         ), //i
    .port_state_in_3_1_5   (port_state_in_3_1_5[2:0]         ), //i
    .port_state_in_3_1_6   (port_state_in_3_1_6[2:0]         ), //i
    .port_state_in_3_1_7   (port_state_in_3_1_7[2:0]         ), //i
    .port_state_in_3_2_0   (port_state_in_3_2_0[2:0]         ), //i
    .port_state_in_3_2_1   (port_state_in_3_2_1[2:0]         ), //i
    .port_state_in_3_2_2   (port_state_in_3_2_2[2:0]         ), //i
    .port_state_in_3_2_3   (port_state_in_3_2_3[2:0]         ), //i
    .port_state_in_3_2_4   (port_state_in_3_2_4[2:0]         ), //i
    .port_state_in_3_2_5   (port_state_in_3_2_5[2:0]         ), //i
    .port_state_in_3_2_6   (port_state_in_3_2_6[2:0]         ), //i
    .port_state_in_3_2_7   (port_state_in_3_2_7[2:0]         ), //i
    .port_state_in_3_3_0   (port_state_in_3_3_0[2:0]         ), //i
    .port_state_in_3_3_1   (port_state_in_3_3_1[2:0]         ), //i
    .port_state_in_3_3_2   (port_state_in_3_3_2[2:0]         ), //i
    .port_state_in_3_3_3   (port_state_in_3_3_3[2:0]         ), //i
    .port_state_in_3_3_4   (port_state_in_3_3_4[2:0]         ), //i
    .port_state_in_3_3_5   (port_state_in_3_3_5[2:0]         ), //i
    .port_state_in_3_3_6   (port_state_in_3_3_6[2:0]         ), //i
    .port_state_in_3_3_7   (port_state_in_3_3_7[2:0]         ), //i
    .port_state_in_4_0_0   (port_state_in_4_0_0[2:0]         ), //i
    .port_state_in_4_0_1   (port_state_in_4_0_1[2:0]         ), //i
    .port_state_in_4_0_2   (port_state_in_4_0_2[2:0]         ), //i
    .port_state_in_4_0_3   (port_state_in_4_0_3[2:0]         ), //i
    .port_state_in_4_0_4   (port_state_in_4_0_4[2:0]         ), //i
    .port_state_in_4_0_5   (port_state_in_4_0_5[2:0]         ), //i
    .port_state_in_4_0_6   (port_state_in_4_0_6[2:0]         ), //i
    .port_state_in_4_0_7   (port_state_in_4_0_7[2:0]         ), //i
    .port_state_in_4_1_0   (port_state_in_4_1_0[2:0]         ), //i
    .port_state_in_4_1_1   (port_state_in_4_1_1[2:0]         ), //i
    .port_state_in_4_1_2   (port_state_in_4_1_2[2:0]         ), //i
    .port_state_in_4_1_3   (port_state_in_4_1_3[2:0]         ), //i
    .port_state_in_4_1_4   (port_state_in_4_1_4[2:0]         ), //i
    .port_state_in_4_1_5   (port_state_in_4_1_5[2:0]         ), //i
    .port_state_in_4_1_6   (port_state_in_4_1_6[2:0]         ), //i
    .port_state_in_4_1_7   (port_state_in_4_1_7[2:0]         ), //i
    .port_state_in_4_2_0   (port_state_in_4_2_0[2:0]         ), //i
    .port_state_in_4_2_1   (port_state_in_4_2_1[2:0]         ), //i
    .port_state_in_4_2_2   (port_state_in_4_2_2[2:0]         ), //i
    .port_state_in_4_2_3   (port_state_in_4_2_3[2:0]         ), //i
    .port_state_in_4_2_4   (port_state_in_4_2_4[2:0]         ), //i
    .port_state_in_4_2_5   (port_state_in_4_2_5[2:0]         ), //i
    .port_state_in_4_2_6   (port_state_in_4_2_6[2:0]         ), //i
    .port_state_in_4_2_7   (port_state_in_4_2_7[2:0]         ), //i
    .port_state_in_4_3_0   (port_state_in_4_3_0[2:0]         ), //i
    .port_state_in_4_3_1   (port_state_in_4_3_1[2:0]         ), //i
    .port_state_in_4_3_2   (port_state_in_4_3_2[2:0]         ), //i
    .port_state_in_4_3_3   (port_state_in_4_3_3[2:0]         ), //i
    .port_state_in_4_3_4   (port_state_in_4_3_4[2:0]         ), //i
    .port_state_in_4_3_5   (port_state_in_4_3_5[2:0]         ), //i
    .port_state_in_4_3_6   (port_state_in_4_3_6[2:0]         ), //i
    .port_state_in_4_3_7   (port_state_in_4_3_7[2:0]         ), //i
    .port_state_in_5_0_0   (port_state_in_5_0_0[2:0]         ), //i
    .port_state_in_5_0_1   (port_state_in_5_0_1[2:0]         ), //i
    .port_state_in_5_0_2   (port_state_in_5_0_2[2:0]         ), //i
    .port_state_in_5_0_3   (port_state_in_5_0_3[2:0]         ), //i
    .port_state_in_5_0_4   (port_state_in_5_0_4[2:0]         ), //i
    .port_state_in_5_0_5   (port_state_in_5_0_5[2:0]         ), //i
    .port_state_in_5_0_6   (port_state_in_5_0_6[2:0]         ), //i
    .port_state_in_5_0_7   (port_state_in_5_0_7[2:0]         ), //i
    .port_state_in_5_1_0   (port_state_in_5_1_0[2:0]         ), //i
    .port_state_in_5_1_1   (port_state_in_5_1_1[2:0]         ), //i
    .port_state_in_5_1_2   (port_state_in_5_1_2[2:0]         ), //i
    .port_state_in_5_1_3   (port_state_in_5_1_3[2:0]         ), //i
    .port_state_in_5_1_4   (port_state_in_5_1_4[2:0]         ), //i
    .port_state_in_5_1_5   (port_state_in_5_1_5[2:0]         ), //i
    .port_state_in_5_1_6   (port_state_in_5_1_6[2:0]         ), //i
    .port_state_in_5_1_7   (port_state_in_5_1_7[2:0]         ), //i
    .port_state_in_5_2_0   (port_state_in_5_2_0[2:0]         ), //i
    .port_state_in_5_2_1   (port_state_in_5_2_1[2:0]         ), //i
    .port_state_in_5_2_2   (port_state_in_5_2_2[2:0]         ), //i
    .port_state_in_5_2_3   (port_state_in_5_2_3[2:0]         ), //i
    .port_state_in_5_2_4   (port_state_in_5_2_4[2:0]         ), //i
    .port_state_in_5_2_5   (port_state_in_5_2_5[2:0]         ), //i
    .port_state_in_5_2_6   (port_state_in_5_2_6[2:0]         ), //i
    .port_state_in_5_2_7   (port_state_in_5_2_7[2:0]         ), //i
    .port_state_in_5_3_0   (port_state_in_5_3_0[2:0]         ), //i
    .port_state_in_5_3_1   (port_state_in_5_3_1[2:0]         ), //i
    .port_state_in_5_3_2   (port_state_in_5_3_2[2:0]         ), //i
    .port_state_in_5_3_3   (port_state_in_5_3_3[2:0]         ), //i
    .port_state_in_5_3_4   (port_state_in_5_3_4[2:0]         ), //i
    .port_state_in_5_3_5   (port_state_in_5_3_5[2:0]         ), //i
    .port_state_in_5_3_6   (port_state_in_5_3_6[2:0]         ), //i
    .port_state_in_5_3_7   (port_state_in_5_3_7[2:0]         ), //i
    .port_state_in_6_0_0   (port_state_in_6_0_0[2:0]         ), //i
    .port_state_in_6_0_1   (port_state_in_6_0_1[2:0]         ), //i
    .port_state_in_6_0_2   (port_state_in_6_0_2[2:0]         ), //i
    .port_state_in_6_0_3   (port_state_in_6_0_3[2:0]         ), //i
    .port_state_in_6_0_4   (port_state_in_6_0_4[2:0]         ), //i
    .port_state_in_6_0_5   (port_state_in_6_0_5[2:0]         ), //i
    .port_state_in_6_0_6   (port_state_in_6_0_6[2:0]         ), //i
    .port_state_in_6_0_7   (port_state_in_6_0_7[2:0]         ), //i
    .port_state_in_6_1_0   (port_state_in_6_1_0[2:0]         ), //i
    .port_state_in_6_1_1   (port_state_in_6_1_1[2:0]         ), //i
    .port_state_in_6_1_2   (port_state_in_6_1_2[2:0]         ), //i
    .port_state_in_6_1_3   (port_state_in_6_1_3[2:0]         ), //i
    .port_state_in_6_1_4   (port_state_in_6_1_4[2:0]         ), //i
    .port_state_in_6_1_5   (port_state_in_6_1_5[2:0]         ), //i
    .port_state_in_6_1_6   (port_state_in_6_1_6[2:0]         ), //i
    .port_state_in_6_1_7   (port_state_in_6_1_7[2:0]         ), //i
    .port_state_in_6_2_0   (port_state_in_6_2_0[2:0]         ), //i
    .port_state_in_6_2_1   (port_state_in_6_2_1[2:0]         ), //i
    .port_state_in_6_2_2   (port_state_in_6_2_2[2:0]         ), //i
    .port_state_in_6_2_3   (port_state_in_6_2_3[2:0]         ), //i
    .port_state_in_6_2_4   (port_state_in_6_2_4[2:0]         ), //i
    .port_state_in_6_2_5   (port_state_in_6_2_5[2:0]         ), //i
    .port_state_in_6_2_6   (port_state_in_6_2_6[2:0]         ), //i
    .port_state_in_6_2_7   (port_state_in_6_2_7[2:0]         ), //i
    .port_state_in_6_3_0   (port_state_in_6_3_0[2:0]         ), //i
    .port_state_in_6_3_1   (port_state_in_6_3_1[2:0]         ), //i
    .port_state_in_6_3_2   (port_state_in_6_3_2[2:0]         ), //i
    .port_state_in_6_3_3   (port_state_in_6_3_3[2:0]         ), //i
    .port_state_in_6_3_4   (port_state_in_6_3_4[2:0]         ), //i
    .port_state_in_6_3_5   (port_state_in_6_3_5[2:0]         ), //i
    .port_state_in_6_3_6   (port_state_in_6_3_6[2:0]         ), //i
    .port_state_in_6_3_7   (port_state_in_6_3_7[2:0]         ), //i
    .port_state_in_7_0_0   (port_state_in_7_0_0[2:0]         ), //i
    .port_state_in_7_0_1   (port_state_in_7_0_1[2:0]         ), //i
    .port_state_in_7_0_2   (port_state_in_7_0_2[2:0]         ), //i
    .port_state_in_7_0_3   (port_state_in_7_0_3[2:0]         ), //i
    .port_state_in_7_0_4   (port_state_in_7_0_4[2:0]         ), //i
    .port_state_in_7_0_5   (port_state_in_7_0_5[2:0]         ), //i
    .port_state_in_7_0_6   (port_state_in_7_0_6[2:0]         ), //i
    .port_state_in_7_0_7   (port_state_in_7_0_7[2:0]         ), //i
    .port_state_in_7_1_0   (port_state_in_7_1_0[2:0]         ), //i
    .port_state_in_7_1_1   (port_state_in_7_1_1[2:0]         ), //i
    .port_state_in_7_1_2   (port_state_in_7_1_2[2:0]         ), //i
    .port_state_in_7_1_3   (port_state_in_7_1_3[2:0]         ), //i
    .port_state_in_7_1_4   (port_state_in_7_1_4[2:0]         ), //i
    .port_state_in_7_1_5   (port_state_in_7_1_5[2:0]         ), //i
    .port_state_in_7_1_6   (port_state_in_7_1_6[2:0]         ), //i
    .port_state_in_7_1_7   (port_state_in_7_1_7[2:0]         ), //i
    .port_state_in_7_2_0   (port_state_in_7_2_0[2:0]         ), //i
    .port_state_in_7_2_1   (port_state_in_7_2_1[2:0]         ), //i
    .port_state_in_7_2_2   (port_state_in_7_2_2[2:0]         ), //i
    .port_state_in_7_2_3   (port_state_in_7_2_3[2:0]         ), //i
    .port_state_in_7_2_4   (port_state_in_7_2_4[2:0]         ), //i
    .port_state_in_7_2_5   (port_state_in_7_2_5[2:0]         ), //i
    .port_state_in_7_2_6   (port_state_in_7_2_6[2:0]         ), //i
    .port_state_in_7_2_7   (port_state_in_7_2_7[2:0]         ), //i
    .port_state_in_7_3_0   (port_state_in_7_3_0[2:0]         ), //i
    .port_state_in_7_3_1   (port_state_in_7_3_1[2:0]         ), //i
    .port_state_in_7_3_2   (port_state_in_7_3_2[2:0]         ), //i
    .port_state_in_7_3_3   (port_state_in_7_3_3[2:0]         ), //i
    .port_state_in_7_3_4   (port_state_in_7_3_4[2:0]         ), //i
    .port_state_in_7_3_5   (port_state_in_7_3_5[2:0]         ), //i
    .port_state_in_7_3_6   (port_state_in_7_3_6[2:0]         ), //i
    .port_state_in_7_3_7   (port_state_in_7_3_7[2:0]         ), //i
    .port_state_in_8_0_0   (port_state_in_8_0_0[2:0]         ), //i
    .port_state_in_8_0_1   (port_state_in_8_0_1[2:0]         ), //i
    .port_state_in_8_0_2   (port_state_in_8_0_2[2:0]         ), //i
    .port_state_in_8_0_3   (port_state_in_8_0_3[2:0]         ), //i
    .port_state_in_8_0_4   (port_state_in_8_0_4[2:0]         ), //i
    .port_state_in_8_0_5   (port_state_in_8_0_5[2:0]         ), //i
    .port_state_in_8_0_6   (port_state_in_8_0_6[2:0]         ), //i
    .port_state_in_8_0_7   (port_state_in_8_0_7[2:0]         ), //i
    .port_state_in_8_1_0   (port_state_in_8_1_0[2:0]         ), //i
    .port_state_in_8_1_1   (port_state_in_8_1_1[2:0]         ), //i
    .port_state_in_8_1_2   (port_state_in_8_1_2[2:0]         ), //i
    .port_state_in_8_1_3   (port_state_in_8_1_3[2:0]         ), //i
    .port_state_in_8_1_4   (port_state_in_8_1_4[2:0]         ), //i
    .port_state_in_8_1_5   (port_state_in_8_1_5[2:0]         ), //i
    .port_state_in_8_1_6   (port_state_in_8_1_6[2:0]         ), //i
    .port_state_in_8_1_7   (port_state_in_8_1_7[2:0]         ), //i
    .port_state_in_8_2_0   (port_state_in_8_2_0[2:0]         ), //i
    .port_state_in_8_2_1   (port_state_in_8_2_1[2:0]         ), //i
    .port_state_in_8_2_2   (port_state_in_8_2_2[2:0]         ), //i
    .port_state_in_8_2_3   (port_state_in_8_2_3[2:0]         ), //i
    .port_state_in_8_2_4   (port_state_in_8_2_4[2:0]         ), //i
    .port_state_in_8_2_5   (port_state_in_8_2_5[2:0]         ), //i
    .port_state_in_8_2_6   (port_state_in_8_2_6[2:0]         ), //i
    .port_state_in_8_2_7   (port_state_in_8_2_7[2:0]         ), //i
    .port_state_in_8_3_0   (port_state_in_8_3_0[2:0]         ), //i
    .port_state_in_8_3_1   (port_state_in_8_3_1[2:0]         ), //i
    .port_state_in_8_3_2   (port_state_in_8_3_2[2:0]         ), //i
    .port_state_in_8_3_3   (port_state_in_8_3_3[2:0]         ), //i
    .port_state_in_8_3_4   (port_state_in_8_3_4[2:0]         ), //i
    .port_state_in_8_3_5   (port_state_in_8_3_5[2:0]         ), //i
    .port_state_in_8_3_6   (port_state_in_8_3_6[2:0]         ), //i
    .port_state_in_8_3_7   (port_state_in_8_3_7[2:0]         ), //i
    .port_state_in_9_0_0   (port_state_in_9_0_0[2:0]         ), //i
    .port_state_in_9_0_1   (port_state_in_9_0_1[2:0]         ), //i
    .port_state_in_9_0_2   (port_state_in_9_0_2[2:0]         ), //i
    .port_state_in_9_0_3   (port_state_in_9_0_3[2:0]         ), //i
    .port_state_in_9_0_4   (port_state_in_9_0_4[2:0]         ), //i
    .port_state_in_9_0_5   (port_state_in_9_0_5[2:0]         ), //i
    .port_state_in_9_0_6   (port_state_in_9_0_6[2:0]         ), //i
    .port_state_in_9_0_7   (port_state_in_9_0_7[2:0]         ), //i
    .port_state_in_9_1_0   (port_state_in_9_1_0[2:0]         ), //i
    .port_state_in_9_1_1   (port_state_in_9_1_1[2:0]         ), //i
    .port_state_in_9_1_2   (port_state_in_9_1_2[2:0]         ), //i
    .port_state_in_9_1_3   (port_state_in_9_1_3[2:0]         ), //i
    .port_state_in_9_1_4   (port_state_in_9_1_4[2:0]         ), //i
    .port_state_in_9_1_5   (port_state_in_9_1_5[2:0]         ), //i
    .port_state_in_9_1_6   (port_state_in_9_1_6[2:0]         ), //i
    .port_state_in_9_1_7   (port_state_in_9_1_7[2:0]         ), //i
    .port_state_in_9_2_0   (port_state_in_9_2_0[2:0]         ), //i
    .port_state_in_9_2_1   (port_state_in_9_2_1[2:0]         ), //i
    .port_state_in_9_2_2   (port_state_in_9_2_2[2:0]         ), //i
    .port_state_in_9_2_3   (port_state_in_9_2_3[2:0]         ), //i
    .port_state_in_9_2_4   (port_state_in_9_2_4[2:0]         ), //i
    .port_state_in_9_2_5   (port_state_in_9_2_5[2:0]         ), //i
    .port_state_in_9_2_6   (port_state_in_9_2_6[2:0]         ), //i
    .port_state_in_9_2_7   (port_state_in_9_2_7[2:0]         ), //i
    .port_state_in_9_3_0   (port_state_in_9_3_0[2:0]         ), //i
    .port_state_in_9_3_1   (port_state_in_9_3_1[2:0]         ), //i
    .port_state_in_9_3_2   (port_state_in_9_3_2[2:0]         ), //i
    .port_state_in_9_3_3   (port_state_in_9_3_3[2:0]         ), //i
    .port_state_in_9_3_4   (port_state_in_9_3_4[2:0]         ), //i
    .port_state_in_9_3_5   (port_state_in_9_3_5[2:0]         ), //i
    .port_state_in_9_3_6   (port_state_in_9_3_6[2:0]         ), //i
    .port_state_in_9_3_7   (port_state_in_9_3_7[2:0]         ), //i
    .port_state_in_10_0_0  (port_state_in_10_0_0[2:0]        ), //i
    .port_state_in_10_0_1  (port_state_in_10_0_1[2:0]        ), //i
    .port_state_in_10_0_2  (port_state_in_10_0_2[2:0]        ), //i
    .port_state_in_10_0_3  (port_state_in_10_0_3[2:0]        ), //i
    .port_state_in_10_0_4  (port_state_in_10_0_4[2:0]        ), //i
    .port_state_in_10_0_5  (port_state_in_10_0_5[2:0]        ), //i
    .port_state_in_10_0_6  (port_state_in_10_0_6[2:0]        ), //i
    .port_state_in_10_0_7  (port_state_in_10_0_7[2:0]        ), //i
    .port_state_in_10_1_0  (port_state_in_10_1_0[2:0]        ), //i
    .port_state_in_10_1_1  (port_state_in_10_1_1[2:0]        ), //i
    .port_state_in_10_1_2  (port_state_in_10_1_2[2:0]        ), //i
    .port_state_in_10_1_3  (port_state_in_10_1_3[2:0]        ), //i
    .port_state_in_10_1_4  (port_state_in_10_1_4[2:0]        ), //i
    .port_state_in_10_1_5  (port_state_in_10_1_5[2:0]        ), //i
    .port_state_in_10_1_6  (port_state_in_10_1_6[2:0]        ), //i
    .port_state_in_10_1_7  (port_state_in_10_1_7[2:0]        ), //i
    .port_state_in_10_2_0  (port_state_in_10_2_0[2:0]        ), //i
    .port_state_in_10_2_1  (port_state_in_10_2_1[2:0]        ), //i
    .port_state_in_10_2_2  (port_state_in_10_2_2[2:0]        ), //i
    .port_state_in_10_2_3  (port_state_in_10_2_3[2:0]        ), //i
    .port_state_in_10_2_4  (port_state_in_10_2_4[2:0]        ), //i
    .port_state_in_10_2_5  (port_state_in_10_2_5[2:0]        ), //i
    .port_state_in_10_2_6  (port_state_in_10_2_6[2:0]        ), //i
    .port_state_in_10_2_7  (port_state_in_10_2_7[2:0]        ), //i
    .port_state_in_10_3_0  (port_state_in_10_3_0[2:0]        ), //i
    .port_state_in_10_3_1  (port_state_in_10_3_1[2:0]        ), //i
    .port_state_in_10_3_2  (port_state_in_10_3_2[2:0]        ), //i
    .port_state_in_10_3_3  (port_state_in_10_3_3[2:0]        ), //i
    .port_state_in_10_3_4  (port_state_in_10_3_4[2:0]        ), //i
    .port_state_in_10_3_5  (port_state_in_10_3_5[2:0]        ), //i
    .port_state_in_10_3_6  (port_state_in_10_3_6[2:0]        ), //i
    .port_state_in_10_3_7  (port_state_in_10_3_7[2:0]        ), //i
    .port_state_in_11_0_0  (port_state_in_11_0_0[2:0]        ), //i
    .port_state_in_11_0_1  (port_state_in_11_0_1[2:0]        ), //i
    .port_state_in_11_0_2  (port_state_in_11_0_2[2:0]        ), //i
    .port_state_in_11_0_3  (port_state_in_11_0_3[2:0]        ), //i
    .port_state_in_11_0_4  (port_state_in_11_0_4[2:0]        ), //i
    .port_state_in_11_0_5  (port_state_in_11_0_5[2:0]        ), //i
    .port_state_in_11_0_6  (port_state_in_11_0_6[2:0]        ), //i
    .port_state_in_11_0_7  (port_state_in_11_0_7[2:0]        ), //i
    .port_state_in_11_1_0  (port_state_in_11_1_0[2:0]        ), //i
    .port_state_in_11_1_1  (port_state_in_11_1_1[2:0]        ), //i
    .port_state_in_11_1_2  (port_state_in_11_1_2[2:0]        ), //i
    .port_state_in_11_1_3  (port_state_in_11_1_3[2:0]        ), //i
    .port_state_in_11_1_4  (port_state_in_11_1_4[2:0]        ), //i
    .port_state_in_11_1_5  (port_state_in_11_1_5[2:0]        ), //i
    .port_state_in_11_1_6  (port_state_in_11_1_6[2:0]        ), //i
    .port_state_in_11_1_7  (port_state_in_11_1_7[2:0]        ), //i
    .port_state_in_11_2_0  (port_state_in_11_2_0[2:0]        ), //i
    .port_state_in_11_2_1  (port_state_in_11_2_1[2:0]        ), //i
    .port_state_in_11_2_2  (port_state_in_11_2_2[2:0]        ), //i
    .port_state_in_11_2_3  (port_state_in_11_2_3[2:0]        ), //i
    .port_state_in_11_2_4  (port_state_in_11_2_4[2:0]        ), //i
    .port_state_in_11_2_5  (port_state_in_11_2_5[2:0]        ), //i
    .port_state_in_11_2_6  (port_state_in_11_2_6[2:0]        ), //i
    .port_state_in_11_2_7  (port_state_in_11_2_7[2:0]        ), //i
    .port_state_in_11_3_0  (port_state_in_11_3_0[2:0]        ), //i
    .port_state_in_11_3_1  (port_state_in_11_3_1[2:0]        ), //i
    .port_state_in_11_3_2  (port_state_in_11_3_2[2:0]        ), //i
    .port_state_in_11_3_3  (port_state_in_11_3_3[2:0]        ), //i
    .port_state_in_11_3_4  (port_state_in_11_3_4[2:0]        ), //i
    .port_state_in_11_3_5  (port_state_in_11_3_5[2:0]        ), //i
    .port_state_in_11_3_6  (port_state_in_11_3_6[2:0]        ), //i
    .port_state_in_11_3_7  (port_state_in_11_3_7[2:0]        ), //i
    .port_state_in_12_0_0  (port_state_in_12_0_0[2:0]        ), //i
    .port_state_in_12_0_1  (port_state_in_12_0_1[2:0]        ), //i
    .port_state_in_12_0_2  (port_state_in_12_0_2[2:0]        ), //i
    .port_state_in_12_0_3  (port_state_in_12_0_3[2:0]        ), //i
    .port_state_in_12_0_4  (port_state_in_12_0_4[2:0]        ), //i
    .port_state_in_12_0_5  (port_state_in_12_0_5[2:0]        ), //i
    .port_state_in_12_0_6  (port_state_in_12_0_6[2:0]        ), //i
    .port_state_in_12_0_7  (port_state_in_12_0_7[2:0]        ), //i
    .port_state_in_12_1_0  (port_state_in_12_1_0[2:0]        ), //i
    .port_state_in_12_1_1  (port_state_in_12_1_1[2:0]        ), //i
    .port_state_in_12_1_2  (port_state_in_12_1_2[2:0]        ), //i
    .port_state_in_12_1_3  (port_state_in_12_1_3[2:0]        ), //i
    .port_state_in_12_1_4  (port_state_in_12_1_4[2:0]        ), //i
    .port_state_in_12_1_5  (port_state_in_12_1_5[2:0]        ), //i
    .port_state_in_12_1_6  (port_state_in_12_1_6[2:0]        ), //i
    .port_state_in_12_1_7  (port_state_in_12_1_7[2:0]        ), //i
    .port_state_in_12_2_0  (port_state_in_12_2_0[2:0]        ), //i
    .port_state_in_12_2_1  (port_state_in_12_2_1[2:0]        ), //i
    .port_state_in_12_2_2  (port_state_in_12_2_2[2:0]        ), //i
    .port_state_in_12_2_3  (port_state_in_12_2_3[2:0]        ), //i
    .port_state_in_12_2_4  (port_state_in_12_2_4[2:0]        ), //i
    .port_state_in_12_2_5  (port_state_in_12_2_5[2:0]        ), //i
    .port_state_in_12_2_6  (port_state_in_12_2_6[2:0]        ), //i
    .port_state_in_12_2_7  (port_state_in_12_2_7[2:0]        ), //i
    .port_state_in_12_3_0  (port_state_in_12_3_0[2:0]        ), //i
    .port_state_in_12_3_1  (port_state_in_12_3_1[2:0]        ), //i
    .port_state_in_12_3_2  (port_state_in_12_3_2[2:0]        ), //i
    .port_state_in_12_3_3  (port_state_in_12_3_3[2:0]        ), //i
    .port_state_in_12_3_4  (port_state_in_12_3_4[2:0]        ), //i
    .port_state_in_12_3_5  (port_state_in_12_3_5[2:0]        ), //i
    .port_state_in_12_3_6  (port_state_in_12_3_6[2:0]        ), //i
    .port_state_in_12_3_7  (port_state_in_12_3_7[2:0]        ), //i
    .port_state_in_13_0_0  (port_state_in_13_0_0[2:0]        ), //i
    .port_state_in_13_0_1  (port_state_in_13_0_1[2:0]        ), //i
    .port_state_in_13_0_2  (port_state_in_13_0_2[2:0]        ), //i
    .port_state_in_13_0_3  (port_state_in_13_0_3[2:0]        ), //i
    .port_state_in_13_0_4  (port_state_in_13_0_4[2:0]        ), //i
    .port_state_in_13_0_5  (port_state_in_13_0_5[2:0]        ), //i
    .port_state_in_13_0_6  (port_state_in_13_0_6[2:0]        ), //i
    .port_state_in_13_0_7  (port_state_in_13_0_7[2:0]        ), //i
    .port_state_in_13_1_0  (port_state_in_13_1_0[2:0]        ), //i
    .port_state_in_13_1_1  (port_state_in_13_1_1[2:0]        ), //i
    .port_state_in_13_1_2  (port_state_in_13_1_2[2:0]        ), //i
    .port_state_in_13_1_3  (port_state_in_13_1_3[2:0]        ), //i
    .port_state_in_13_1_4  (port_state_in_13_1_4[2:0]        ), //i
    .port_state_in_13_1_5  (port_state_in_13_1_5[2:0]        ), //i
    .port_state_in_13_1_6  (port_state_in_13_1_6[2:0]        ), //i
    .port_state_in_13_1_7  (port_state_in_13_1_7[2:0]        ), //i
    .port_state_in_13_2_0  (port_state_in_13_2_0[2:0]        ), //i
    .port_state_in_13_2_1  (port_state_in_13_2_1[2:0]        ), //i
    .port_state_in_13_2_2  (port_state_in_13_2_2[2:0]        ), //i
    .port_state_in_13_2_3  (port_state_in_13_2_3[2:0]        ), //i
    .port_state_in_13_2_4  (port_state_in_13_2_4[2:0]        ), //i
    .port_state_in_13_2_5  (port_state_in_13_2_5[2:0]        ), //i
    .port_state_in_13_2_6  (port_state_in_13_2_6[2:0]        ), //i
    .port_state_in_13_2_7  (port_state_in_13_2_7[2:0]        ), //i
    .port_state_in_13_3_0  (port_state_in_13_3_0[2:0]        ), //i
    .port_state_in_13_3_1  (port_state_in_13_3_1[2:0]        ), //i
    .port_state_in_13_3_2  (port_state_in_13_3_2[2:0]        ), //i
    .port_state_in_13_3_3  (port_state_in_13_3_3[2:0]        ), //i
    .port_state_in_13_3_4  (port_state_in_13_3_4[2:0]        ), //i
    .port_state_in_13_3_5  (port_state_in_13_3_5[2:0]        ), //i
    .port_state_in_13_3_6  (port_state_in_13_3_6[2:0]        ), //i
    .port_state_in_13_3_7  (port_state_in_13_3_7[2:0]        ), //i
    .port_state_in_14_0_0  (port_state_in_14_0_0[2:0]        ), //i
    .port_state_in_14_0_1  (port_state_in_14_0_1[2:0]        ), //i
    .port_state_in_14_0_2  (port_state_in_14_0_2[2:0]        ), //i
    .port_state_in_14_0_3  (port_state_in_14_0_3[2:0]        ), //i
    .port_state_in_14_0_4  (port_state_in_14_0_4[2:0]        ), //i
    .port_state_in_14_0_5  (port_state_in_14_0_5[2:0]        ), //i
    .port_state_in_14_0_6  (port_state_in_14_0_6[2:0]        ), //i
    .port_state_in_14_0_7  (port_state_in_14_0_7[2:0]        ), //i
    .port_state_in_14_1_0  (port_state_in_14_1_0[2:0]        ), //i
    .port_state_in_14_1_1  (port_state_in_14_1_1[2:0]        ), //i
    .port_state_in_14_1_2  (port_state_in_14_1_2[2:0]        ), //i
    .port_state_in_14_1_3  (port_state_in_14_1_3[2:0]        ), //i
    .port_state_in_14_1_4  (port_state_in_14_1_4[2:0]        ), //i
    .port_state_in_14_1_5  (port_state_in_14_1_5[2:0]        ), //i
    .port_state_in_14_1_6  (port_state_in_14_1_6[2:0]        ), //i
    .port_state_in_14_1_7  (port_state_in_14_1_7[2:0]        ), //i
    .port_state_in_14_2_0  (port_state_in_14_2_0[2:0]        ), //i
    .port_state_in_14_2_1  (port_state_in_14_2_1[2:0]        ), //i
    .port_state_in_14_2_2  (port_state_in_14_2_2[2:0]        ), //i
    .port_state_in_14_2_3  (port_state_in_14_2_3[2:0]        ), //i
    .port_state_in_14_2_4  (port_state_in_14_2_4[2:0]        ), //i
    .port_state_in_14_2_5  (port_state_in_14_2_5[2:0]        ), //i
    .port_state_in_14_2_6  (port_state_in_14_2_6[2:0]        ), //i
    .port_state_in_14_2_7  (port_state_in_14_2_7[2:0]        ), //i
    .port_state_in_14_3_0  (port_state_in_14_3_0[2:0]        ), //i
    .port_state_in_14_3_1  (port_state_in_14_3_1[2:0]        ), //i
    .port_state_in_14_3_2  (port_state_in_14_3_2[2:0]        ), //i
    .port_state_in_14_3_3  (port_state_in_14_3_3[2:0]        ), //i
    .port_state_in_14_3_4  (port_state_in_14_3_4[2:0]        ), //i
    .port_state_in_14_3_5  (port_state_in_14_3_5[2:0]        ), //i
    .port_state_in_14_3_6  (port_state_in_14_3_6[2:0]        ), //i
    .port_state_in_14_3_7  (port_state_in_14_3_7[2:0]        ), //i
    .port_state_in_15_0_0  (port_state_in_15_0_0[2:0]        ), //i
    .port_state_in_15_0_1  (port_state_in_15_0_1[2:0]        ), //i
    .port_state_in_15_0_2  (port_state_in_15_0_2[2:0]        ), //i
    .port_state_in_15_0_3  (port_state_in_15_0_3[2:0]        ), //i
    .port_state_in_15_0_4  (port_state_in_15_0_4[2:0]        ), //i
    .port_state_in_15_0_5  (port_state_in_15_0_5[2:0]        ), //i
    .port_state_in_15_0_6  (port_state_in_15_0_6[2:0]        ), //i
    .port_state_in_15_0_7  (port_state_in_15_0_7[2:0]        ), //i
    .port_state_in_15_1_0  (port_state_in_15_1_0[2:0]        ), //i
    .port_state_in_15_1_1  (port_state_in_15_1_1[2:0]        ), //i
    .port_state_in_15_1_2  (port_state_in_15_1_2[2:0]        ), //i
    .port_state_in_15_1_3  (port_state_in_15_1_3[2:0]        ), //i
    .port_state_in_15_1_4  (port_state_in_15_1_4[2:0]        ), //i
    .port_state_in_15_1_5  (port_state_in_15_1_5[2:0]        ), //i
    .port_state_in_15_1_6  (port_state_in_15_1_6[2:0]        ), //i
    .port_state_in_15_1_7  (port_state_in_15_1_7[2:0]        ), //i
    .port_state_in_15_2_0  (port_state_in_15_2_0[2:0]        ), //i
    .port_state_in_15_2_1  (port_state_in_15_2_1[2:0]        ), //i
    .port_state_in_15_2_2  (port_state_in_15_2_2[2:0]        ), //i
    .port_state_in_15_2_3  (port_state_in_15_2_3[2:0]        ), //i
    .port_state_in_15_2_4  (port_state_in_15_2_4[2:0]        ), //i
    .port_state_in_15_2_5  (port_state_in_15_2_5[2:0]        ), //i
    .port_state_in_15_2_6  (port_state_in_15_2_6[2:0]        ), //i
    .port_state_in_15_2_7  (port_state_in_15_2_7[2:0]        ), //i
    .port_state_in_15_3_0  (port_state_in_15_3_0[2:0]        ), //i
    .port_state_in_15_3_1  (port_state_in_15_3_1[2:0]        ), //i
    .port_state_in_15_3_2  (port_state_in_15_3_2[2:0]        ), //i
    .port_state_in_15_3_3  (port_state_in_15_3_3[2:0]        ), //i
    .port_state_in_15_3_4  (port_state_in_15_3_4[2:0]        ), //i
    .port_state_in_15_3_5  (port_state_in_15_3_5[2:0]        ), //i
    .port_state_in_15_3_6  (port_state_in_15_3_6[2:0]        ), //i
    .port_state_in_15_3_7  (port_state_in_15_3_7[2:0]        ), //i
    .port_key_0_0_0        (port_key_0_0_0[2:0]              ), //i
    .port_key_0_0_1        (port_key_0_0_1[2:0]              ), //i
    .port_key_0_0_2        (port_key_0_0_2[2:0]              ), //i
    .port_key_0_0_3        (port_key_0_0_3[2:0]              ), //i
    .port_key_0_0_4        (port_key_0_0_4[2:0]              ), //i
    .port_key_0_0_5        (port_key_0_0_5[2:0]              ), //i
    .port_key_0_0_6        (port_key_0_0_6[2:0]              ), //i
    .port_key_0_0_7        (port_key_0_0_7[2:0]              ), //i
    .port_key_0_1_0        (port_key_0_1_0[2:0]              ), //i
    .port_key_0_1_1        (port_key_0_1_1[2:0]              ), //i
    .port_key_0_1_2        (port_key_0_1_2[2:0]              ), //i
    .port_key_0_1_3        (port_key_0_1_3[2:0]              ), //i
    .port_key_0_1_4        (port_key_0_1_4[2:0]              ), //i
    .port_key_0_1_5        (port_key_0_1_5[2:0]              ), //i
    .port_key_0_1_6        (port_key_0_1_6[2:0]              ), //i
    .port_key_0_1_7        (port_key_0_1_7[2:0]              ), //i
    .port_key_0_2_0        (port_key_0_2_0[2:0]              ), //i
    .port_key_0_2_1        (port_key_0_2_1[2:0]              ), //i
    .port_key_0_2_2        (port_key_0_2_2[2:0]              ), //i
    .port_key_0_2_3        (port_key_0_2_3[2:0]              ), //i
    .port_key_0_2_4        (port_key_0_2_4[2:0]              ), //i
    .port_key_0_2_5        (port_key_0_2_5[2:0]              ), //i
    .port_key_0_2_6        (port_key_0_2_6[2:0]              ), //i
    .port_key_0_2_7        (port_key_0_2_7[2:0]              ), //i
    .port_key_0_3_0        (port_key_0_3_0[2:0]              ), //i
    .port_key_0_3_1        (port_key_0_3_1[2:0]              ), //i
    .port_key_0_3_2        (port_key_0_3_2[2:0]              ), //i
    .port_key_0_3_3        (port_key_0_3_3[2:0]              ), //i
    .port_key_0_3_4        (port_key_0_3_4[2:0]              ), //i
    .port_key_0_3_5        (port_key_0_3_5[2:0]              ), //i
    .port_key_0_3_6        (port_key_0_3_6[2:0]              ), //i
    .port_key_0_3_7        (port_key_0_3_7[2:0]              ), //i
    .port_key_1_0_0        (port_key_1_0_0[2:0]              ), //i
    .port_key_1_0_1        (port_key_1_0_1[2:0]              ), //i
    .port_key_1_0_2        (port_key_1_0_2[2:0]              ), //i
    .port_key_1_0_3        (port_key_1_0_3[2:0]              ), //i
    .port_key_1_0_4        (port_key_1_0_4[2:0]              ), //i
    .port_key_1_0_5        (port_key_1_0_5[2:0]              ), //i
    .port_key_1_0_6        (port_key_1_0_6[2:0]              ), //i
    .port_key_1_0_7        (port_key_1_0_7[2:0]              ), //i
    .port_key_1_1_0        (port_key_1_1_0[2:0]              ), //i
    .port_key_1_1_1        (port_key_1_1_1[2:0]              ), //i
    .port_key_1_1_2        (port_key_1_1_2[2:0]              ), //i
    .port_key_1_1_3        (port_key_1_1_3[2:0]              ), //i
    .port_key_1_1_4        (port_key_1_1_4[2:0]              ), //i
    .port_key_1_1_5        (port_key_1_1_5[2:0]              ), //i
    .port_key_1_1_6        (port_key_1_1_6[2:0]              ), //i
    .port_key_1_1_7        (port_key_1_1_7[2:0]              ), //i
    .port_key_1_2_0        (port_key_1_2_0[2:0]              ), //i
    .port_key_1_2_1        (port_key_1_2_1[2:0]              ), //i
    .port_key_1_2_2        (port_key_1_2_2[2:0]              ), //i
    .port_key_1_2_3        (port_key_1_2_3[2:0]              ), //i
    .port_key_1_2_4        (port_key_1_2_4[2:0]              ), //i
    .port_key_1_2_5        (port_key_1_2_5[2:0]              ), //i
    .port_key_1_2_6        (port_key_1_2_6[2:0]              ), //i
    .port_key_1_2_7        (port_key_1_2_7[2:0]              ), //i
    .port_key_1_3_0        (port_key_1_3_0[2:0]              ), //i
    .port_key_1_3_1        (port_key_1_3_1[2:0]              ), //i
    .port_key_1_3_2        (port_key_1_3_2[2:0]              ), //i
    .port_key_1_3_3        (port_key_1_3_3[2:0]              ), //i
    .port_key_1_3_4        (port_key_1_3_4[2:0]              ), //i
    .port_key_1_3_5        (port_key_1_3_5[2:0]              ), //i
    .port_key_1_3_6        (port_key_1_3_6[2:0]              ), //i
    .port_key_1_3_7        (port_key_1_3_7[2:0]              ), //i
    .port_key_2_0_0        (port_key_2_0_0[2:0]              ), //i
    .port_key_2_0_1        (port_key_2_0_1[2:0]              ), //i
    .port_key_2_0_2        (port_key_2_0_2[2:0]              ), //i
    .port_key_2_0_3        (port_key_2_0_3[2:0]              ), //i
    .port_key_2_0_4        (port_key_2_0_4[2:0]              ), //i
    .port_key_2_0_5        (port_key_2_0_5[2:0]              ), //i
    .port_key_2_0_6        (port_key_2_0_6[2:0]              ), //i
    .port_key_2_0_7        (port_key_2_0_7[2:0]              ), //i
    .port_key_2_1_0        (port_key_2_1_0[2:0]              ), //i
    .port_key_2_1_1        (port_key_2_1_1[2:0]              ), //i
    .port_key_2_1_2        (port_key_2_1_2[2:0]              ), //i
    .port_key_2_1_3        (port_key_2_1_3[2:0]              ), //i
    .port_key_2_1_4        (port_key_2_1_4[2:0]              ), //i
    .port_key_2_1_5        (port_key_2_1_5[2:0]              ), //i
    .port_key_2_1_6        (port_key_2_1_6[2:0]              ), //i
    .port_key_2_1_7        (port_key_2_1_7[2:0]              ), //i
    .port_key_2_2_0        (port_key_2_2_0[2:0]              ), //i
    .port_key_2_2_1        (port_key_2_2_1[2:0]              ), //i
    .port_key_2_2_2        (port_key_2_2_2[2:0]              ), //i
    .port_key_2_2_3        (port_key_2_2_3[2:0]              ), //i
    .port_key_2_2_4        (port_key_2_2_4[2:0]              ), //i
    .port_key_2_2_5        (port_key_2_2_5[2:0]              ), //i
    .port_key_2_2_6        (port_key_2_2_6[2:0]              ), //i
    .port_key_2_2_7        (port_key_2_2_7[2:0]              ), //i
    .port_key_2_3_0        (port_key_2_3_0[2:0]              ), //i
    .port_key_2_3_1        (port_key_2_3_1[2:0]              ), //i
    .port_key_2_3_2        (port_key_2_3_2[2:0]              ), //i
    .port_key_2_3_3        (port_key_2_3_3[2:0]              ), //i
    .port_key_2_3_4        (port_key_2_3_4[2:0]              ), //i
    .port_key_2_3_5        (port_key_2_3_5[2:0]              ), //i
    .port_key_2_3_6        (port_key_2_3_6[2:0]              ), //i
    .port_key_2_3_7        (port_key_2_3_7[2:0]              ), //i
    .port_key_3_0_0        (port_key_3_0_0[2:0]              ), //i
    .port_key_3_0_1        (port_key_3_0_1[2:0]              ), //i
    .port_key_3_0_2        (port_key_3_0_2[2:0]              ), //i
    .port_key_3_0_3        (port_key_3_0_3[2:0]              ), //i
    .port_key_3_0_4        (port_key_3_0_4[2:0]              ), //i
    .port_key_3_0_5        (port_key_3_0_5[2:0]              ), //i
    .port_key_3_0_6        (port_key_3_0_6[2:0]              ), //i
    .port_key_3_0_7        (port_key_3_0_7[2:0]              ), //i
    .port_key_3_1_0        (port_key_3_1_0[2:0]              ), //i
    .port_key_3_1_1        (port_key_3_1_1[2:0]              ), //i
    .port_key_3_1_2        (port_key_3_1_2[2:0]              ), //i
    .port_key_3_1_3        (port_key_3_1_3[2:0]              ), //i
    .port_key_3_1_4        (port_key_3_1_4[2:0]              ), //i
    .port_key_3_1_5        (port_key_3_1_5[2:0]              ), //i
    .port_key_3_1_6        (port_key_3_1_6[2:0]              ), //i
    .port_key_3_1_7        (port_key_3_1_7[2:0]              ), //i
    .port_key_3_2_0        (port_key_3_2_0[2:0]              ), //i
    .port_key_3_2_1        (port_key_3_2_1[2:0]              ), //i
    .port_key_3_2_2        (port_key_3_2_2[2:0]              ), //i
    .port_key_3_2_3        (port_key_3_2_3[2:0]              ), //i
    .port_key_3_2_4        (port_key_3_2_4[2:0]              ), //i
    .port_key_3_2_5        (port_key_3_2_5[2:0]              ), //i
    .port_key_3_2_6        (port_key_3_2_6[2:0]              ), //i
    .port_key_3_2_7        (port_key_3_2_7[2:0]              ), //i
    .port_key_3_3_0        (port_key_3_3_0[2:0]              ), //i
    .port_key_3_3_1        (port_key_3_3_1[2:0]              ), //i
    .port_key_3_3_2        (port_key_3_3_2[2:0]              ), //i
    .port_key_3_3_3        (port_key_3_3_3[2:0]              ), //i
    .port_key_3_3_4        (port_key_3_3_4[2:0]              ), //i
    .port_key_3_3_5        (port_key_3_3_5[2:0]              ), //i
    .port_key_3_3_6        (port_key_3_3_6[2:0]              ), //i
    .port_key_3_3_7        (port_key_3_3_7[2:0]              ), //i
    .port_key_4_0_0        (port_key_4_0_0[2:0]              ), //i
    .port_key_4_0_1        (port_key_4_0_1[2:0]              ), //i
    .port_key_4_0_2        (port_key_4_0_2[2:0]              ), //i
    .port_key_4_0_3        (port_key_4_0_3[2:0]              ), //i
    .port_key_4_0_4        (port_key_4_0_4[2:0]              ), //i
    .port_key_4_0_5        (port_key_4_0_5[2:0]              ), //i
    .port_key_4_0_6        (port_key_4_0_6[2:0]              ), //i
    .port_key_4_0_7        (port_key_4_0_7[2:0]              ), //i
    .port_key_4_1_0        (port_key_4_1_0[2:0]              ), //i
    .port_key_4_1_1        (port_key_4_1_1[2:0]              ), //i
    .port_key_4_1_2        (port_key_4_1_2[2:0]              ), //i
    .port_key_4_1_3        (port_key_4_1_3[2:0]              ), //i
    .port_key_4_1_4        (port_key_4_1_4[2:0]              ), //i
    .port_key_4_1_5        (port_key_4_1_5[2:0]              ), //i
    .port_key_4_1_6        (port_key_4_1_6[2:0]              ), //i
    .port_key_4_1_7        (port_key_4_1_7[2:0]              ), //i
    .port_key_4_2_0        (port_key_4_2_0[2:0]              ), //i
    .port_key_4_2_1        (port_key_4_2_1[2:0]              ), //i
    .port_key_4_2_2        (port_key_4_2_2[2:0]              ), //i
    .port_key_4_2_3        (port_key_4_2_3[2:0]              ), //i
    .port_key_4_2_4        (port_key_4_2_4[2:0]              ), //i
    .port_key_4_2_5        (port_key_4_2_5[2:0]              ), //i
    .port_key_4_2_6        (port_key_4_2_6[2:0]              ), //i
    .port_key_4_2_7        (port_key_4_2_7[2:0]              ), //i
    .port_key_4_3_0        (port_key_4_3_0[2:0]              ), //i
    .port_key_4_3_1        (port_key_4_3_1[2:0]              ), //i
    .port_key_4_3_2        (port_key_4_3_2[2:0]              ), //i
    .port_key_4_3_3        (port_key_4_3_3[2:0]              ), //i
    .port_key_4_3_4        (port_key_4_3_4[2:0]              ), //i
    .port_key_4_3_5        (port_key_4_3_5[2:0]              ), //i
    .port_key_4_3_6        (port_key_4_3_6[2:0]              ), //i
    .port_key_4_3_7        (port_key_4_3_7[2:0]              ), //i
    .port_key_5_0_0        (port_key_5_0_0[2:0]              ), //i
    .port_key_5_0_1        (port_key_5_0_1[2:0]              ), //i
    .port_key_5_0_2        (port_key_5_0_2[2:0]              ), //i
    .port_key_5_0_3        (port_key_5_0_3[2:0]              ), //i
    .port_key_5_0_4        (port_key_5_0_4[2:0]              ), //i
    .port_key_5_0_5        (port_key_5_0_5[2:0]              ), //i
    .port_key_5_0_6        (port_key_5_0_6[2:0]              ), //i
    .port_key_5_0_7        (port_key_5_0_7[2:0]              ), //i
    .port_key_5_1_0        (port_key_5_1_0[2:0]              ), //i
    .port_key_5_1_1        (port_key_5_1_1[2:0]              ), //i
    .port_key_5_1_2        (port_key_5_1_2[2:0]              ), //i
    .port_key_5_1_3        (port_key_5_1_3[2:0]              ), //i
    .port_key_5_1_4        (port_key_5_1_4[2:0]              ), //i
    .port_key_5_1_5        (port_key_5_1_5[2:0]              ), //i
    .port_key_5_1_6        (port_key_5_1_6[2:0]              ), //i
    .port_key_5_1_7        (port_key_5_1_7[2:0]              ), //i
    .port_key_5_2_0        (port_key_5_2_0[2:0]              ), //i
    .port_key_5_2_1        (port_key_5_2_1[2:0]              ), //i
    .port_key_5_2_2        (port_key_5_2_2[2:0]              ), //i
    .port_key_5_2_3        (port_key_5_2_3[2:0]              ), //i
    .port_key_5_2_4        (port_key_5_2_4[2:0]              ), //i
    .port_key_5_2_5        (port_key_5_2_5[2:0]              ), //i
    .port_key_5_2_6        (port_key_5_2_6[2:0]              ), //i
    .port_key_5_2_7        (port_key_5_2_7[2:0]              ), //i
    .port_key_5_3_0        (port_key_5_3_0[2:0]              ), //i
    .port_key_5_3_1        (port_key_5_3_1[2:0]              ), //i
    .port_key_5_3_2        (port_key_5_3_2[2:0]              ), //i
    .port_key_5_3_3        (port_key_5_3_3[2:0]              ), //i
    .port_key_5_3_4        (port_key_5_3_4[2:0]              ), //i
    .port_key_5_3_5        (port_key_5_3_5[2:0]              ), //i
    .port_key_5_3_6        (port_key_5_3_6[2:0]              ), //i
    .port_key_5_3_7        (port_key_5_3_7[2:0]              ), //i
    .port_key_6_0_0        (port_key_6_0_0[2:0]              ), //i
    .port_key_6_0_1        (port_key_6_0_1[2:0]              ), //i
    .port_key_6_0_2        (port_key_6_0_2[2:0]              ), //i
    .port_key_6_0_3        (port_key_6_0_3[2:0]              ), //i
    .port_key_6_0_4        (port_key_6_0_4[2:0]              ), //i
    .port_key_6_0_5        (port_key_6_0_5[2:0]              ), //i
    .port_key_6_0_6        (port_key_6_0_6[2:0]              ), //i
    .port_key_6_0_7        (port_key_6_0_7[2:0]              ), //i
    .port_key_6_1_0        (port_key_6_1_0[2:0]              ), //i
    .port_key_6_1_1        (port_key_6_1_1[2:0]              ), //i
    .port_key_6_1_2        (port_key_6_1_2[2:0]              ), //i
    .port_key_6_1_3        (port_key_6_1_3[2:0]              ), //i
    .port_key_6_1_4        (port_key_6_1_4[2:0]              ), //i
    .port_key_6_1_5        (port_key_6_1_5[2:0]              ), //i
    .port_key_6_1_6        (port_key_6_1_6[2:0]              ), //i
    .port_key_6_1_7        (port_key_6_1_7[2:0]              ), //i
    .port_key_6_2_0        (port_key_6_2_0[2:0]              ), //i
    .port_key_6_2_1        (port_key_6_2_1[2:0]              ), //i
    .port_key_6_2_2        (port_key_6_2_2[2:0]              ), //i
    .port_key_6_2_3        (port_key_6_2_3[2:0]              ), //i
    .port_key_6_2_4        (port_key_6_2_4[2:0]              ), //i
    .port_key_6_2_5        (port_key_6_2_5[2:0]              ), //i
    .port_key_6_2_6        (port_key_6_2_6[2:0]              ), //i
    .port_key_6_2_7        (port_key_6_2_7[2:0]              ), //i
    .port_key_6_3_0        (port_key_6_3_0[2:0]              ), //i
    .port_key_6_3_1        (port_key_6_3_1[2:0]              ), //i
    .port_key_6_3_2        (port_key_6_3_2[2:0]              ), //i
    .port_key_6_3_3        (port_key_6_3_3[2:0]              ), //i
    .port_key_6_3_4        (port_key_6_3_4[2:0]              ), //i
    .port_key_6_3_5        (port_key_6_3_5[2:0]              ), //i
    .port_key_6_3_6        (port_key_6_3_6[2:0]              ), //i
    .port_key_6_3_7        (port_key_6_3_7[2:0]              ), //i
    .port_key_7_0_0        (port_key_7_0_0[2:0]              ), //i
    .port_key_7_0_1        (port_key_7_0_1[2:0]              ), //i
    .port_key_7_0_2        (port_key_7_0_2[2:0]              ), //i
    .port_key_7_0_3        (port_key_7_0_3[2:0]              ), //i
    .port_key_7_0_4        (port_key_7_0_4[2:0]              ), //i
    .port_key_7_0_5        (port_key_7_0_5[2:0]              ), //i
    .port_key_7_0_6        (port_key_7_0_6[2:0]              ), //i
    .port_key_7_0_7        (port_key_7_0_7[2:0]              ), //i
    .port_key_7_1_0        (port_key_7_1_0[2:0]              ), //i
    .port_key_7_1_1        (port_key_7_1_1[2:0]              ), //i
    .port_key_7_1_2        (port_key_7_1_2[2:0]              ), //i
    .port_key_7_1_3        (port_key_7_1_3[2:0]              ), //i
    .port_key_7_1_4        (port_key_7_1_4[2:0]              ), //i
    .port_key_7_1_5        (port_key_7_1_5[2:0]              ), //i
    .port_key_7_1_6        (port_key_7_1_6[2:0]              ), //i
    .port_key_7_1_7        (port_key_7_1_7[2:0]              ), //i
    .port_key_7_2_0        (port_key_7_2_0[2:0]              ), //i
    .port_key_7_2_1        (port_key_7_2_1[2:0]              ), //i
    .port_key_7_2_2        (port_key_7_2_2[2:0]              ), //i
    .port_key_7_2_3        (port_key_7_2_3[2:0]              ), //i
    .port_key_7_2_4        (port_key_7_2_4[2:0]              ), //i
    .port_key_7_2_5        (port_key_7_2_5[2:0]              ), //i
    .port_key_7_2_6        (port_key_7_2_6[2:0]              ), //i
    .port_key_7_2_7        (port_key_7_2_7[2:0]              ), //i
    .port_key_7_3_0        (port_key_7_3_0[2:0]              ), //i
    .port_key_7_3_1        (port_key_7_3_1[2:0]              ), //i
    .port_key_7_3_2        (port_key_7_3_2[2:0]              ), //i
    .port_key_7_3_3        (port_key_7_3_3[2:0]              ), //i
    .port_key_7_3_4        (port_key_7_3_4[2:0]              ), //i
    .port_key_7_3_5        (port_key_7_3_5[2:0]              ), //i
    .port_key_7_3_6        (port_key_7_3_6[2:0]              ), //i
    .port_key_7_3_7        (port_key_7_3_7[2:0]              ), //i
    .port_key_8_0_0        (port_key_8_0_0[2:0]              ), //i
    .port_key_8_0_1        (port_key_8_0_1[2:0]              ), //i
    .port_key_8_0_2        (port_key_8_0_2[2:0]              ), //i
    .port_key_8_0_3        (port_key_8_0_3[2:0]              ), //i
    .port_key_8_0_4        (port_key_8_0_4[2:0]              ), //i
    .port_key_8_0_5        (port_key_8_0_5[2:0]              ), //i
    .port_key_8_0_6        (port_key_8_0_6[2:0]              ), //i
    .port_key_8_0_7        (port_key_8_0_7[2:0]              ), //i
    .port_key_8_1_0        (port_key_8_1_0[2:0]              ), //i
    .port_key_8_1_1        (port_key_8_1_1[2:0]              ), //i
    .port_key_8_1_2        (port_key_8_1_2[2:0]              ), //i
    .port_key_8_1_3        (port_key_8_1_3[2:0]              ), //i
    .port_key_8_1_4        (port_key_8_1_4[2:0]              ), //i
    .port_key_8_1_5        (port_key_8_1_5[2:0]              ), //i
    .port_key_8_1_6        (port_key_8_1_6[2:0]              ), //i
    .port_key_8_1_7        (port_key_8_1_7[2:0]              ), //i
    .port_key_8_2_0        (port_key_8_2_0[2:0]              ), //i
    .port_key_8_2_1        (port_key_8_2_1[2:0]              ), //i
    .port_key_8_2_2        (port_key_8_2_2[2:0]              ), //i
    .port_key_8_2_3        (port_key_8_2_3[2:0]              ), //i
    .port_key_8_2_4        (port_key_8_2_4[2:0]              ), //i
    .port_key_8_2_5        (port_key_8_2_5[2:0]              ), //i
    .port_key_8_2_6        (port_key_8_2_6[2:0]              ), //i
    .port_key_8_2_7        (port_key_8_2_7[2:0]              ), //i
    .port_key_8_3_0        (port_key_8_3_0[2:0]              ), //i
    .port_key_8_3_1        (port_key_8_3_1[2:0]              ), //i
    .port_key_8_3_2        (port_key_8_3_2[2:0]              ), //i
    .port_key_8_3_3        (port_key_8_3_3[2:0]              ), //i
    .port_key_8_3_4        (port_key_8_3_4[2:0]              ), //i
    .port_key_8_3_5        (port_key_8_3_5[2:0]              ), //i
    .port_key_8_3_6        (port_key_8_3_6[2:0]              ), //i
    .port_key_8_3_7        (port_key_8_3_7[2:0]              ), //i
    .port_key_9_0_0        (port_key_9_0_0[2:0]              ), //i
    .port_key_9_0_1        (port_key_9_0_1[2:0]              ), //i
    .port_key_9_0_2        (port_key_9_0_2[2:0]              ), //i
    .port_key_9_0_3        (port_key_9_0_3[2:0]              ), //i
    .port_key_9_0_4        (port_key_9_0_4[2:0]              ), //i
    .port_key_9_0_5        (port_key_9_0_5[2:0]              ), //i
    .port_key_9_0_6        (port_key_9_0_6[2:0]              ), //i
    .port_key_9_0_7        (port_key_9_0_7[2:0]              ), //i
    .port_key_9_1_0        (port_key_9_1_0[2:0]              ), //i
    .port_key_9_1_1        (port_key_9_1_1[2:0]              ), //i
    .port_key_9_1_2        (port_key_9_1_2[2:0]              ), //i
    .port_key_9_1_3        (port_key_9_1_3[2:0]              ), //i
    .port_key_9_1_4        (port_key_9_1_4[2:0]              ), //i
    .port_key_9_1_5        (port_key_9_1_5[2:0]              ), //i
    .port_key_9_1_6        (port_key_9_1_6[2:0]              ), //i
    .port_key_9_1_7        (port_key_9_1_7[2:0]              ), //i
    .port_key_9_2_0        (port_key_9_2_0[2:0]              ), //i
    .port_key_9_2_1        (port_key_9_2_1[2:0]              ), //i
    .port_key_9_2_2        (port_key_9_2_2[2:0]              ), //i
    .port_key_9_2_3        (port_key_9_2_3[2:0]              ), //i
    .port_key_9_2_4        (port_key_9_2_4[2:0]              ), //i
    .port_key_9_2_5        (port_key_9_2_5[2:0]              ), //i
    .port_key_9_2_6        (port_key_9_2_6[2:0]              ), //i
    .port_key_9_2_7        (port_key_9_2_7[2:0]              ), //i
    .port_key_9_3_0        (port_key_9_3_0[2:0]              ), //i
    .port_key_9_3_1        (port_key_9_3_1[2:0]              ), //i
    .port_key_9_3_2        (port_key_9_3_2[2:0]              ), //i
    .port_key_9_3_3        (port_key_9_3_3[2:0]              ), //i
    .port_key_9_3_4        (port_key_9_3_4[2:0]              ), //i
    .port_key_9_3_5        (port_key_9_3_5[2:0]              ), //i
    .port_key_9_3_6        (port_key_9_3_6[2:0]              ), //i
    .port_key_9_3_7        (port_key_9_3_7[2:0]              ), //i
    .port_key_10_0_0       (port_key_10_0_0[2:0]             ), //i
    .port_key_10_0_1       (port_key_10_0_1[2:0]             ), //i
    .port_key_10_0_2       (port_key_10_0_2[2:0]             ), //i
    .port_key_10_0_3       (port_key_10_0_3[2:0]             ), //i
    .port_key_10_0_4       (port_key_10_0_4[2:0]             ), //i
    .port_key_10_0_5       (port_key_10_0_5[2:0]             ), //i
    .port_key_10_0_6       (port_key_10_0_6[2:0]             ), //i
    .port_key_10_0_7       (port_key_10_0_7[2:0]             ), //i
    .port_key_10_1_0       (port_key_10_1_0[2:0]             ), //i
    .port_key_10_1_1       (port_key_10_1_1[2:0]             ), //i
    .port_key_10_1_2       (port_key_10_1_2[2:0]             ), //i
    .port_key_10_1_3       (port_key_10_1_3[2:0]             ), //i
    .port_key_10_1_4       (port_key_10_1_4[2:0]             ), //i
    .port_key_10_1_5       (port_key_10_1_5[2:0]             ), //i
    .port_key_10_1_6       (port_key_10_1_6[2:0]             ), //i
    .port_key_10_1_7       (port_key_10_1_7[2:0]             ), //i
    .port_key_10_2_0       (port_key_10_2_0[2:0]             ), //i
    .port_key_10_2_1       (port_key_10_2_1[2:0]             ), //i
    .port_key_10_2_2       (port_key_10_2_2[2:0]             ), //i
    .port_key_10_2_3       (port_key_10_2_3[2:0]             ), //i
    .port_key_10_2_4       (port_key_10_2_4[2:0]             ), //i
    .port_key_10_2_5       (port_key_10_2_5[2:0]             ), //i
    .port_key_10_2_6       (port_key_10_2_6[2:0]             ), //i
    .port_key_10_2_7       (port_key_10_2_7[2:0]             ), //i
    .port_key_10_3_0       (port_key_10_3_0[2:0]             ), //i
    .port_key_10_3_1       (port_key_10_3_1[2:0]             ), //i
    .port_key_10_3_2       (port_key_10_3_2[2:0]             ), //i
    .port_key_10_3_3       (port_key_10_3_3[2:0]             ), //i
    .port_key_10_3_4       (port_key_10_3_4[2:0]             ), //i
    .port_key_10_3_5       (port_key_10_3_5[2:0]             ), //i
    .port_key_10_3_6       (port_key_10_3_6[2:0]             ), //i
    .port_key_10_3_7       (port_key_10_3_7[2:0]             ), //i
    .port_key_11_0_0       (port_key_11_0_0[2:0]             ), //i
    .port_key_11_0_1       (port_key_11_0_1[2:0]             ), //i
    .port_key_11_0_2       (port_key_11_0_2[2:0]             ), //i
    .port_key_11_0_3       (port_key_11_0_3[2:0]             ), //i
    .port_key_11_0_4       (port_key_11_0_4[2:0]             ), //i
    .port_key_11_0_5       (port_key_11_0_5[2:0]             ), //i
    .port_key_11_0_6       (port_key_11_0_6[2:0]             ), //i
    .port_key_11_0_7       (port_key_11_0_7[2:0]             ), //i
    .port_key_11_1_0       (port_key_11_1_0[2:0]             ), //i
    .port_key_11_1_1       (port_key_11_1_1[2:0]             ), //i
    .port_key_11_1_2       (port_key_11_1_2[2:0]             ), //i
    .port_key_11_1_3       (port_key_11_1_3[2:0]             ), //i
    .port_key_11_1_4       (port_key_11_1_4[2:0]             ), //i
    .port_key_11_1_5       (port_key_11_1_5[2:0]             ), //i
    .port_key_11_1_6       (port_key_11_1_6[2:0]             ), //i
    .port_key_11_1_7       (port_key_11_1_7[2:0]             ), //i
    .port_key_11_2_0       (port_key_11_2_0[2:0]             ), //i
    .port_key_11_2_1       (port_key_11_2_1[2:0]             ), //i
    .port_key_11_2_2       (port_key_11_2_2[2:0]             ), //i
    .port_key_11_2_3       (port_key_11_2_3[2:0]             ), //i
    .port_key_11_2_4       (port_key_11_2_4[2:0]             ), //i
    .port_key_11_2_5       (port_key_11_2_5[2:0]             ), //i
    .port_key_11_2_6       (port_key_11_2_6[2:0]             ), //i
    .port_key_11_2_7       (port_key_11_2_7[2:0]             ), //i
    .port_key_11_3_0       (port_key_11_3_0[2:0]             ), //i
    .port_key_11_3_1       (port_key_11_3_1[2:0]             ), //i
    .port_key_11_3_2       (port_key_11_3_2[2:0]             ), //i
    .port_key_11_3_3       (port_key_11_3_3[2:0]             ), //i
    .port_key_11_3_4       (port_key_11_3_4[2:0]             ), //i
    .port_key_11_3_5       (port_key_11_3_5[2:0]             ), //i
    .port_key_11_3_6       (port_key_11_3_6[2:0]             ), //i
    .port_key_11_3_7       (port_key_11_3_7[2:0]             ), //i
    .port_key_12_0_0       (port_key_12_0_0[2:0]             ), //i
    .port_key_12_0_1       (port_key_12_0_1[2:0]             ), //i
    .port_key_12_0_2       (port_key_12_0_2[2:0]             ), //i
    .port_key_12_0_3       (port_key_12_0_3[2:0]             ), //i
    .port_key_12_0_4       (port_key_12_0_4[2:0]             ), //i
    .port_key_12_0_5       (port_key_12_0_5[2:0]             ), //i
    .port_key_12_0_6       (port_key_12_0_6[2:0]             ), //i
    .port_key_12_0_7       (port_key_12_0_7[2:0]             ), //i
    .port_key_12_1_0       (port_key_12_1_0[2:0]             ), //i
    .port_key_12_1_1       (port_key_12_1_1[2:0]             ), //i
    .port_key_12_1_2       (port_key_12_1_2[2:0]             ), //i
    .port_key_12_1_3       (port_key_12_1_3[2:0]             ), //i
    .port_key_12_1_4       (port_key_12_1_4[2:0]             ), //i
    .port_key_12_1_5       (port_key_12_1_5[2:0]             ), //i
    .port_key_12_1_6       (port_key_12_1_6[2:0]             ), //i
    .port_key_12_1_7       (port_key_12_1_7[2:0]             ), //i
    .port_key_12_2_0       (port_key_12_2_0[2:0]             ), //i
    .port_key_12_2_1       (port_key_12_2_1[2:0]             ), //i
    .port_key_12_2_2       (port_key_12_2_2[2:0]             ), //i
    .port_key_12_2_3       (port_key_12_2_3[2:0]             ), //i
    .port_key_12_2_4       (port_key_12_2_4[2:0]             ), //i
    .port_key_12_2_5       (port_key_12_2_5[2:0]             ), //i
    .port_key_12_2_6       (port_key_12_2_6[2:0]             ), //i
    .port_key_12_2_7       (port_key_12_2_7[2:0]             ), //i
    .port_key_12_3_0       (port_key_12_3_0[2:0]             ), //i
    .port_key_12_3_1       (port_key_12_3_1[2:0]             ), //i
    .port_key_12_3_2       (port_key_12_3_2[2:0]             ), //i
    .port_key_12_3_3       (port_key_12_3_3[2:0]             ), //i
    .port_key_12_3_4       (port_key_12_3_4[2:0]             ), //i
    .port_key_12_3_5       (port_key_12_3_5[2:0]             ), //i
    .port_key_12_3_6       (port_key_12_3_6[2:0]             ), //i
    .port_key_12_3_7       (port_key_12_3_7[2:0]             ), //i
    .port_key_13_0_0       (port_key_13_0_0[2:0]             ), //i
    .port_key_13_0_1       (port_key_13_0_1[2:0]             ), //i
    .port_key_13_0_2       (port_key_13_0_2[2:0]             ), //i
    .port_key_13_0_3       (port_key_13_0_3[2:0]             ), //i
    .port_key_13_0_4       (port_key_13_0_4[2:0]             ), //i
    .port_key_13_0_5       (port_key_13_0_5[2:0]             ), //i
    .port_key_13_0_6       (port_key_13_0_6[2:0]             ), //i
    .port_key_13_0_7       (port_key_13_0_7[2:0]             ), //i
    .port_key_13_1_0       (port_key_13_1_0[2:0]             ), //i
    .port_key_13_1_1       (port_key_13_1_1[2:0]             ), //i
    .port_key_13_1_2       (port_key_13_1_2[2:0]             ), //i
    .port_key_13_1_3       (port_key_13_1_3[2:0]             ), //i
    .port_key_13_1_4       (port_key_13_1_4[2:0]             ), //i
    .port_key_13_1_5       (port_key_13_1_5[2:0]             ), //i
    .port_key_13_1_6       (port_key_13_1_6[2:0]             ), //i
    .port_key_13_1_7       (port_key_13_1_7[2:0]             ), //i
    .port_key_13_2_0       (port_key_13_2_0[2:0]             ), //i
    .port_key_13_2_1       (port_key_13_2_1[2:0]             ), //i
    .port_key_13_2_2       (port_key_13_2_2[2:0]             ), //i
    .port_key_13_2_3       (port_key_13_2_3[2:0]             ), //i
    .port_key_13_2_4       (port_key_13_2_4[2:0]             ), //i
    .port_key_13_2_5       (port_key_13_2_5[2:0]             ), //i
    .port_key_13_2_6       (port_key_13_2_6[2:0]             ), //i
    .port_key_13_2_7       (port_key_13_2_7[2:0]             ), //i
    .port_key_13_3_0       (port_key_13_3_0[2:0]             ), //i
    .port_key_13_3_1       (port_key_13_3_1[2:0]             ), //i
    .port_key_13_3_2       (port_key_13_3_2[2:0]             ), //i
    .port_key_13_3_3       (port_key_13_3_3[2:0]             ), //i
    .port_key_13_3_4       (port_key_13_3_4[2:0]             ), //i
    .port_key_13_3_5       (port_key_13_3_5[2:0]             ), //i
    .port_key_13_3_6       (port_key_13_3_6[2:0]             ), //i
    .port_key_13_3_7       (port_key_13_3_7[2:0]             ), //i
    .port_key_14_0_0       (port_key_14_0_0[2:0]             ), //i
    .port_key_14_0_1       (port_key_14_0_1[2:0]             ), //i
    .port_key_14_0_2       (port_key_14_0_2[2:0]             ), //i
    .port_key_14_0_3       (port_key_14_0_3[2:0]             ), //i
    .port_key_14_0_4       (port_key_14_0_4[2:0]             ), //i
    .port_key_14_0_5       (port_key_14_0_5[2:0]             ), //i
    .port_key_14_0_6       (port_key_14_0_6[2:0]             ), //i
    .port_key_14_0_7       (port_key_14_0_7[2:0]             ), //i
    .port_key_14_1_0       (port_key_14_1_0[2:0]             ), //i
    .port_key_14_1_1       (port_key_14_1_1[2:0]             ), //i
    .port_key_14_1_2       (port_key_14_1_2[2:0]             ), //i
    .port_key_14_1_3       (port_key_14_1_3[2:0]             ), //i
    .port_key_14_1_4       (port_key_14_1_4[2:0]             ), //i
    .port_key_14_1_5       (port_key_14_1_5[2:0]             ), //i
    .port_key_14_1_6       (port_key_14_1_6[2:0]             ), //i
    .port_key_14_1_7       (port_key_14_1_7[2:0]             ), //i
    .port_key_14_2_0       (port_key_14_2_0[2:0]             ), //i
    .port_key_14_2_1       (port_key_14_2_1[2:0]             ), //i
    .port_key_14_2_2       (port_key_14_2_2[2:0]             ), //i
    .port_key_14_2_3       (port_key_14_2_3[2:0]             ), //i
    .port_key_14_2_4       (port_key_14_2_4[2:0]             ), //i
    .port_key_14_2_5       (port_key_14_2_5[2:0]             ), //i
    .port_key_14_2_6       (port_key_14_2_6[2:0]             ), //i
    .port_key_14_2_7       (port_key_14_2_7[2:0]             ), //i
    .port_key_14_3_0       (port_key_14_3_0[2:0]             ), //i
    .port_key_14_3_1       (port_key_14_3_1[2:0]             ), //i
    .port_key_14_3_2       (port_key_14_3_2[2:0]             ), //i
    .port_key_14_3_3       (port_key_14_3_3[2:0]             ), //i
    .port_key_14_3_4       (port_key_14_3_4[2:0]             ), //i
    .port_key_14_3_5       (port_key_14_3_5[2:0]             ), //i
    .port_key_14_3_6       (port_key_14_3_6[2:0]             ), //i
    .port_key_14_3_7       (port_key_14_3_7[2:0]             ), //i
    .port_key_15_0_0       (port_key_15_0_0[2:0]             ), //i
    .port_key_15_0_1       (port_key_15_0_1[2:0]             ), //i
    .port_key_15_0_2       (port_key_15_0_2[2:0]             ), //i
    .port_key_15_0_3       (port_key_15_0_3[2:0]             ), //i
    .port_key_15_0_4       (port_key_15_0_4[2:0]             ), //i
    .port_key_15_0_5       (port_key_15_0_5[2:0]             ), //i
    .port_key_15_0_6       (port_key_15_0_6[2:0]             ), //i
    .port_key_15_0_7       (port_key_15_0_7[2:0]             ), //i
    .port_key_15_1_0       (port_key_15_1_0[2:0]             ), //i
    .port_key_15_1_1       (port_key_15_1_1[2:0]             ), //i
    .port_key_15_1_2       (port_key_15_1_2[2:0]             ), //i
    .port_key_15_1_3       (port_key_15_1_3[2:0]             ), //i
    .port_key_15_1_4       (port_key_15_1_4[2:0]             ), //i
    .port_key_15_1_5       (port_key_15_1_5[2:0]             ), //i
    .port_key_15_1_6       (port_key_15_1_6[2:0]             ), //i
    .port_key_15_1_7       (port_key_15_1_7[2:0]             ), //i
    .port_key_15_2_0       (port_key_15_2_0[2:0]             ), //i
    .port_key_15_2_1       (port_key_15_2_1[2:0]             ), //i
    .port_key_15_2_2       (port_key_15_2_2[2:0]             ), //i
    .port_key_15_2_3       (port_key_15_2_3[2:0]             ), //i
    .port_key_15_2_4       (port_key_15_2_4[2:0]             ), //i
    .port_key_15_2_5       (port_key_15_2_5[2:0]             ), //i
    .port_key_15_2_6       (port_key_15_2_6[2:0]             ), //i
    .port_key_15_2_7       (port_key_15_2_7[2:0]             ), //i
    .port_key_15_3_0       (port_key_15_3_0[2:0]             ), //i
    .port_key_15_3_1       (port_key_15_3_1[2:0]             ), //i
    .port_key_15_3_2       (port_key_15_3_2[2:0]             ), //i
    .port_key_15_3_3       (port_key_15_3_3[2:0]             ), //i
    .port_key_15_3_4       (port_key_15_3_4[2:0]             ), //i
    .port_key_15_3_5       (port_key_15_3_5[2:0]             ), //i
    .port_key_15_3_6       (port_key_15_3_6[2:0]             ), //i
    .port_key_15_3_7       (port_key_15_3_7[2:0]             ), //i
    .port_state_out_0_0_0  (keyAdd_port_state_out_0_0_0[2:0] ), //o
    .port_state_out_0_0_1  (keyAdd_port_state_out_0_0_1[2:0] ), //o
    .port_state_out_0_0_2  (keyAdd_port_state_out_0_0_2[2:0] ), //o
    .port_state_out_0_0_3  (keyAdd_port_state_out_0_0_3[2:0] ), //o
    .port_state_out_0_0_4  (keyAdd_port_state_out_0_0_4[2:0] ), //o
    .port_state_out_0_0_5  (keyAdd_port_state_out_0_0_5[2:0] ), //o
    .port_state_out_0_0_6  (keyAdd_port_state_out_0_0_6[2:0] ), //o
    .port_state_out_0_0_7  (keyAdd_port_state_out_0_0_7[2:0] ), //o
    .port_state_out_0_1_0  (keyAdd_port_state_out_0_1_0[2:0] ), //o
    .port_state_out_0_1_1  (keyAdd_port_state_out_0_1_1[2:0] ), //o
    .port_state_out_0_1_2  (keyAdd_port_state_out_0_1_2[2:0] ), //o
    .port_state_out_0_1_3  (keyAdd_port_state_out_0_1_3[2:0] ), //o
    .port_state_out_0_1_4  (keyAdd_port_state_out_0_1_4[2:0] ), //o
    .port_state_out_0_1_5  (keyAdd_port_state_out_0_1_5[2:0] ), //o
    .port_state_out_0_1_6  (keyAdd_port_state_out_0_1_6[2:0] ), //o
    .port_state_out_0_1_7  (keyAdd_port_state_out_0_1_7[2:0] ), //o
    .port_state_out_0_2_0  (keyAdd_port_state_out_0_2_0[2:0] ), //o
    .port_state_out_0_2_1  (keyAdd_port_state_out_0_2_1[2:0] ), //o
    .port_state_out_0_2_2  (keyAdd_port_state_out_0_2_2[2:0] ), //o
    .port_state_out_0_2_3  (keyAdd_port_state_out_0_2_3[2:0] ), //o
    .port_state_out_0_2_4  (keyAdd_port_state_out_0_2_4[2:0] ), //o
    .port_state_out_0_2_5  (keyAdd_port_state_out_0_2_5[2:0] ), //o
    .port_state_out_0_2_6  (keyAdd_port_state_out_0_2_6[2:0] ), //o
    .port_state_out_0_2_7  (keyAdd_port_state_out_0_2_7[2:0] ), //o
    .port_state_out_0_3_0  (keyAdd_port_state_out_0_3_0[2:0] ), //o
    .port_state_out_0_3_1  (keyAdd_port_state_out_0_3_1[2:0] ), //o
    .port_state_out_0_3_2  (keyAdd_port_state_out_0_3_2[2:0] ), //o
    .port_state_out_0_3_3  (keyAdd_port_state_out_0_3_3[2:0] ), //o
    .port_state_out_0_3_4  (keyAdd_port_state_out_0_3_4[2:0] ), //o
    .port_state_out_0_3_5  (keyAdd_port_state_out_0_3_5[2:0] ), //o
    .port_state_out_0_3_6  (keyAdd_port_state_out_0_3_6[2:0] ), //o
    .port_state_out_0_3_7  (keyAdd_port_state_out_0_3_7[2:0] ), //o
    .port_state_out_1_0_0  (keyAdd_port_state_out_1_0_0[2:0] ), //o
    .port_state_out_1_0_1  (keyAdd_port_state_out_1_0_1[2:0] ), //o
    .port_state_out_1_0_2  (keyAdd_port_state_out_1_0_2[2:0] ), //o
    .port_state_out_1_0_3  (keyAdd_port_state_out_1_0_3[2:0] ), //o
    .port_state_out_1_0_4  (keyAdd_port_state_out_1_0_4[2:0] ), //o
    .port_state_out_1_0_5  (keyAdd_port_state_out_1_0_5[2:0] ), //o
    .port_state_out_1_0_6  (keyAdd_port_state_out_1_0_6[2:0] ), //o
    .port_state_out_1_0_7  (keyAdd_port_state_out_1_0_7[2:0] ), //o
    .port_state_out_1_1_0  (keyAdd_port_state_out_1_1_0[2:0] ), //o
    .port_state_out_1_1_1  (keyAdd_port_state_out_1_1_1[2:0] ), //o
    .port_state_out_1_1_2  (keyAdd_port_state_out_1_1_2[2:0] ), //o
    .port_state_out_1_1_3  (keyAdd_port_state_out_1_1_3[2:0] ), //o
    .port_state_out_1_1_4  (keyAdd_port_state_out_1_1_4[2:0] ), //o
    .port_state_out_1_1_5  (keyAdd_port_state_out_1_1_5[2:0] ), //o
    .port_state_out_1_1_6  (keyAdd_port_state_out_1_1_6[2:0] ), //o
    .port_state_out_1_1_7  (keyAdd_port_state_out_1_1_7[2:0] ), //o
    .port_state_out_1_2_0  (keyAdd_port_state_out_1_2_0[2:0] ), //o
    .port_state_out_1_2_1  (keyAdd_port_state_out_1_2_1[2:0] ), //o
    .port_state_out_1_2_2  (keyAdd_port_state_out_1_2_2[2:0] ), //o
    .port_state_out_1_2_3  (keyAdd_port_state_out_1_2_3[2:0] ), //o
    .port_state_out_1_2_4  (keyAdd_port_state_out_1_2_4[2:0] ), //o
    .port_state_out_1_2_5  (keyAdd_port_state_out_1_2_5[2:0] ), //o
    .port_state_out_1_2_6  (keyAdd_port_state_out_1_2_6[2:0] ), //o
    .port_state_out_1_2_7  (keyAdd_port_state_out_1_2_7[2:0] ), //o
    .port_state_out_1_3_0  (keyAdd_port_state_out_1_3_0[2:0] ), //o
    .port_state_out_1_3_1  (keyAdd_port_state_out_1_3_1[2:0] ), //o
    .port_state_out_1_3_2  (keyAdd_port_state_out_1_3_2[2:0] ), //o
    .port_state_out_1_3_3  (keyAdd_port_state_out_1_3_3[2:0] ), //o
    .port_state_out_1_3_4  (keyAdd_port_state_out_1_3_4[2:0] ), //o
    .port_state_out_1_3_5  (keyAdd_port_state_out_1_3_5[2:0] ), //o
    .port_state_out_1_3_6  (keyAdd_port_state_out_1_3_6[2:0] ), //o
    .port_state_out_1_3_7  (keyAdd_port_state_out_1_3_7[2:0] ), //o
    .port_state_out_2_0_0  (keyAdd_port_state_out_2_0_0[2:0] ), //o
    .port_state_out_2_0_1  (keyAdd_port_state_out_2_0_1[2:0] ), //o
    .port_state_out_2_0_2  (keyAdd_port_state_out_2_0_2[2:0] ), //o
    .port_state_out_2_0_3  (keyAdd_port_state_out_2_0_3[2:0] ), //o
    .port_state_out_2_0_4  (keyAdd_port_state_out_2_0_4[2:0] ), //o
    .port_state_out_2_0_5  (keyAdd_port_state_out_2_0_5[2:0] ), //o
    .port_state_out_2_0_6  (keyAdd_port_state_out_2_0_6[2:0] ), //o
    .port_state_out_2_0_7  (keyAdd_port_state_out_2_0_7[2:0] ), //o
    .port_state_out_2_1_0  (keyAdd_port_state_out_2_1_0[2:0] ), //o
    .port_state_out_2_1_1  (keyAdd_port_state_out_2_1_1[2:0] ), //o
    .port_state_out_2_1_2  (keyAdd_port_state_out_2_1_2[2:0] ), //o
    .port_state_out_2_1_3  (keyAdd_port_state_out_2_1_3[2:0] ), //o
    .port_state_out_2_1_4  (keyAdd_port_state_out_2_1_4[2:0] ), //o
    .port_state_out_2_1_5  (keyAdd_port_state_out_2_1_5[2:0] ), //o
    .port_state_out_2_1_6  (keyAdd_port_state_out_2_1_6[2:0] ), //o
    .port_state_out_2_1_7  (keyAdd_port_state_out_2_1_7[2:0] ), //o
    .port_state_out_2_2_0  (keyAdd_port_state_out_2_2_0[2:0] ), //o
    .port_state_out_2_2_1  (keyAdd_port_state_out_2_2_1[2:0] ), //o
    .port_state_out_2_2_2  (keyAdd_port_state_out_2_2_2[2:0] ), //o
    .port_state_out_2_2_3  (keyAdd_port_state_out_2_2_3[2:0] ), //o
    .port_state_out_2_2_4  (keyAdd_port_state_out_2_2_4[2:0] ), //o
    .port_state_out_2_2_5  (keyAdd_port_state_out_2_2_5[2:0] ), //o
    .port_state_out_2_2_6  (keyAdd_port_state_out_2_2_6[2:0] ), //o
    .port_state_out_2_2_7  (keyAdd_port_state_out_2_2_7[2:0] ), //o
    .port_state_out_2_3_0  (keyAdd_port_state_out_2_3_0[2:0] ), //o
    .port_state_out_2_3_1  (keyAdd_port_state_out_2_3_1[2:0] ), //o
    .port_state_out_2_3_2  (keyAdd_port_state_out_2_3_2[2:0] ), //o
    .port_state_out_2_3_3  (keyAdd_port_state_out_2_3_3[2:0] ), //o
    .port_state_out_2_3_4  (keyAdd_port_state_out_2_3_4[2:0] ), //o
    .port_state_out_2_3_5  (keyAdd_port_state_out_2_3_5[2:0] ), //o
    .port_state_out_2_3_6  (keyAdd_port_state_out_2_3_6[2:0] ), //o
    .port_state_out_2_3_7  (keyAdd_port_state_out_2_3_7[2:0] ), //o
    .port_state_out_3_0_0  (keyAdd_port_state_out_3_0_0[2:0] ), //o
    .port_state_out_3_0_1  (keyAdd_port_state_out_3_0_1[2:0] ), //o
    .port_state_out_3_0_2  (keyAdd_port_state_out_3_0_2[2:0] ), //o
    .port_state_out_3_0_3  (keyAdd_port_state_out_3_0_3[2:0] ), //o
    .port_state_out_3_0_4  (keyAdd_port_state_out_3_0_4[2:0] ), //o
    .port_state_out_3_0_5  (keyAdd_port_state_out_3_0_5[2:0] ), //o
    .port_state_out_3_0_6  (keyAdd_port_state_out_3_0_6[2:0] ), //o
    .port_state_out_3_0_7  (keyAdd_port_state_out_3_0_7[2:0] ), //o
    .port_state_out_3_1_0  (keyAdd_port_state_out_3_1_0[2:0] ), //o
    .port_state_out_3_1_1  (keyAdd_port_state_out_3_1_1[2:0] ), //o
    .port_state_out_3_1_2  (keyAdd_port_state_out_3_1_2[2:0] ), //o
    .port_state_out_3_1_3  (keyAdd_port_state_out_3_1_3[2:0] ), //o
    .port_state_out_3_1_4  (keyAdd_port_state_out_3_1_4[2:0] ), //o
    .port_state_out_3_1_5  (keyAdd_port_state_out_3_1_5[2:0] ), //o
    .port_state_out_3_1_6  (keyAdd_port_state_out_3_1_6[2:0] ), //o
    .port_state_out_3_1_7  (keyAdd_port_state_out_3_1_7[2:0] ), //o
    .port_state_out_3_2_0  (keyAdd_port_state_out_3_2_0[2:0] ), //o
    .port_state_out_3_2_1  (keyAdd_port_state_out_3_2_1[2:0] ), //o
    .port_state_out_3_2_2  (keyAdd_port_state_out_3_2_2[2:0] ), //o
    .port_state_out_3_2_3  (keyAdd_port_state_out_3_2_3[2:0] ), //o
    .port_state_out_3_2_4  (keyAdd_port_state_out_3_2_4[2:0] ), //o
    .port_state_out_3_2_5  (keyAdd_port_state_out_3_2_5[2:0] ), //o
    .port_state_out_3_2_6  (keyAdd_port_state_out_3_2_6[2:0] ), //o
    .port_state_out_3_2_7  (keyAdd_port_state_out_3_2_7[2:0] ), //o
    .port_state_out_3_3_0  (keyAdd_port_state_out_3_3_0[2:0] ), //o
    .port_state_out_3_3_1  (keyAdd_port_state_out_3_3_1[2:0] ), //o
    .port_state_out_3_3_2  (keyAdd_port_state_out_3_3_2[2:0] ), //o
    .port_state_out_3_3_3  (keyAdd_port_state_out_3_3_3[2:0] ), //o
    .port_state_out_3_3_4  (keyAdd_port_state_out_3_3_4[2:0] ), //o
    .port_state_out_3_3_5  (keyAdd_port_state_out_3_3_5[2:0] ), //o
    .port_state_out_3_3_6  (keyAdd_port_state_out_3_3_6[2:0] ), //o
    .port_state_out_3_3_7  (keyAdd_port_state_out_3_3_7[2:0] ), //o
    .port_state_out_4_0_0  (keyAdd_port_state_out_4_0_0[2:0] ), //o
    .port_state_out_4_0_1  (keyAdd_port_state_out_4_0_1[2:0] ), //o
    .port_state_out_4_0_2  (keyAdd_port_state_out_4_0_2[2:0] ), //o
    .port_state_out_4_0_3  (keyAdd_port_state_out_4_0_3[2:0] ), //o
    .port_state_out_4_0_4  (keyAdd_port_state_out_4_0_4[2:0] ), //o
    .port_state_out_4_0_5  (keyAdd_port_state_out_4_0_5[2:0] ), //o
    .port_state_out_4_0_6  (keyAdd_port_state_out_4_0_6[2:0] ), //o
    .port_state_out_4_0_7  (keyAdd_port_state_out_4_0_7[2:0] ), //o
    .port_state_out_4_1_0  (keyAdd_port_state_out_4_1_0[2:0] ), //o
    .port_state_out_4_1_1  (keyAdd_port_state_out_4_1_1[2:0] ), //o
    .port_state_out_4_1_2  (keyAdd_port_state_out_4_1_2[2:0] ), //o
    .port_state_out_4_1_3  (keyAdd_port_state_out_4_1_3[2:0] ), //o
    .port_state_out_4_1_4  (keyAdd_port_state_out_4_1_4[2:0] ), //o
    .port_state_out_4_1_5  (keyAdd_port_state_out_4_1_5[2:0] ), //o
    .port_state_out_4_1_6  (keyAdd_port_state_out_4_1_6[2:0] ), //o
    .port_state_out_4_1_7  (keyAdd_port_state_out_4_1_7[2:0] ), //o
    .port_state_out_4_2_0  (keyAdd_port_state_out_4_2_0[2:0] ), //o
    .port_state_out_4_2_1  (keyAdd_port_state_out_4_2_1[2:0] ), //o
    .port_state_out_4_2_2  (keyAdd_port_state_out_4_2_2[2:0] ), //o
    .port_state_out_4_2_3  (keyAdd_port_state_out_4_2_3[2:0] ), //o
    .port_state_out_4_2_4  (keyAdd_port_state_out_4_2_4[2:0] ), //o
    .port_state_out_4_2_5  (keyAdd_port_state_out_4_2_5[2:0] ), //o
    .port_state_out_4_2_6  (keyAdd_port_state_out_4_2_6[2:0] ), //o
    .port_state_out_4_2_7  (keyAdd_port_state_out_4_2_7[2:0] ), //o
    .port_state_out_4_3_0  (keyAdd_port_state_out_4_3_0[2:0] ), //o
    .port_state_out_4_3_1  (keyAdd_port_state_out_4_3_1[2:0] ), //o
    .port_state_out_4_3_2  (keyAdd_port_state_out_4_3_2[2:0] ), //o
    .port_state_out_4_3_3  (keyAdd_port_state_out_4_3_3[2:0] ), //o
    .port_state_out_4_3_4  (keyAdd_port_state_out_4_3_4[2:0] ), //o
    .port_state_out_4_3_5  (keyAdd_port_state_out_4_3_5[2:0] ), //o
    .port_state_out_4_3_6  (keyAdd_port_state_out_4_3_6[2:0] ), //o
    .port_state_out_4_3_7  (keyAdd_port_state_out_4_3_7[2:0] ), //o
    .port_state_out_5_0_0  (keyAdd_port_state_out_5_0_0[2:0] ), //o
    .port_state_out_5_0_1  (keyAdd_port_state_out_5_0_1[2:0] ), //o
    .port_state_out_5_0_2  (keyAdd_port_state_out_5_0_2[2:0] ), //o
    .port_state_out_5_0_3  (keyAdd_port_state_out_5_0_3[2:0] ), //o
    .port_state_out_5_0_4  (keyAdd_port_state_out_5_0_4[2:0] ), //o
    .port_state_out_5_0_5  (keyAdd_port_state_out_5_0_5[2:0] ), //o
    .port_state_out_5_0_6  (keyAdd_port_state_out_5_0_6[2:0] ), //o
    .port_state_out_5_0_7  (keyAdd_port_state_out_5_0_7[2:0] ), //o
    .port_state_out_5_1_0  (keyAdd_port_state_out_5_1_0[2:0] ), //o
    .port_state_out_5_1_1  (keyAdd_port_state_out_5_1_1[2:0] ), //o
    .port_state_out_5_1_2  (keyAdd_port_state_out_5_1_2[2:0] ), //o
    .port_state_out_5_1_3  (keyAdd_port_state_out_5_1_3[2:0] ), //o
    .port_state_out_5_1_4  (keyAdd_port_state_out_5_1_4[2:0] ), //o
    .port_state_out_5_1_5  (keyAdd_port_state_out_5_1_5[2:0] ), //o
    .port_state_out_5_1_6  (keyAdd_port_state_out_5_1_6[2:0] ), //o
    .port_state_out_5_1_7  (keyAdd_port_state_out_5_1_7[2:0] ), //o
    .port_state_out_5_2_0  (keyAdd_port_state_out_5_2_0[2:0] ), //o
    .port_state_out_5_2_1  (keyAdd_port_state_out_5_2_1[2:0] ), //o
    .port_state_out_5_2_2  (keyAdd_port_state_out_5_2_2[2:0] ), //o
    .port_state_out_5_2_3  (keyAdd_port_state_out_5_2_3[2:0] ), //o
    .port_state_out_5_2_4  (keyAdd_port_state_out_5_2_4[2:0] ), //o
    .port_state_out_5_2_5  (keyAdd_port_state_out_5_2_5[2:0] ), //o
    .port_state_out_5_2_6  (keyAdd_port_state_out_5_2_6[2:0] ), //o
    .port_state_out_5_2_7  (keyAdd_port_state_out_5_2_7[2:0] ), //o
    .port_state_out_5_3_0  (keyAdd_port_state_out_5_3_0[2:0] ), //o
    .port_state_out_5_3_1  (keyAdd_port_state_out_5_3_1[2:0] ), //o
    .port_state_out_5_3_2  (keyAdd_port_state_out_5_3_2[2:0] ), //o
    .port_state_out_5_3_3  (keyAdd_port_state_out_5_3_3[2:0] ), //o
    .port_state_out_5_3_4  (keyAdd_port_state_out_5_3_4[2:0] ), //o
    .port_state_out_5_3_5  (keyAdd_port_state_out_5_3_5[2:0] ), //o
    .port_state_out_5_3_6  (keyAdd_port_state_out_5_3_6[2:0] ), //o
    .port_state_out_5_3_7  (keyAdd_port_state_out_5_3_7[2:0] ), //o
    .port_state_out_6_0_0  (keyAdd_port_state_out_6_0_0[2:0] ), //o
    .port_state_out_6_0_1  (keyAdd_port_state_out_6_0_1[2:0] ), //o
    .port_state_out_6_0_2  (keyAdd_port_state_out_6_0_2[2:0] ), //o
    .port_state_out_6_0_3  (keyAdd_port_state_out_6_0_3[2:0] ), //o
    .port_state_out_6_0_4  (keyAdd_port_state_out_6_0_4[2:0] ), //o
    .port_state_out_6_0_5  (keyAdd_port_state_out_6_0_5[2:0] ), //o
    .port_state_out_6_0_6  (keyAdd_port_state_out_6_0_6[2:0] ), //o
    .port_state_out_6_0_7  (keyAdd_port_state_out_6_0_7[2:0] ), //o
    .port_state_out_6_1_0  (keyAdd_port_state_out_6_1_0[2:0] ), //o
    .port_state_out_6_1_1  (keyAdd_port_state_out_6_1_1[2:0] ), //o
    .port_state_out_6_1_2  (keyAdd_port_state_out_6_1_2[2:0] ), //o
    .port_state_out_6_1_3  (keyAdd_port_state_out_6_1_3[2:0] ), //o
    .port_state_out_6_1_4  (keyAdd_port_state_out_6_1_4[2:0] ), //o
    .port_state_out_6_1_5  (keyAdd_port_state_out_6_1_5[2:0] ), //o
    .port_state_out_6_1_6  (keyAdd_port_state_out_6_1_6[2:0] ), //o
    .port_state_out_6_1_7  (keyAdd_port_state_out_6_1_7[2:0] ), //o
    .port_state_out_6_2_0  (keyAdd_port_state_out_6_2_0[2:0] ), //o
    .port_state_out_6_2_1  (keyAdd_port_state_out_6_2_1[2:0] ), //o
    .port_state_out_6_2_2  (keyAdd_port_state_out_6_2_2[2:0] ), //o
    .port_state_out_6_2_3  (keyAdd_port_state_out_6_2_3[2:0] ), //o
    .port_state_out_6_2_4  (keyAdd_port_state_out_6_2_4[2:0] ), //o
    .port_state_out_6_2_5  (keyAdd_port_state_out_6_2_5[2:0] ), //o
    .port_state_out_6_2_6  (keyAdd_port_state_out_6_2_6[2:0] ), //o
    .port_state_out_6_2_7  (keyAdd_port_state_out_6_2_7[2:0] ), //o
    .port_state_out_6_3_0  (keyAdd_port_state_out_6_3_0[2:0] ), //o
    .port_state_out_6_3_1  (keyAdd_port_state_out_6_3_1[2:0] ), //o
    .port_state_out_6_3_2  (keyAdd_port_state_out_6_3_2[2:0] ), //o
    .port_state_out_6_3_3  (keyAdd_port_state_out_6_3_3[2:0] ), //o
    .port_state_out_6_3_4  (keyAdd_port_state_out_6_3_4[2:0] ), //o
    .port_state_out_6_3_5  (keyAdd_port_state_out_6_3_5[2:0] ), //o
    .port_state_out_6_3_6  (keyAdd_port_state_out_6_3_6[2:0] ), //o
    .port_state_out_6_3_7  (keyAdd_port_state_out_6_3_7[2:0] ), //o
    .port_state_out_7_0_0  (keyAdd_port_state_out_7_0_0[2:0] ), //o
    .port_state_out_7_0_1  (keyAdd_port_state_out_7_0_1[2:0] ), //o
    .port_state_out_7_0_2  (keyAdd_port_state_out_7_0_2[2:0] ), //o
    .port_state_out_7_0_3  (keyAdd_port_state_out_7_0_3[2:0] ), //o
    .port_state_out_7_0_4  (keyAdd_port_state_out_7_0_4[2:0] ), //o
    .port_state_out_7_0_5  (keyAdd_port_state_out_7_0_5[2:0] ), //o
    .port_state_out_7_0_6  (keyAdd_port_state_out_7_0_6[2:0] ), //o
    .port_state_out_7_0_7  (keyAdd_port_state_out_7_0_7[2:0] ), //o
    .port_state_out_7_1_0  (keyAdd_port_state_out_7_1_0[2:0] ), //o
    .port_state_out_7_1_1  (keyAdd_port_state_out_7_1_1[2:0] ), //o
    .port_state_out_7_1_2  (keyAdd_port_state_out_7_1_2[2:0] ), //o
    .port_state_out_7_1_3  (keyAdd_port_state_out_7_1_3[2:0] ), //o
    .port_state_out_7_1_4  (keyAdd_port_state_out_7_1_4[2:0] ), //o
    .port_state_out_7_1_5  (keyAdd_port_state_out_7_1_5[2:0] ), //o
    .port_state_out_7_1_6  (keyAdd_port_state_out_7_1_6[2:0] ), //o
    .port_state_out_7_1_7  (keyAdd_port_state_out_7_1_7[2:0] ), //o
    .port_state_out_7_2_0  (keyAdd_port_state_out_7_2_0[2:0] ), //o
    .port_state_out_7_2_1  (keyAdd_port_state_out_7_2_1[2:0] ), //o
    .port_state_out_7_2_2  (keyAdd_port_state_out_7_2_2[2:0] ), //o
    .port_state_out_7_2_3  (keyAdd_port_state_out_7_2_3[2:0] ), //o
    .port_state_out_7_2_4  (keyAdd_port_state_out_7_2_4[2:0] ), //o
    .port_state_out_7_2_5  (keyAdd_port_state_out_7_2_5[2:0] ), //o
    .port_state_out_7_2_6  (keyAdd_port_state_out_7_2_6[2:0] ), //o
    .port_state_out_7_2_7  (keyAdd_port_state_out_7_2_7[2:0] ), //o
    .port_state_out_7_3_0  (keyAdd_port_state_out_7_3_0[2:0] ), //o
    .port_state_out_7_3_1  (keyAdd_port_state_out_7_3_1[2:0] ), //o
    .port_state_out_7_3_2  (keyAdd_port_state_out_7_3_2[2:0] ), //o
    .port_state_out_7_3_3  (keyAdd_port_state_out_7_3_3[2:0] ), //o
    .port_state_out_7_3_4  (keyAdd_port_state_out_7_3_4[2:0] ), //o
    .port_state_out_7_3_5  (keyAdd_port_state_out_7_3_5[2:0] ), //o
    .port_state_out_7_3_6  (keyAdd_port_state_out_7_3_6[2:0] ), //o
    .port_state_out_7_3_7  (keyAdd_port_state_out_7_3_7[2:0] ), //o
    .port_state_out_8_0_0  (keyAdd_port_state_out_8_0_0[2:0] ), //o
    .port_state_out_8_0_1  (keyAdd_port_state_out_8_0_1[2:0] ), //o
    .port_state_out_8_0_2  (keyAdd_port_state_out_8_0_2[2:0] ), //o
    .port_state_out_8_0_3  (keyAdd_port_state_out_8_0_3[2:0] ), //o
    .port_state_out_8_0_4  (keyAdd_port_state_out_8_0_4[2:0] ), //o
    .port_state_out_8_0_5  (keyAdd_port_state_out_8_0_5[2:0] ), //o
    .port_state_out_8_0_6  (keyAdd_port_state_out_8_0_6[2:0] ), //o
    .port_state_out_8_0_7  (keyAdd_port_state_out_8_0_7[2:0] ), //o
    .port_state_out_8_1_0  (keyAdd_port_state_out_8_1_0[2:0] ), //o
    .port_state_out_8_1_1  (keyAdd_port_state_out_8_1_1[2:0] ), //o
    .port_state_out_8_1_2  (keyAdd_port_state_out_8_1_2[2:0] ), //o
    .port_state_out_8_1_3  (keyAdd_port_state_out_8_1_3[2:0] ), //o
    .port_state_out_8_1_4  (keyAdd_port_state_out_8_1_4[2:0] ), //o
    .port_state_out_8_1_5  (keyAdd_port_state_out_8_1_5[2:0] ), //o
    .port_state_out_8_1_6  (keyAdd_port_state_out_8_1_6[2:0] ), //o
    .port_state_out_8_1_7  (keyAdd_port_state_out_8_1_7[2:0] ), //o
    .port_state_out_8_2_0  (keyAdd_port_state_out_8_2_0[2:0] ), //o
    .port_state_out_8_2_1  (keyAdd_port_state_out_8_2_1[2:0] ), //o
    .port_state_out_8_2_2  (keyAdd_port_state_out_8_2_2[2:0] ), //o
    .port_state_out_8_2_3  (keyAdd_port_state_out_8_2_3[2:0] ), //o
    .port_state_out_8_2_4  (keyAdd_port_state_out_8_2_4[2:0] ), //o
    .port_state_out_8_2_5  (keyAdd_port_state_out_8_2_5[2:0] ), //o
    .port_state_out_8_2_6  (keyAdd_port_state_out_8_2_6[2:0] ), //o
    .port_state_out_8_2_7  (keyAdd_port_state_out_8_2_7[2:0] ), //o
    .port_state_out_8_3_0  (keyAdd_port_state_out_8_3_0[2:0] ), //o
    .port_state_out_8_3_1  (keyAdd_port_state_out_8_3_1[2:0] ), //o
    .port_state_out_8_3_2  (keyAdd_port_state_out_8_3_2[2:0] ), //o
    .port_state_out_8_3_3  (keyAdd_port_state_out_8_3_3[2:0] ), //o
    .port_state_out_8_3_4  (keyAdd_port_state_out_8_3_4[2:0] ), //o
    .port_state_out_8_3_5  (keyAdd_port_state_out_8_3_5[2:0] ), //o
    .port_state_out_8_3_6  (keyAdd_port_state_out_8_3_6[2:0] ), //o
    .port_state_out_8_3_7  (keyAdd_port_state_out_8_3_7[2:0] ), //o
    .port_state_out_9_0_0  (keyAdd_port_state_out_9_0_0[2:0] ), //o
    .port_state_out_9_0_1  (keyAdd_port_state_out_9_0_1[2:0] ), //o
    .port_state_out_9_0_2  (keyAdd_port_state_out_9_0_2[2:0] ), //o
    .port_state_out_9_0_3  (keyAdd_port_state_out_9_0_3[2:0] ), //o
    .port_state_out_9_0_4  (keyAdd_port_state_out_9_0_4[2:0] ), //o
    .port_state_out_9_0_5  (keyAdd_port_state_out_9_0_5[2:0] ), //o
    .port_state_out_9_0_6  (keyAdd_port_state_out_9_0_6[2:0] ), //o
    .port_state_out_9_0_7  (keyAdd_port_state_out_9_0_7[2:0] ), //o
    .port_state_out_9_1_0  (keyAdd_port_state_out_9_1_0[2:0] ), //o
    .port_state_out_9_1_1  (keyAdd_port_state_out_9_1_1[2:0] ), //o
    .port_state_out_9_1_2  (keyAdd_port_state_out_9_1_2[2:0] ), //o
    .port_state_out_9_1_3  (keyAdd_port_state_out_9_1_3[2:0] ), //o
    .port_state_out_9_1_4  (keyAdd_port_state_out_9_1_4[2:0] ), //o
    .port_state_out_9_1_5  (keyAdd_port_state_out_9_1_5[2:0] ), //o
    .port_state_out_9_1_6  (keyAdd_port_state_out_9_1_6[2:0] ), //o
    .port_state_out_9_1_7  (keyAdd_port_state_out_9_1_7[2:0] ), //o
    .port_state_out_9_2_0  (keyAdd_port_state_out_9_2_0[2:0] ), //o
    .port_state_out_9_2_1  (keyAdd_port_state_out_9_2_1[2:0] ), //o
    .port_state_out_9_2_2  (keyAdd_port_state_out_9_2_2[2:0] ), //o
    .port_state_out_9_2_3  (keyAdd_port_state_out_9_2_3[2:0] ), //o
    .port_state_out_9_2_4  (keyAdd_port_state_out_9_2_4[2:0] ), //o
    .port_state_out_9_2_5  (keyAdd_port_state_out_9_2_5[2:0] ), //o
    .port_state_out_9_2_6  (keyAdd_port_state_out_9_2_6[2:0] ), //o
    .port_state_out_9_2_7  (keyAdd_port_state_out_9_2_7[2:0] ), //o
    .port_state_out_9_3_0  (keyAdd_port_state_out_9_3_0[2:0] ), //o
    .port_state_out_9_3_1  (keyAdd_port_state_out_9_3_1[2:0] ), //o
    .port_state_out_9_3_2  (keyAdd_port_state_out_9_3_2[2:0] ), //o
    .port_state_out_9_3_3  (keyAdd_port_state_out_9_3_3[2:0] ), //o
    .port_state_out_9_3_4  (keyAdd_port_state_out_9_3_4[2:0] ), //o
    .port_state_out_9_3_5  (keyAdd_port_state_out_9_3_5[2:0] ), //o
    .port_state_out_9_3_6  (keyAdd_port_state_out_9_3_6[2:0] ), //o
    .port_state_out_9_3_7  (keyAdd_port_state_out_9_3_7[2:0] ), //o
    .port_state_out_10_0_0 (keyAdd_port_state_out_10_0_0[2:0]), //o
    .port_state_out_10_0_1 (keyAdd_port_state_out_10_0_1[2:0]), //o
    .port_state_out_10_0_2 (keyAdd_port_state_out_10_0_2[2:0]), //o
    .port_state_out_10_0_3 (keyAdd_port_state_out_10_0_3[2:0]), //o
    .port_state_out_10_0_4 (keyAdd_port_state_out_10_0_4[2:0]), //o
    .port_state_out_10_0_5 (keyAdd_port_state_out_10_0_5[2:0]), //o
    .port_state_out_10_0_6 (keyAdd_port_state_out_10_0_6[2:0]), //o
    .port_state_out_10_0_7 (keyAdd_port_state_out_10_0_7[2:0]), //o
    .port_state_out_10_1_0 (keyAdd_port_state_out_10_1_0[2:0]), //o
    .port_state_out_10_1_1 (keyAdd_port_state_out_10_1_1[2:0]), //o
    .port_state_out_10_1_2 (keyAdd_port_state_out_10_1_2[2:0]), //o
    .port_state_out_10_1_3 (keyAdd_port_state_out_10_1_3[2:0]), //o
    .port_state_out_10_1_4 (keyAdd_port_state_out_10_1_4[2:0]), //o
    .port_state_out_10_1_5 (keyAdd_port_state_out_10_1_5[2:0]), //o
    .port_state_out_10_1_6 (keyAdd_port_state_out_10_1_6[2:0]), //o
    .port_state_out_10_1_7 (keyAdd_port_state_out_10_1_7[2:0]), //o
    .port_state_out_10_2_0 (keyAdd_port_state_out_10_2_0[2:0]), //o
    .port_state_out_10_2_1 (keyAdd_port_state_out_10_2_1[2:0]), //o
    .port_state_out_10_2_2 (keyAdd_port_state_out_10_2_2[2:0]), //o
    .port_state_out_10_2_3 (keyAdd_port_state_out_10_2_3[2:0]), //o
    .port_state_out_10_2_4 (keyAdd_port_state_out_10_2_4[2:0]), //o
    .port_state_out_10_2_5 (keyAdd_port_state_out_10_2_5[2:0]), //o
    .port_state_out_10_2_6 (keyAdd_port_state_out_10_2_6[2:0]), //o
    .port_state_out_10_2_7 (keyAdd_port_state_out_10_2_7[2:0]), //o
    .port_state_out_10_3_0 (keyAdd_port_state_out_10_3_0[2:0]), //o
    .port_state_out_10_3_1 (keyAdd_port_state_out_10_3_1[2:0]), //o
    .port_state_out_10_3_2 (keyAdd_port_state_out_10_3_2[2:0]), //o
    .port_state_out_10_3_3 (keyAdd_port_state_out_10_3_3[2:0]), //o
    .port_state_out_10_3_4 (keyAdd_port_state_out_10_3_4[2:0]), //o
    .port_state_out_10_3_5 (keyAdd_port_state_out_10_3_5[2:0]), //o
    .port_state_out_10_3_6 (keyAdd_port_state_out_10_3_6[2:0]), //o
    .port_state_out_10_3_7 (keyAdd_port_state_out_10_3_7[2:0]), //o
    .port_state_out_11_0_0 (keyAdd_port_state_out_11_0_0[2:0]), //o
    .port_state_out_11_0_1 (keyAdd_port_state_out_11_0_1[2:0]), //o
    .port_state_out_11_0_2 (keyAdd_port_state_out_11_0_2[2:0]), //o
    .port_state_out_11_0_3 (keyAdd_port_state_out_11_0_3[2:0]), //o
    .port_state_out_11_0_4 (keyAdd_port_state_out_11_0_4[2:0]), //o
    .port_state_out_11_0_5 (keyAdd_port_state_out_11_0_5[2:0]), //o
    .port_state_out_11_0_6 (keyAdd_port_state_out_11_0_6[2:0]), //o
    .port_state_out_11_0_7 (keyAdd_port_state_out_11_0_7[2:0]), //o
    .port_state_out_11_1_0 (keyAdd_port_state_out_11_1_0[2:0]), //o
    .port_state_out_11_1_1 (keyAdd_port_state_out_11_1_1[2:0]), //o
    .port_state_out_11_1_2 (keyAdd_port_state_out_11_1_2[2:0]), //o
    .port_state_out_11_1_3 (keyAdd_port_state_out_11_1_3[2:0]), //o
    .port_state_out_11_1_4 (keyAdd_port_state_out_11_1_4[2:0]), //o
    .port_state_out_11_1_5 (keyAdd_port_state_out_11_1_5[2:0]), //o
    .port_state_out_11_1_6 (keyAdd_port_state_out_11_1_6[2:0]), //o
    .port_state_out_11_1_7 (keyAdd_port_state_out_11_1_7[2:0]), //o
    .port_state_out_11_2_0 (keyAdd_port_state_out_11_2_0[2:0]), //o
    .port_state_out_11_2_1 (keyAdd_port_state_out_11_2_1[2:0]), //o
    .port_state_out_11_2_2 (keyAdd_port_state_out_11_2_2[2:0]), //o
    .port_state_out_11_2_3 (keyAdd_port_state_out_11_2_3[2:0]), //o
    .port_state_out_11_2_4 (keyAdd_port_state_out_11_2_4[2:0]), //o
    .port_state_out_11_2_5 (keyAdd_port_state_out_11_2_5[2:0]), //o
    .port_state_out_11_2_6 (keyAdd_port_state_out_11_2_6[2:0]), //o
    .port_state_out_11_2_7 (keyAdd_port_state_out_11_2_7[2:0]), //o
    .port_state_out_11_3_0 (keyAdd_port_state_out_11_3_0[2:0]), //o
    .port_state_out_11_3_1 (keyAdd_port_state_out_11_3_1[2:0]), //o
    .port_state_out_11_3_2 (keyAdd_port_state_out_11_3_2[2:0]), //o
    .port_state_out_11_3_3 (keyAdd_port_state_out_11_3_3[2:0]), //o
    .port_state_out_11_3_4 (keyAdd_port_state_out_11_3_4[2:0]), //o
    .port_state_out_11_3_5 (keyAdd_port_state_out_11_3_5[2:0]), //o
    .port_state_out_11_3_6 (keyAdd_port_state_out_11_3_6[2:0]), //o
    .port_state_out_11_3_7 (keyAdd_port_state_out_11_3_7[2:0]), //o
    .port_state_out_12_0_0 (keyAdd_port_state_out_12_0_0[2:0]), //o
    .port_state_out_12_0_1 (keyAdd_port_state_out_12_0_1[2:0]), //o
    .port_state_out_12_0_2 (keyAdd_port_state_out_12_0_2[2:0]), //o
    .port_state_out_12_0_3 (keyAdd_port_state_out_12_0_3[2:0]), //o
    .port_state_out_12_0_4 (keyAdd_port_state_out_12_0_4[2:0]), //o
    .port_state_out_12_0_5 (keyAdd_port_state_out_12_0_5[2:0]), //o
    .port_state_out_12_0_6 (keyAdd_port_state_out_12_0_6[2:0]), //o
    .port_state_out_12_0_7 (keyAdd_port_state_out_12_0_7[2:0]), //o
    .port_state_out_12_1_0 (keyAdd_port_state_out_12_1_0[2:0]), //o
    .port_state_out_12_1_1 (keyAdd_port_state_out_12_1_1[2:0]), //o
    .port_state_out_12_1_2 (keyAdd_port_state_out_12_1_2[2:0]), //o
    .port_state_out_12_1_3 (keyAdd_port_state_out_12_1_3[2:0]), //o
    .port_state_out_12_1_4 (keyAdd_port_state_out_12_1_4[2:0]), //o
    .port_state_out_12_1_5 (keyAdd_port_state_out_12_1_5[2:0]), //o
    .port_state_out_12_1_6 (keyAdd_port_state_out_12_1_6[2:0]), //o
    .port_state_out_12_1_7 (keyAdd_port_state_out_12_1_7[2:0]), //o
    .port_state_out_12_2_0 (keyAdd_port_state_out_12_2_0[2:0]), //o
    .port_state_out_12_2_1 (keyAdd_port_state_out_12_2_1[2:0]), //o
    .port_state_out_12_2_2 (keyAdd_port_state_out_12_2_2[2:0]), //o
    .port_state_out_12_2_3 (keyAdd_port_state_out_12_2_3[2:0]), //o
    .port_state_out_12_2_4 (keyAdd_port_state_out_12_2_4[2:0]), //o
    .port_state_out_12_2_5 (keyAdd_port_state_out_12_2_5[2:0]), //o
    .port_state_out_12_2_6 (keyAdd_port_state_out_12_2_6[2:0]), //o
    .port_state_out_12_2_7 (keyAdd_port_state_out_12_2_7[2:0]), //o
    .port_state_out_12_3_0 (keyAdd_port_state_out_12_3_0[2:0]), //o
    .port_state_out_12_3_1 (keyAdd_port_state_out_12_3_1[2:0]), //o
    .port_state_out_12_3_2 (keyAdd_port_state_out_12_3_2[2:0]), //o
    .port_state_out_12_3_3 (keyAdd_port_state_out_12_3_3[2:0]), //o
    .port_state_out_12_3_4 (keyAdd_port_state_out_12_3_4[2:0]), //o
    .port_state_out_12_3_5 (keyAdd_port_state_out_12_3_5[2:0]), //o
    .port_state_out_12_3_6 (keyAdd_port_state_out_12_3_6[2:0]), //o
    .port_state_out_12_3_7 (keyAdd_port_state_out_12_3_7[2:0]), //o
    .port_state_out_13_0_0 (keyAdd_port_state_out_13_0_0[2:0]), //o
    .port_state_out_13_0_1 (keyAdd_port_state_out_13_0_1[2:0]), //o
    .port_state_out_13_0_2 (keyAdd_port_state_out_13_0_2[2:0]), //o
    .port_state_out_13_0_3 (keyAdd_port_state_out_13_0_3[2:0]), //o
    .port_state_out_13_0_4 (keyAdd_port_state_out_13_0_4[2:0]), //o
    .port_state_out_13_0_5 (keyAdd_port_state_out_13_0_5[2:0]), //o
    .port_state_out_13_0_6 (keyAdd_port_state_out_13_0_6[2:0]), //o
    .port_state_out_13_0_7 (keyAdd_port_state_out_13_0_7[2:0]), //o
    .port_state_out_13_1_0 (keyAdd_port_state_out_13_1_0[2:0]), //o
    .port_state_out_13_1_1 (keyAdd_port_state_out_13_1_1[2:0]), //o
    .port_state_out_13_1_2 (keyAdd_port_state_out_13_1_2[2:0]), //o
    .port_state_out_13_1_3 (keyAdd_port_state_out_13_1_3[2:0]), //o
    .port_state_out_13_1_4 (keyAdd_port_state_out_13_1_4[2:0]), //o
    .port_state_out_13_1_5 (keyAdd_port_state_out_13_1_5[2:0]), //o
    .port_state_out_13_1_6 (keyAdd_port_state_out_13_1_6[2:0]), //o
    .port_state_out_13_1_7 (keyAdd_port_state_out_13_1_7[2:0]), //o
    .port_state_out_13_2_0 (keyAdd_port_state_out_13_2_0[2:0]), //o
    .port_state_out_13_2_1 (keyAdd_port_state_out_13_2_1[2:0]), //o
    .port_state_out_13_2_2 (keyAdd_port_state_out_13_2_2[2:0]), //o
    .port_state_out_13_2_3 (keyAdd_port_state_out_13_2_3[2:0]), //o
    .port_state_out_13_2_4 (keyAdd_port_state_out_13_2_4[2:0]), //o
    .port_state_out_13_2_5 (keyAdd_port_state_out_13_2_5[2:0]), //o
    .port_state_out_13_2_6 (keyAdd_port_state_out_13_2_6[2:0]), //o
    .port_state_out_13_2_7 (keyAdd_port_state_out_13_2_7[2:0]), //o
    .port_state_out_13_3_0 (keyAdd_port_state_out_13_3_0[2:0]), //o
    .port_state_out_13_3_1 (keyAdd_port_state_out_13_3_1[2:0]), //o
    .port_state_out_13_3_2 (keyAdd_port_state_out_13_3_2[2:0]), //o
    .port_state_out_13_3_3 (keyAdd_port_state_out_13_3_3[2:0]), //o
    .port_state_out_13_3_4 (keyAdd_port_state_out_13_3_4[2:0]), //o
    .port_state_out_13_3_5 (keyAdd_port_state_out_13_3_5[2:0]), //o
    .port_state_out_13_3_6 (keyAdd_port_state_out_13_3_6[2:0]), //o
    .port_state_out_13_3_7 (keyAdd_port_state_out_13_3_7[2:0]), //o
    .port_state_out_14_0_0 (keyAdd_port_state_out_14_0_0[2:0]), //o
    .port_state_out_14_0_1 (keyAdd_port_state_out_14_0_1[2:0]), //o
    .port_state_out_14_0_2 (keyAdd_port_state_out_14_0_2[2:0]), //o
    .port_state_out_14_0_3 (keyAdd_port_state_out_14_0_3[2:0]), //o
    .port_state_out_14_0_4 (keyAdd_port_state_out_14_0_4[2:0]), //o
    .port_state_out_14_0_5 (keyAdd_port_state_out_14_0_5[2:0]), //o
    .port_state_out_14_0_6 (keyAdd_port_state_out_14_0_6[2:0]), //o
    .port_state_out_14_0_7 (keyAdd_port_state_out_14_0_7[2:0]), //o
    .port_state_out_14_1_0 (keyAdd_port_state_out_14_1_0[2:0]), //o
    .port_state_out_14_1_1 (keyAdd_port_state_out_14_1_1[2:0]), //o
    .port_state_out_14_1_2 (keyAdd_port_state_out_14_1_2[2:0]), //o
    .port_state_out_14_1_3 (keyAdd_port_state_out_14_1_3[2:0]), //o
    .port_state_out_14_1_4 (keyAdd_port_state_out_14_1_4[2:0]), //o
    .port_state_out_14_1_5 (keyAdd_port_state_out_14_1_5[2:0]), //o
    .port_state_out_14_1_6 (keyAdd_port_state_out_14_1_6[2:0]), //o
    .port_state_out_14_1_7 (keyAdd_port_state_out_14_1_7[2:0]), //o
    .port_state_out_14_2_0 (keyAdd_port_state_out_14_2_0[2:0]), //o
    .port_state_out_14_2_1 (keyAdd_port_state_out_14_2_1[2:0]), //o
    .port_state_out_14_2_2 (keyAdd_port_state_out_14_2_2[2:0]), //o
    .port_state_out_14_2_3 (keyAdd_port_state_out_14_2_3[2:0]), //o
    .port_state_out_14_2_4 (keyAdd_port_state_out_14_2_4[2:0]), //o
    .port_state_out_14_2_5 (keyAdd_port_state_out_14_2_5[2:0]), //o
    .port_state_out_14_2_6 (keyAdd_port_state_out_14_2_6[2:0]), //o
    .port_state_out_14_2_7 (keyAdd_port_state_out_14_2_7[2:0]), //o
    .port_state_out_14_3_0 (keyAdd_port_state_out_14_3_0[2:0]), //o
    .port_state_out_14_3_1 (keyAdd_port_state_out_14_3_1[2:0]), //o
    .port_state_out_14_3_2 (keyAdd_port_state_out_14_3_2[2:0]), //o
    .port_state_out_14_3_3 (keyAdd_port_state_out_14_3_3[2:0]), //o
    .port_state_out_14_3_4 (keyAdd_port_state_out_14_3_4[2:0]), //o
    .port_state_out_14_3_5 (keyAdd_port_state_out_14_3_5[2:0]), //o
    .port_state_out_14_3_6 (keyAdd_port_state_out_14_3_6[2:0]), //o
    .port_state_out_14_3_7 (keyAdd_port_state_out_14_3_7[2:0]), //o
    .port_state_out_15_0_0 (keyAdd_port_state_out_15_0_0[2:0]), //o
    .port_state_out_15_0_1 (keyAdd_port_state_out_15_0_1[2:0]), //o
    .port_state_out_15_0_2 (keyAdd_port_state_out_15_0_2[2:0]), //o
    .port_state_out_15_0_3 (keyAdd_port_state_out_15_0_3[2:0]), //o
    .port_state_out_15_0_4 (keyAdd_port_state_out_15_0_4[2:0]), //o
    .port_state_out_15_0_5 (keyAdd_port_state_out_15_0_5[2:0]), //o
    .port_state_out_15_0_6 (keyAdd_port_state_out_15_0_6[2:0]), //o
    .port_state_out_15_0_7 (keyAdd_port_state_out_15_0_7[2:0]), //o
    .port_state_out_15_1_0 (keyAdd_port_state_out_15_1_0[2:0]), //o
    .port_state_out_15_1_1 (keyAdd_port_state_out_15_1_1[2:0]), //o
    .port_state_out_15_1_2 (keyAdd_port_state_out_15_1_2[2:0]), //o
    .port_state_out_15_1_3 (keyAdd_port_state_out_15_1_3[2:0]), //o
    .port_state_out_15_1_4 (keyAdd_port_state_out_15_1_4[2:0]), //o
    .port_state_out_15_1_5 (keyAdd_port_state_out_15_1_5[2:0]), //o
    .port_state_out_15_1_6 (keyAdd_port_state_out_15_1_6[2:0]), //o
    .port_state_out_15_1_7 (keyAdd_port_state_out_15_1_7[2:0]), //o
    .port_state_out_15_2_0 (keyAdd_port_state_out_15_2_0[2:0]), //o
    .port_state_out_15_2_1 (keyAdd_port_state_out_15_2_1[2:0]), //o
    .port_state_out_15_2_2 (keyAdd_port_state_out_15_2_2[2:0]), //o
    .port_state_out_15_2_3 (keyAdd_port_state_out_15_2_3[2:0]), //o
    .port_state_out_15_2_4 (keyAdd_port_state_out_15_2_4[2:0]), //o
    .port_state_out_15_2_5 (keyAdd_port_state_out_15_2_5[2:0]), //o
    .port_state_out_15_2_6 (keyAdd_port_state_out_15_2_6[2:0]), //o
    .port_state_out_15_2_7 (keyAdd_port_state_out_15_2_7[2:0]), //o
    .port_state_out_15_3_0 (keyAdd_port_state_out_15_3_0[2:0]), //o
    .port_state_out_15_3_1 (keyAdd_port_state_out_15_3_1[2:0]), //o
    .port_state_out_15_3_2 (keyAdd_port_state_out_15_3_2[2:0]), //o
    .port_state_out_15_3_3 (keyAdd_port_state_out_15_3_3[2:0]), //o
    .port_state_out_15_3_4 (keyAdd_port_state_out_15_3_4[2:0]), //o
    .port_state_out_15_3_5 (keyAdd_port_state_out_15_3_5[2:0]), //o
    .port_state_out_15_3_6 (keyAdd_port_state_out_15_3_6[2:0]), //o
    .port_state_out_15_3_7 (keyAdd_port_state_out_15_3_7[2:0])  //o
  );
  Sbox_AES_BoyarPeralta sbox_AES_BoyarPeralta_16 (
    .port_i_0_0 (keyAdd_port_state_out_0_0_0[2:0]        ), //i
    .port_i_0_1 (keyAdd_port_state_out_0_0_1[2:0]        ), //i
    .port_i_0_2 (keyAdd_port_state_out_0_0_2[2:0]        ), //i
    .port_i_0_3 (keyAdd_port_state_out_0_0_3[2:0]        ), //i
    .port_i_0_4 (keyAdd_port_state_out_0_0_4[2:0]        ), //i
    .port_i_0_5 (keyAdd_port_state_out_0_0_5[2:0]        ), //i
    .port_i_0_6 (keyAdd_port_state_out_0_0_6[2:0]        ), //i
    .port_i_0_7 (keyAdd_port_state_out_0_0_7[2:0]        ), //i
    .port_i_1_0 (keyAdd_port_state_out_0_1_0[2:0]        ), //i
    .port_i_1_1 (keyAdd_port_state_out_0_1_1[2:0]        ), //i
    .port_i_1_2 (keyAdd_port_state_out_0_1_2[2:0]        ), //i
    .port_i_1_3 (keyAdd_port_state_out_0_1_3[2:0]        ), //i
    .port_i_1_4 (keyAdd_port_state_out_0_1_4[2:0]        ), //i
    .port_i_1_5 (keyAdd_port_state_out_0_1_5[2:0]        ), //i
    .port_i_1_6 (keyAdd_port_state_out_0_1_6[2:0]        ), //i
    .port_i_1_7 (keyAdd_port_state_out_0_1_7[2:0]        ), //i
    .port_i_2_0 (keyAdd_port_state_out_0_2_0[2:0]        ), //i
    .port_i_2_1 (keyAdd_port_state_out_0_2_1[2:0]        ), //i
    .port_i_2_2 (keyAdd_port_state_out_0_2_2[2:0]        ), //i
    .port_i_2_3 (keyAdd_port_state_out_0_2_3[2:0]        ), //i
    .port_i_2_4 (keyAdd_port_state_out_0_2_4[2:0]        ), //i
    .port_i_2_5 (keyAdd_port_state_out_0_2_5[2:0]        ), //i
    .port_i_2_6 (keyAdd_port_state_out_0_2_6[2:0]        ), //i
    .port_i_2_7 (keyAdd_port_state_out_0_2_7[2:0]        ), //i
    .port_i_3_0 (keyAdd_port_state_out_0_3_0[2:0]        ), //i
    .port_i_3_1 (keyAdd_port_state_out_0_3_1[2:0]        ), //i
    .port_i_3_2 (keyAdd_port_state_out_0_3_2[2:0]        ), //i
    .port_i_3_3 (keyAdd_port_state_out_0_3_3[2:0]        ), //i
    .port_i_3_4 (keyAdd_port_state_out_0_3_4[2:0]        ), //i
    .port_i_3_5 (keyAdd_port_state_out_0_3_5[2:0]        ), //i
    .port_i_3_6 (keyAdd_port_state_out_0_3_6[2:0]        ), //i
    .port_i_3_7 (keyAdd_port_state_out_0_3_7[2:0]        ), //i
    .port_o_0_0 (sbox_AES_BoyarPeralta_16_port_o_0_0[2:0]), //o
    .port_o_0_1 (sbox_AES_BoyarPeralta_16_port_o_0_1[2:0]), //o
    .port_o_0_2 (sbox_AES_BoyarPeralta_16_port_o_0_2[2:0]), //o
    .port_o_0_3 (sbox_AES_BoyarPeralta_16_port_o_0_3[2:0]), //o
    .port_o_0_4 (sbox_AES_BoyarPeralta_16_port_o_0_4[2:0]), //o
    .port_o_0_5 (sbox_AES_BoyarPeralta_16_port_o_0_5[2:0]), //o
    .port_o_0_6 (sbox_AES_BoyarPeralta_16_port_o_0_6[2:0]), //o
    .port_o_0_7 (sbox_AES_BoyarPeralta_16_port_o_0_7[2:0]), //o
    .port_o_1_0 (sbox_AES_BoyarPeralta_16_port_o_1_0[2:0]), //o
    .port_o_1_1 (sbox_AES_BoyarPeralta_16_port_o_1_1[2:0]), //o
    .port_o_1_2 (sbox_AES_BoyarPeralta_16_port_o_1_2[2:0]), //o
    .port_o_1_3 (sbox_AES_BoyarPeralta_16_port_o_1_3[2:0]), //o
    .port_o_1_4 (sbox_AES_BoyarPeralta_16_port_o_1_4[2:0]), //o
    .port_o_1_5 (sbox_AES_BoyarPeralta_16_port_o_1_5[2:0]), //o
    .port_o_1_6 (sbox_AES_BoyarPeralta_16_port_o_1_6[2:0]), //o
    .port_o_1_7 (sbox_AES_BoyarPeralta_16_port_o_1_7[2:0]), //o
    .port_o_2_0 (sbox_AES_BoyarPeralta_16_port_o_2_0[2:0]), //o
    .port_o_2_1 (sbox_AES_BoyarPeralta_16_port_o_2_1[2:0]), //o
    .port_o_2_2 (sbox_AES_BoyarPeralta_16_port_o_2_2[2:0]), //o
    .port_o_2_3 (sbox_AES_BoyarPeralta_16_port_o_2_3[2:0]), //o
    .port_o_2_4 (sbox_AES_BoyarPeralta_16_port_o_2_4[2:0]), //o
    .port_o_2_5 (sbox_AES_BoyarPeralta_16_port_o_2_5[2:0]), //o
    .port_o_2_6 (sbox_AES_BoyarPeralta_16_port_o_2_6[2:0]), //o
    .port_o_2_7 (sbox_AES_BoyarPeralta_16_port_o_2_7[2:0]), //o
    .port_o_3_0 (sbox_AES_BoyarPeralta_16_port_o_3_0[2:0]), //o
    .port_o_3_1 (sbox_AES_BoyarPeralta_16_port_o_3_1[2:0]), //o
    .port_o_3_2 (sbox_AES_BoyarPeralta_16_port_o_3_2[2:0]), //o
    .port_o_3_3 (sbox_AES_BoyarPeralta_16_port_o_3_3[2:0]), //o
    .port_o_3_4 (sbox_AES_BoyarPeralta_16_port_o_3_4[2:0]), //o
    .port_o_3_5 (sbox_AES_BoyarPeralta_16_port_o_3_5[2:0]), //o
    .port_o_3_6 (sbox_AES_BoyarPeralta_16_port_o_3_6[2:0]), //o
    .port_o_3_7 (sbox_AES_BoyarPeralta_16_port_o_3_7[2:0]), //o
    .clk        (clk                                     ), //i
    .reset      (reset                                   )  //i
  );
  Sbox_AES_BoyarPeralta sbox_AES_BoyarPeralta_17 (
    .port_i_0_0 (keyAdd_port_state_out_1_0_0[2:0]        ), //i
    .port_i_0_1 (keyAdd_port_state_out_1_0_1[2:0]        ), //i
    .port_i_0_2 (keyAdd_port_state_out_1_0_2[2:0]        ), //i
    .port_i_0_3 (keyAdd_port_state_out_1_0_3[2:0]        ), //i
    .port_i_0_4 (keyAdd_port_state_out_1_0_4[2:0]        ), //i
    .port_i_0_5 (keyAdd_port_state_out_1_0_5[2:0]        ), //i
    .port_i_0_6 (keyAdd_port_state_out_1_0_6[2:0]        ), //i
    .port_i_0_7 (keyAdd_port_state_out_1_0_7[2:0]        ), //i
    .port_i_1_0 (keyAdd_port_state_out_1_1_0[2:0]        ), //i
    .port_i_1_1 (keyAdd_port_state_out_1_1_1[2:0]        ), //i
    .port_i_1_2 (keyAdd_port_state_out_1_1_2[2:0]        ), //i
    .port_i_1_3 (keyAdd_port_state_out_1_1_3[2:0]        ), //i
    .port_i_1_4 (keyAdd_port_state_out_1_1_4[2:0]        ), //i
    .port_i_1_5 (keyAdd_port_state_out_1_1_5[2:0]        ), //i
    .port_i_1_6 (keyAdd_port_state_out_1_1_6[2:0]        ), //i
    .port_i_1_7 (keyAdd_port_state_out_1_1_7[2:0]        ), //i
    .port_i_2_0 (keyAdd_port_state_out_1_2_0[2:0]        ), //i
    .port_i_2_1 (keyAdd_port_state_out_1_2_1[2:0]        ), //i
    .port_i_2_2 (keyAdd_port_state_out_1_2_2[2:0]        ), //i
    .port_i_2_3 (keyAdd_port_state_out_1_2_3[2:0]        ), //i
    .port_i_2_4 (keyAdd_port_state_out_1_2_4[2:0]        ), //i
    .port_i_2_5 (keyAdd_port_state_out_1_2_5[2:0]        ), //i
    .port_i_2_6 (keyAdd_port_state_out_1_2_6[2:0]        ), //i
    .port_i_2_7 (keyAdd_port_state_out_1_2_7[2:0]        ), //i
    .port_i_3_0 (keyAdd_port_state_out_1_3_0[2:0]        ), //i
    .port_i_3_1 (keyAdd_port_state_out_1_3_1[2:0]        ), //i
    .port_i_3_2 (keyAdd_port_state_out_1_3_2[2:0]        ), //i
    .port_i_3_3 (keyAdd_port_state_out_1_3_3[2:0]        ), //i
    .port_i_3_4 (keyAdd_port_state_out_1_3_4[2:0]        ), //i
    .port_i_3_5 (keyAdd_port_state_out_1_3_5[2:0]        ), //i
    .port_i_3_6 (keyAdd_port_state_out_1_3_6[2:0]        ), //i
    .port_i_3_7 (keyAdd_port_state_out_1_3_7[2:0]        ), //i
    .port_o_0_0 (sbox_AES_BoyarPeralta_17_port_o_0_0[2:0]), //o
    .port_o_0_1 (sbox_AES_BoyarPeralta_17_port_o_0_1[2:0]), //o
    .port_o_0_2 (sbox_AES_BoyarPeralta_17_port_o_0_2[2:0]), //o
    .port_o_0_3 (sbox_AES_BoyarPeralta_17_port_o_0_3[2:0]), //o
    .port_o_0_4 (sbox_AES_BoyarPeralta_17_port_o_0_4[2:0]), //o
    .port_o_0_5 (sbox_AES_BoyarPeralta_17_port_o_0_5[2:0]), //o
    .port_o_0_6 (sbox_AES_BoyarPeralta_17_port_o_0_6[2:0]), //o
    .port_o_0_7 (sbox_AES_BoyarPeralta_17_port_o_0_7[2:0]), //o
    .port_o_1_0 (sbox_AES_BoyarPeralta_17_port_o_1_0[2:0]), //o
    .port_o_1_1 (sbox_AES_BoyarPeralta_17_port_o_1_1[2:0]), //o
    .port_o_1_2 (sbox_AES_BoyarPeralta_17_port_o_1_2[2:0]), //o
    .port_o_1_3 (sbox_AES_BoyarPeralta_17_port_o_1_3[2:0]), //o
    .port_o_1_4 (sbox_AES_BoyarPeralta_17_port_o_1_4[2:0]), //o
    .port_o_1_5 (sbox_AES_BoyarPeralta_17_port_o_1_5[2:0]), //o
    .port_o_1_6 (sbox_AES_BoyarPeralta_17_port_o_1_6[2:0]), //o
    .port_o_1_7 (sbox_AES_BoyarPeralta_17_port_o_1_7[2:0]), //o
    .port_o_2_0 (sbox_AES_BoyarPeralta_17_port_o_2_0[2:0]), //o
    .port_o_2_1 (sbox_AES_BoyarPeralta_17_port_o_2_1[2:0]), //o
    .port_o_2_2 (sbox_AES_BoyarPeralta_17_port_o_2_2[2:0]), //o
    .port_o_2_3 (sbox_AES_BoyarPeralta_17_port_o_2_3[2:0]), //o
    .port_o_2_4 (sbox_AES_BoyarPeralta_17_port_o_2_4[2:0]), //o
    .port_o_2_5 (sbox_AES_BoyarPeralta_17_port_o_2_5[2:0]), //o
    .port_o_2_6 (sbox_AES_BoyarPeralta_17_port_o_2_6[2:0]), //o
    .port_o_2_7 (sbox_AES_BoyarPeralta_17_port_o_2_7[2:0]), //o
    .port_o_3_0 (sbox_AES_BoyarPeralta_17_port_o_3_0[2:0]), //o
    .port_o_3_1 (sbox_AES_BoyarPeralta_17_port_o_3_1[2:0]), //o
    .port_o_3_2 (sbox_AES_BoyarPeralta_17_port_o_3_2[2:0]), //o
    .port_o_3_3 (sbox_AES_BoyarPeralta_17_port_o_3_3[2:0]), //o
    .port_o_3_4 (sbox_AES_BoyarPeralta_17_port_o_3_4[2:0]), //o
    .port_o_3_5 (sbox_AES_BoyarPeralta_17_port_o_3_5[2:0]), //o
    .port_o_3_6 (sbox_AES_BoyarPeralta_17_port_o_3_6[2:0]), //o
    .port_o_3_7 (sbox_AES_BoyarPeralta_17_port_o_3_7[2:0]), //o
    .clk        (clk                                     ), //i
    .reset      (reset                                   )  //i
  );
  Sbox_AES_BoyarPeralta sbox_AES_BoyarPeralta_18 (
    .port_i_0_0 (keyAdd_port_state_out_2_0_0[2:0]        ), //i
    .port_i_0_1 (keyAdd_port_state_out_2_0_1[2:0]        ), //i
    .port_i_0_2 (keyAdd_port_state_out_2_0_2[2:0]        ), //i
    .port_i_0_3 (keyAdd_port_state_out_2_0_3[2:0]        ), //i
    .port_i_0_4 (keyAdd_port_state_out_2_0_4[2:0]        ), //i
    .port_i_0_5 (keyAdd_port_state_out_2_0_5[2:0]        ), //i
    .port_i_0_6 (keyAdd_port_state_out_2_0_6[2:0]        ), //i
    .port_i_0_7 (keyAdd_port_state_out_2_0_7[2:0]        ), //i
    .port_i_1_0 (keyAdd_port_state_out_2_1_0[2:0]        ), //i
    .port_i_1_1 (keyAdd_port_state_out_2_1_1[2:0]        ), //i
    .port_i_1_2 (keyAdd_port_state_out_2_1_2[2:0]        ), //i
    .port_i_1_3 (keyAdd_port_state_out_2_1_3[2:0]        ), //i
    .port_i_1_4 (keyAdd_port_state_out_2_1_4[2:0]        ), //i
    .port_i_1_5 (keyAdd_port_state_out_2_1_5[2:0]        ), //i
    .port_i_1_6 (keyAdd_port_state_out_2_1_6[2:0]        ), //i
    .port_i_1_7 (keyAdd_port_state_out_2_1_7[2:0]        ), //i
    .port_i_2_0 (keyAdd_port_state_out_2_2_0[2:0]        ), //i
    .port_i_2_1 (keyAdd_port_state_out_2_2_1[2:0]        ), //i
    .port_i_2_2 (keyAdd_port_state_out_2_2_2[2:0]        ), //i
    .port_i_2_3 (keyAdd_port_state_out_2_2_3[2:0]        ), //i
    .port_i_2_4 (keyAdd_port_state_out_2_2_4[2:0]        ), //i
    .port_i_2_5 (keyAdd_port_state_out_2_2_5[2:0]        ), //i
    .port_i_2_6 (keyAdd_port_state_out_2_2_6[2:0]        ), //i
    .port_i_2_7 (keyAdd_port_state_out_2_2_7[2:0]        ), //i
    .port_i_3_0 (keyAdd_port_state_out_2_3_0[2:0]        ), //i
    .port_i_3_1 (keyAdd_port_state_out_2_3_1[2:0]        ), //i
    .port_i_3_2 (keyAdd_port_state_out_2_3_2[2:0]        ), //i
    .port_i_3_3 (keyAdd_port_state_out_2_3_3[2:0]        ), //i
    .port_i_3_4 (keyAdd_port_state_out_2_3_4[2:0]        ), //i
    .port_i_3_5 (keyAdd_port_state_out_2_3_5[2:0]        ), //i
    .port_i_3_6 (keyAdd_port_state_out_2_3_6[2:0]        ), //i
    .port_i_3_7 (keyAdd_port_state_out_2_3_7[2:0]        ), //i
    .port_o_0_0 (sbox_AES_BoyarPeralta_18_port_o_0_0[2:0]), //o
    .port_o_0_1 (sbox_AES_BoyarPeralta_18_port_o_0_1[2:0]), //o
    .port_o_0_2 (sbox_AES_BoyarPeralta_18_port_o_0_2[2:0]), //o
    .port_o_0_3 (sbox_AES_BoyarPeralta_18_port_o_0_3[2:0]), //o
    .port_o_0_4 (sbox_AES_BoyarPeralta_18_port_o_0_4[2:0]), //o
    .port_o_0_5 (sbox_AES_BoyarPeralta_18_port_o_0_5[2:0]), //o
    .port_o_0_6 (sbox_AES_BoyarPeralta_18_port_o_0_6[2:0]), //o
    .port_o_0_7 (sbox_AES_BoyarPeralta_18_port_o_0_7[2:0]), //o
    .port_o_1_0 (sbox_AES_BoyarPeralta_18_port_o_1_0[2:0]), //o
    .port_o_1_1 (sbox_AES_BoyarPeralta_18_port_o_1_1[2:0]), //o
    .port_o_1_2 (sbox_AES_BoyarPeralta_18_port_o_1_2[2:0]), //o
    .port_o_1_3 (sbox_AES_BoyarPeralta_18_port_o_1_3[2:0]), //o
    .port_o_1_4 (sbox_AES_BoyarPeralta_18_port_o_1_4[2:0]), //o
    .port_o_1_5 (sbox_AES_BoyarPeralta_18_port_o_1_5[2:0]), //o
    .port_o_1_6 (sbox_AES_BoyarPeralta_18_port_o_1_6[2:0]), //o
    .port_o_1_7 (sbox_AES_BoyarPeralta_18_port_o_1_7[2:0]), //o
    .port_o_2_0 (sbox_AES_BoyarPeralta_18_port_o_2_0[2:0]), //o
    .port_o_2_1 (sbox_AES_BoyarPeralta_18_port_o_2_1[2:0]), //o
    .port_o_2_2 (sbox_AES_BoyarPeralta_18_port_o_2_2[2:0]), //o
    .port_o_2_3 (sbox_AES_BoyarPeralta_18_port_o_2_3[2:0]), //o
    .port_o_2_4 (sbox_AES_BoyarPeralta_18_port_o_2_4[2:0]), //o
    .port_o_2_5 (sbox_AES_BoyarPeralta_18_port_o_2_5[2:0]), //o
    .port_o_2_6 (sbox_AES_BoyarPeralta_18_port_o_2_6[2:0]), //o
    .port_o_2_7 (sbox_AES_BoyarPeralta_18_port_o_2_7[2:0]), //o
    .port_o_3_0 (sbox_AES_BoyarPeralta_18_port_o_3_0[2:0]), //o
    .port_o_3_1 (sbox_AES_BoyarPeralta_18_port_o_3_1[2:0]), //o
    .port_o_3_2 (sbox_AES_BoyarPeralta_18_port_o_3_2[2:0]), //o
    .port_o_3_3 (sbox_AES_BoyarPeralta_18_port_o_3_3[2:0]), //o
    .port_o_3_4 (sbox_AES_BoyarPeralta_18_port_o_3_4[2:0]), //o
    .port_o_3_5 (sbox_AES_BoyarPeralta_18_port_o_3_5[2:0]), //o
    .port_o_3_6 (sbox_AES_BoyarPeralta_18_port_o_3_6[2:0]), //o
    .port_o_3_7 (sbox_AES_BoyarPeralta_18_port_o_3_7[2:0]), //o
    .clk        (clk                                     ), //i
    .reset      (reset                                   )  //i
  );
  Sbox_AES_BoyarPeralta sbox_AES_BoyarPeralta_19 (
    .port_i_0_0 (keyAdd_port_state_out_3_0_0[2:0]        ), //i
    .port_i_0_1 (keyAdd_port_state_out_3_0_1[2:0]        ), //i
    .port_i_0_2 (keyAdd_port_state_out_3_0_2[2:0]        ), //i
    .port_i_0_3 (keyAdd_port_state_out_3_0_3[2:0]        ), //i
    .port_i_0_4 (keyAdd_port_state_out_3_0_4[2:0]        ), //i
    .port_i_0_5 (keyAdd_port_state_out_3_0_5[2:0]        ), //i
    .port_i_0_6 (keyAdd_port_state_out_3_0_6[2:0]        ), //i
    .port_i_0_7 (keyAdd_port_state_out_3_0_7[2:0]        ), //i
    .port_i_1_0 (keyAdd_port_state_out_3_1_0[2:0]        ), //i
    .port_i_1_1 (keyAdd_port_state_out_3_1_1[2:0]        ), //i
    .port_i_1_2 (keyAdd_port_state_out_3_1_2[2:0]        ), //i
    .port_i_1_3 (keyAdd_port_state_out_3_1_3[2:0]        ), //i
    .port_i_1_4 (keyAdd_port_state_out_3_1_4[2:0]        ), //i
    .port_i_1_5 (keyAdd_port_state_out_3_1_5[2:0]        ), //i
    .port_i_1_6 (keyAdd_port_state_out_3_1_6[2:0]        ), //i
    .port_i_1_7 (keyAdd_port_state_out_3_1_7[2:0]        ), //i
    .port_i_2_0 (keyAdd_port_state_out_3_2_0[2:0]        ), //i
    .port_i_2_1 (keyAdd_port_state_out_3_2_1[2:0]        ), //i
    .port_i_2_2 (keyAdd_port_state_out_3_2_2[2:0]        ), //i
    .port_i_2_3 (keyAdd_port_state_out_3_2_3[2:0]        ), //i
    .port_i_2_4 (keyAdd_port_state_out_3_2_4[2:0]        ), //i
    .port_i_2_5 (keyAdd_port_state_out_3_2_5[2:0]        ), //i
    .port_i_2_6 (keyAdd_port_state_out_3_2_6[2:0]        ), //i
    .port_i_2_7 (keyAdd_port_state_out_3_2_7[2:0]        ), //i
    .port_i_3_0 (keyAdd_port_state_out_3_3_0[2:0]        ), //i
    .port_i_3_1 (keyAdd_port_state_out_3_3_1[2:0]        ), //i
    .port_i_3_2 (keyAdd_port_state_out_3_3_2[2:0]        ), //i
    .port_i_3_3 (keyAdd_port_state_out_3_3_3[2:0]        ), //i
    .port_i_3_4 (keyAdd_port_state_out_3_3_4[2:0]        ), //i
    .port_i_3_5 (keyAdd_port_state_out_3_3_5[2:0]        ), //i
    .port_i_3_6 (keyAdd_port_state_out_3_3_6[2:0]        ), //i
    .port_i_3_7 (keyAdd_port_state_out_3_3_7[2:0]        ), //i
    .port_o_0_0 (sbox_AES_BoyarPeralta_19_port_o_0_0[2:0]), //o
    .port_o_0_1 (sbox_AES_BoyarPeralta_19_port_o_0_1[2:0]), //o
    .port_o_0_2 (sbox_AES_BoyarPeralta_19_port_o_0_2[2:0]), //o
    .port_o_0_3 (sbox_AES_BoyarPeralta_19_port_o_0_3[2:0]), //o
    .port_o_0_4 (sbox_AES_BoyarPeralta_19_port_o_0_4[2:0]), //o
    .port_o_0_5 (sbox_AES_BoyarPeralta_19_port_o_0_5[2:0]), //o
    .port_o_0_6 (sbox_AES_BoyarPeralta_19_port_o_0_6[2:0]), //o
    .port_o_0_7 (sbox_AES_BoyarPeralta_19_port_o_0_7[2:0]), //o
    .port_o_1_0 (sbox_AES_BoyarPeralta_19_port_o_1_0[2:0]), //o
    .port_o_1_1 (sbox_AES_BoyarPeralta_19_port_o_1_1[2:0]), //o
    .port_o_1_2 (sbox_AES_BoyarPeralta_19_port_o_1_2[2:0]), //o
    .port_o_1_3 (sbox_AES_BoyarPeralta_19_port_o_1_3[2:0]), //o
    .port_o_1_4 (sbox_AES_BoyarPeralta_19_port_o_1_4[2:0]), //o
    .port_o_1_5 (sbox_AES_BoyarPeralta_19_port_o_1_5[2:0]), //o
    .port_o_1_6 (sbox_AES_BoyarPeralta_19_port_o_1_6[2:0]), //o
    .port_o_1_7 (sbox_AES_BoyarPeralta_19_port_o_1_7[2:0]), //o
    .port_o_2_0 (sbox_AES_BoyarPeralta_19_port_o_2_0[2:0]), //o
    .port_o_2_1 (sbox_AES_BoyarPeralta_19_port_o_2_1[2:0]), //o
    .port_o_2_2 (sbox_AES_BoyarPeralta_19_port_o_2_2[2:0]), //o
    .port_o_2_3 (sbox_AES_BoyarPeralta_19_port_o_2_3[2:0]), //o
    .port_o_2_4 (sbox_AES_BoyarPeralta_19_port_o_2_4[2:0]), //o
    .port_o_2_5 (sbox_AES_BoyarPeralta_19_port_o_2_5[2:0]), //o
    .port_o_2_6 (sbox_AES_BoyarPeralta_19_port_o_2_6[2:0]), //o
    .port_o_2_7 (sbox_AES_BoyarPeralta_19_port_o_2_7[2:0]), //o
    .port_o_3_0 (sbox_AES_BoyarPeralta_19_port_o_3_0[2:0]), //o
    .port_o_3_1 (sbox_AES_BoyarPeralta_19_port_o_3_1[2:0]), //o
    .port_o_3_2 (sbox_AES_BoyarPeralta_19_port_o_3_2[2:0]), //o
    .port_o_3_3 (sbox_AES_BoyarPeralta_19_port_o_3_3[2:0]), //o
    .port_o_3_4 (sbox_AES_BoyarPeralta_19_port_o_3_4[2:0]), //o
    .port_o_3_5 (sbox_AES_BoyarPeralta_19_port_o_3_5[2:0]), //o
    .port_o_3_6 (sbox_AES_BoyarPeralta_19_port_o_3_6[2:0]), //o
    .port_o_3_7 (sbox_AES_BoyarPeralta_19_port_o_3_7[2:0]), //o
    .clk        (clk                                     ), //i
    .reset      (reset                                   )  //i
  );
  Sbox_AES_BoyarPeralta sbox_AES_BoyarPeralta_20 (
    .port_i_0_0 (keyAdd_port_state_out_4_0_0[2:0]        ), //i
    .port_i_0_1 (keyAdd_port_state_out_4_0_1[2:0]        ), //i
    .port_i_0_2 (keyAdd_port_state_out_4_0_2[2:0]        ), //i
    .port_i_0_3 (keyAdd_port_state_out_4_0_3[2:0]        ), //i
    .port_i_0_4 (keyAdd_port_state_out_4_0_4[2:0]        ), //i
    .port_i_0_5 (keyAdd_port_state_out_4_0_5[2:0]        ), //i
    .port_i_0_6 (keyAdd_port_state_out_4_0_6[2:0]        ), //i
    .port_i_0_7 (keyAdd_port_state_out_4_0_7[2:0]        ), //i
    .port_i_1_0 (keyAdd_port_state_out_4_1_0[2:0]        ), //i
    .port_i_1_1 (keyAdd_port_state_out_4_1_1[2:0]        ), //i
    .port_i_1_2 (keyAdd_port_state_out_4_1_2[2:0]        ), //i
    .port_i_1_3 (keyAdd_port_state_out_4_1_3[2:0]        ), //i
    .port_i_1_4 (keyAdd_port_state_out_4_1_4[2:0]        ), //i
    .port_i_1_5 (keyAdd_port_state_out_4_1_5[2:0]        ), //i
    .port_i_1_6 (keyAdd_port_state_out_4_1_6[2:0]        ), //i
    .port_i_1_7 (keyAdd_port_state_out_4_1_7[2:0]        ), //i
    .port_i_2_0 (keyAdd_port_state_out_4_2_0[2:0]        ), //i
    .port_i_2_1 (keyAdd_port_state_out_4_2_1[2:0]        ), //i
    .port_i_2_2 (keyAdd_port_state_out_4_2_2[2:0]        ), //i
    .port_i_2_3 (keyAdd_port_state_out_4_2_3[2:0]        ), //i
    .port_i_2_4 (keyAdd_port_state_out_4_2_4[2:0]        ), //i
    .port_i_2_5 (keyAdd_port_state_out_4_2_5[2:0]        ), //i
    .port_i_2_6 (keyAdd_port_state_out_4_2_6[2:0]        ), //i
    .port_i_2_7 (keyAdd_port_state_out_4_2_7[2:0]        ), //i
    .port_i_3_0 (keyAdd_port_state_out_4_3_0[2:0]        ), //i
    .port_i_3_1 (keyAdd_port_state_out_4_3_1[2:0]        ), //i
    .port_i_3_2 (keyAdd_port_state_out_4_3_2[2:0]        ), //i
    .port_i_3_3 (keyAdd_port_state_out_4_3_3[2:0]        ), //i
    .port_i_3_4 (keyAdd_port_state_out_4_3_4[2:0]        ), //i
    .port_i_3_5 (keyAdd_port_state_out_4_3_5[2:0]        ), //i
    .port_i_3_6 (keyAdd_port_state_out_4_3_6[2:0]        ), //i
    .port_i_3_7 (keyAdd_port_state_out_4_3_7[2:0]        ), //i
    .port_o_0_0 (sbox_AES_BoyarPeralta_20_port_o_0_0[2:0]), //o
    .port_o_0_1 (sbox_AES_BoyarPeralta_20_port_o_0_1[2:0]), //o
    .port_o_0_2 (sbox_AES_BoyarPeralta_20_port_o_0_2[2:0]), //o
    .port_o_0_3 (sbox_AES_BoyarPeralta_20_port_o_0_3[2:0]), //o
    .port_o_0_4 (sbox_AES_BoyarPeralta_20_port_o_0_4[2:0]), //o
    .port_o_0_5 (sbox_AES_BoyarPeralta_20_port_o_0_5[2:0]), //o
    .port_o_0_6 (sbox_AES_BoyarPeralta_20_port_o_0_6[2:0]), //o
    .port_o_0_7 (sbox_AES_BoyarPeralta_20_port_o_0_7[2:0]), //o
    .port_o_1_0 (sbox_AES_BoyarPeralta_20_port_o_1_0[2:0]), //o
    .port_o_1_1 (sbox_AES_BoyarPeralta_20_port_o_1_1[2:0]), //o
    .port_o_1_2 (sbox_AES_BoyarPeralta_20_port_o_1_2[2:0]), //o
    .port_o_1_3 (sbox_AES_BoyarPeralta_20_port_o_1_3[2:0]), //o
    .port_o_1_4 (sbox_AES_BoyarPeralta_20_port_o_1_4[2:0]), //o
    .port_o_1_5 (sbox_AES_BoyarPeralta_20_port_o_1_5[2:0]), //o
    .port_o_1_6 (sbox_AES_BoyarPeralta_20_port_o_1_6[2:0]), //o
    .port_o_1_7 (sbox_AES_BoyarPeralta_20_port_o_1_7[2:0]), //o
    .port_o_2_0 (sbox_AES_BoyarPeralta_20_port_o_2_0[2:0]), //o
    .port_o_2_1 (sbox_AES_BoyarPeralta_20_port_o_2_1[2:0]), //o
    .port_o_2_2 (sbox_AES_BoyarPeralta_20_port_o_2_2[2:0]), //o
    .port_o_2_3 (sbox_AES_BoyarPeralta_20_port_o_2_3[2:0]), //o
    .port_o_2_4 (sbox_AES_BoyarPeralta_20_port_o_2_4[2:0]), //o
    .port_o_2_5 (sbox_AES_BoyarPeralta_20_port_o_2_5[2:0]), //o
    .port_o_2_6 (sbox_AES_BoyarPeralta_20_port_o_2_6[2:0]), //o
    .port_o_2_7 (sbox_AES_BoyarPeralta_20_port_o_2_7[2:0]), //o
    .port_o_3_0 (sbox_AES_BoyarPeralta_20_port_o_3_0[2:0]), //o
    .port_o_3_1 (sbox_AES_BoyarPeralta_20_port_o_3_1[2:0]), //o
    .port_o_3_2 (sbox_AES_BoyarPeralta_20_port_o_3_2[2:0]), //o
    .port_o_3_3 (sbox_AES_BoyarPeralta_20_port_o_3_3[2:0]), //o
    .port_o_3_4 (sbox_AES_BoyarPeralta_20_port_o_3_4[2:0]), //o
    .port_o_3_5 (sbox_AES_BoyarPeralta_20_port_o_3_5[2:0]), //o
    .port_o_3_6 (sbox_AES_BoyarPeralta_20_port_o_3_6[2:0]), //o
    .port_o_3_7 (sbox_AES_BoyarPeralta_20_port_o_3_7[2:0]), //o
    .clk        (clk                                     ), //i
    .reset      (reset                                   )  //i
  );
  Sbox_AES_BoyarPeralta sbox_AES_BoyarPeralta_21 (
    .port_i_0_0 (keyAdd_port_state_out_5_0_0[2:0]        ), //i
    .port_i_0_1 (keyAdd_port_state_out_5_0_1[2:0]        ), //i
    .port_i_0_2 (keyAdd_port_state_out_5_0_2[2:0]        ), //i
    .port_i_0_3 (keyAdd_port_state_out_5_0_3[2:0]        ), //i
    .port_i_0_4 (keyAdd_port_state_out_5_0_4[2:0]        ), //i
    .port_i_0_5 (keyAdd_port_state_out_5_0_5[2:0]        ), //i
    .port_i_0_6 (keyAdd_port_state_out_5_0_6[2:0]        ), //i
    .port_i_0_7 (keyAdd_port_state_out_5_0_7[2:0]        ), //i
    .port_i_1_0 (keyAdd_port_state_out_5_1_0[2:0]        ), //i
    .port_i_1_1 (keyAdd_port_state_out_5_1_1[2:0]        ), //i
    .port_i_1_2 (keyAdd_port_state_out_5_1_2[2:0]        ), //i
    .port_i_1_3 (keyAdd_port_state_out_5_1_3[2:0]        ), //i
    .port_i_1_4 (keyAdd_port_state_out_5_1_4[2:0]        ), //i
    .port_i_1_5 (keyAdd_port_state_out_5_1_5[2:0]        ), //i
    .port_i_1_6 (keyAdd_port_state_out_5_1_6[2:0]        ), //i
    .port_i_1_7 (keyAdd_port_state_out_5_1_7[2:0]        ), //i
    .port_i_2_0 (keyAdd_port_state_out_5_2_0[2:0]        ), //i
    .port_i_2_1 (keyAdd_port_state_out_5_2_1[2:0]        ), //i
    .port_i_2_2 (keyAdd_port_state_out_5_2_2[2:0]        ), //i
    .port_i_2_3 (keyAdd_port_state_out_5_2_3[2:0]        ), //i
    .port_i_2_4 (keyAdd_port_state_out_5_2_4[2:0]        ), //i
    .port_i_2_5 (keyAdd_port_state_out_5_2_5[2:0]        ), //i
    .port_i_2_6 (keyAdd_port_state_out_5_2_6[2:0]        ), //i
    .port_i_2_7 (keyAdd_port_state_out_5_2_7[2:0]        ), //i
    .port_i_3_0 (keyAdd_port_state_out_5_3_0[2:0]        ), //i
    .port_i_3_1 (keyAdd_port_state_out_5_3_1[2:0]        ), //i
    .port_i_3_2 (keyAdd_port_state_out_5_3_2[2:0]        ), //i
    .port_i_3_3 (keyAdd_port_state_out_5_3_3[2:0]        ), //i
    .port_i_3_4 (keyAdd_port_state_out_5_3_4[2:0]        ), //i
    .port_i_3_5 (keyAdd_port_state_out_5_3_5[2:0]        ), //i
    .port_i_3_6 (keyAdd_port_state_out_5_3_6[2:0]        ), //i
    .port_i_3_7 (keyAdd_port_state_out_5_3_7[2:0]        ), //i
    .port_o_0_0 (sbox_AES_BoyarPeralta_21_port_o_0_0[2:0]), //o
    .port_o_0_1 (sbox_AES_BoyarPeralta_21_port_o_0_1[2:0]), //o
    .port_o_0_2 (sbox_AES_BoyarPeralta_21_port_o_0_2[2:0]), //o
    .port_o_0_3 (sbox_AES_BoyarPeralta_21_port_o_0_3[2:0]), //o
    .port_o_0_4 (sbox_AES_BoyarPeralta_21_port_o_0_4[2:0]), //o
    .port_o_0_5 (sbox_AES_BoyarPeralta_21_port_o_0_5[2:0]), //o
    .port_o_0_6 (sbox_AES_BoyarPeralta_21_port_o_0_6[2:0]), //o
    .port_o_0_7 (sbox_AES_BoyarPeralta_21_port_o_0_7[2:0]), //o
    .port_o_1_0 (sbox_AES_BoyarPeralta_21_port_o_1_0[2:0]), //o
    .port_o_1_1 (sbox_AES_BoyarPeralta_21_port_o_1_1[2:0]), //o
    .port_o_1_2 (sbox_AES_BoyarPeralta_21_port_o_1_2[2:0]), //o
    .port_o_1_3 (sbox_AES_BoyarPeralta_21_port_o_1_3[2:0]), //o
    .port_o_1_4 (sbox_AES_BoyarPeralta_21_port_o_1_4[2:0]), //o
    .port_o_1_5 (sbox_AES_BoyarPeralta_21_port_o_1_5[2:0]), //o
    .port_o_1_6 (sbox_AES_BoyarPeralta_21_port_o_1_6[2:0]), //o
    .port_o_1_7 (sbox_AES_BoyarPeralta_21_port_o_1_7[2:0]), //o
    .port_o_2_0 (sbox_AES_BoyarPeralta_21_port_o_2_0[2:0]), //o
    .port_o_2_1 (sbox_AES_BoyarPeralta_21_port_o_2_1[2:0]), //o
    .port_o_2_2 (sbox_AES_BoyarPeralta_21_port_o_2_2[2:0]), //o
    .port_o_2_3 (sbox_AES_BoyarPeralta_21_port_o_2_3[2:0]), //o
    .port_o_2_4 (sbox_AES_BoyarPeralta_21_port_o_2_4[2:0]), //o
    .port_o_2_5 (sbox_AES_BoyarPeralta_21_port_o_2_5[2:0]), //o
    .port_o_2_6 (sbox_AES_BoyarPeralta_21_port_o_2_6[2:0]), //o
    .port_o_2_7 (sbox_AES_BoyarPeralta_21_port_o_2_7[2:0]), //o
    .port_o_3_0 (sbox_AES_BoyarPeralta_21_port_o_3_0[2:0]), //o
    .port_o_3_1 (sbox_AES_BoyarPeralta_21_port_o_3_1[2:0]), //o
    .port_o_3_2 (sbox_AES_BoyarPeralta_21_port_o_3_2[2:0]), //o
    .port_o_3_3 (sbox_AES_BoyarPeralta_21_port_o_3_3[2:0]), //o
    .port_o_3_4 (sbox_AES_BoyarPeralta_21_port_o_3_4[2:0]), //o
    .port_o_3_5 (sbox_AES_BoyarPeralta_21_port_o_3_5[2:0]), //o
    .port_o_3_6 (sbox_AES_BoyarPeralta_21_port_o_3_6[2:0]), //o
    .port_o_3_7 (sbox_AES_BoyarPeralta_21_port_o_3_7[2:0]), //o
    .clk        (clk                                     ), //i
    .reset      (reset                                   )  //i
  );
  Sbox_AES_BoyarPeralta sbox_AES_BoyarPeralta_22 (
    .port_i_0_0 (keyAdd_port_state_out_6_0_0[2:0]        ), //i
    .port_i_0_1 (keyAdd_port_state_out_6_0_1[2:0]        ), //i
    .port_i_0_2 (keyAdd_port_state_out_6_0_2[2:0]        ), //i
    .port_i_0_3 (keyAdd_port_state_out_6_0_3[2:0]        ), //i
    .port_i_0_4 (keyAdd_port_state_out_6_0_4[2:0]        ), //i
    .port_i_0_5 (keyAdd_port_state_out_6_0_5[2:0]        ), //i
    .port_i_0_6 (keyAdd_port_state_out_6_0_6[2:0]        ), //i
    .port_i_0_7 (keyAdd_port_state_out_6_0_7[2:0]        ), //i
    .port_i_1_0 (keyAdd_port_state_out_6_1_0[2:0]        ), //i
    .port_i_1_1 (keyAdd_port_state_out_6_1_1[2:0]        ), //i
    .port_i_1_2 (keyAdd_port_state_out_6_1_2[2:0]        ), //i
    .port_i_1_3 (keyAdd_port_state_out_6_1_3[2:0]        ), //i
    .port_i_1_4 (keyAdd_port_state_out_6_1_4[2:0]        ), //i
    .port_i_1_5 (keyAdd_port_state_out_6_1_5[2:0]        ), //i
    .port_i_1_6 (keyAdd_port_state_out_6_1_6[2:0]        ), //i
    .port_i_1_7 (keyAdd_port_state_out_6_1_7[2:0]        ), //i
    .port_i_2_0 (keyAdd_port_state_out_6_2_0[2:0]        ), //i
    .port_i_2_1 (keyAdd_port_state_out_6_2_1[2:0]        ), //i
    .port_i_2_2 (keyAdd_port_state_out_6_2_2[2:0]        ), //i
    .port_i_2_3 (keyAdd_port_state_out_6_2_3[2:0]        ), //i
    .port_i_2_4 (keyAdd_port_state_out_6_2_4[2:0]        ), //i
    .port_i_2_5 (keyAdd_port_state_out_6_2_5[2:0]        ), //i
    .port_i_2_6 (keyAdd_port_state_out_6_2_6[2:0]        ), //i
    .port_i_2_7 (keyAdd_port_state_out_6_2_7[2:0]        ), //i
    .port_i_3_0 (keyAdd_port_state_out_6_3_0[2:0]        ), //i
    .port_i_3_1 (keyAdd_port_state_out_6_3_1[2:0]        ), //i
    .port_i_3_2 (keyAdd_port_state_out_6_3_2[2:0]        ), //i
    .port_i_3_3 (keyAdd_port_state_out_6_3_3[2:0]        ), //i
    .port_i_3_4 (keyAdd_port_state_out_6_3_4[2:0]        ), //i
    .port_i_3_5 (keyAdd_port_state_out_6_3_5[2:0]        ), //i
    .port_i_3_6 (keyAdd_port_state_out_6_3_6[2:0]        ), //i
    .port_i_3_7 (keyAdd_port_state_out_6_3_7[2:0]        ), //i
    .port_o_0_0 (sbox_AES_BoyarPeralta_22_port_o_0_0[2:0]), //o
    .port_o_0_1 (sbox_AES_BoyarPeralta_22_port_o_0_1[2:0]), //o
    .port_o_0_2 (sbox_AES_BoyarPeralta_22_port_o_0_2[2:0]), //o
    .port_o_0_3 (sbox_AES_BoyarPeralta_22_port_o_0_3[2:0]), //o
    .port_o_0_4 (sbox_AES_BoyarPeralta_22_port_o_0_4[2:0]), //o
    .port_o_0_5 (sbox_AES_BoyarPeralta_22_port_o_0_5[2:0]), //o
    .port_o_0_6 (sbox_AES_BoyarPeralta_22_port_o_0_6[2:0]), //o
    .port_o_0_7 (sbox_AES_BoyarPeralta_22_port_o_0_7[2:0]), //o
    .port_o_1_0 (sbox_AES_BoyarPeralta_22_port_o_1_0[2:0]), //o
    .port_o_1_1 (sbox_AES_BoyarPeralta_22_port_o_1_1[2:0]), //o
    .port_o_1_2 (sbox_AES_BoyarPeralta_22_port_o_1_2[2:0]), //o
    .port_o_1_3 (sbox_AES_BoyarPeralta_22_port_o_1_3[2:0]), //o
    .port_o_1_4 (sbox_AES_BoyarPeralta_22_port_o_1_4[2:0]), //o
    .port_o_1_5 (sbox_AES_BoyarPeralta_22_port_o_1_5[2:0]), //o
    .port_o_1_6 (sbox_AES_BoyarPeralta_22_port_o_1_6[2:0]), //o
    .port_o_1_7 (sbox_AES_BoyarPeralta_22_port_o_1_7[2:0]), //o
    .port_o_2_0 (sbox_AES_BoyarPeralta_22_port_o_2_0[2:0]), //o
    .port_o_2_1 (sbox_AES_BoyarPeralta_22_port_o_2_1[2:0]), //o
    .port_o_2_2 (sbox_AES_BoyarPeralta_22_port_o_2_2[2:0]), //o
    .port_o_2_3 (sbox_AES_BoyarPeralta_22_port_o_2_3[2:0]), //o
    .port_o_2_4 (sbox_AES_BoyarPeralta_22_port_o_2_4[2:0]), //o
    .port_o_2_5 (sbox_AES_BoyarPeralta_22_port_o_2_5[2:0]), //o
    .port_o_2_6 (sbox_AES_BoyarPeralta_22_port_o_2_6[2:0]), //o
    .port_o_2_7 (sbox_AES_BoyarPeralta_22_port_o_2_7[2:0]), //o
    .port_o_3_0 (sbox_AES_BoyarPeralta_22_port_o_3_0[2:0]), //o
    .port_o_3_1 (sbox_AES_BoyarPeralta_22_port_o_3_1[2:0]), //o
    .port_o_3_2 (sbox_AES_BoyarPeralta_22_port_o_3_2[2:0]), //o
    .port_o_3_3 (sbox_AES_BoyarPeralta_22_port_o_3_3[2:0]), //o
    .port_o_3_4 (sbox_AES_BoyarPeralta_22_port_o_3_4[2:0]), //o
    .port_o_3_5 (sbox_AES_BoyarPeralta_22_port_o_3_5[2:0]), //o
    .port_o_3_6 (sbox_AES_BoyarPeralta_22_port_o_3_6[2:0]), //o
    .port_o_3_7 (sbox_AES_BoyarPeralta_22_port_o_3_7[2:0]), //o
    .clk        (clk                                     ), //i
    .reset      (reset                                   )  //i
  );
  Sbox_AES_BoyarPeralta sbox_AES_BoyarPeralta_23 (
    .port_i_0_0 (keyAdd_port_state_out_7_0_0[2:0]        ), //i
    .port_i_0_1 (keyAdd_port_state_out_7_0_1[2:0]        ), //i
    .port_i_0_2 (keyAdd_port_state_out_7_0_2[2:0]        ), //i
    .port_i_0_3 (keyAdd_port_state_out_7_0_3[2:0]        ), //i
    .port_i_0_4 (keyAdd_port_state_out_7_0_4[2:0]        ), //i
    .port_i_0_5 (keyAdd_port_state_out_7_0_5[2:0]        ), //i
    .port_i_0_6 (keyAdd_port_state_out_7_0_6[2:0]        ), //i
    .port_i_0_7 (keyAdd_port_state_out_7_0_7[2:0]        ), //i
    .port_i_1_0 (keyAdd_port_state_out_7_1_0[2:0]        ), //i
    .port_i_1_1 (keyAdd_port_state_out_7_1_1[2:0]        ), //i
    .port_i_1_2 (keyAdd_port_state_out_7_1_2[2:0]        ), //i
    .port_i_1_3 (keyAdd_port_state_out_7_1_3[2:0]        ), //i
    .port_i_1_4 (keyAdd_port_state_out_7_1_4[2:0]        ), //i
    .port_i_1_5 (keyAdd_port_state_out_7_1_5[2:0]        ), //i
    .port_i_1_6 (keyAdd_port_state_out_7_1_6[2:0]        ), //i
    .port_i_1_7 (keyAdd_port_state_out_7_1_7[2:0]        ), //i
    .port_i_2_0 (keyAdd_port_state_out_7_2_0[2:0]        ), //i
    .port_i_2_1 (keyAdd_port_state_out_7_2_1[2:0]        ), //i
    .port_i_2_2 (keyAdd_port_state_out_7_2_2[2:0]        ), //i
    .port_i_2_3 (keyAdd_port_state_out_7_2_3[2:0]        ), //i
    .port_i_2_4 (keyAdd_port_state_out_7_2_4[2:0]        ), //i
    .port_i_2_5 (keyAdd_port_state_out_7_2_5[2:0]        ), //i
    .port_i_2_6 (keyAdd_port_state_out_7_2_6[2:0]        ), //i
    .port_i_2_7 (keyAdd_port_state_out_7_2_7[2:0]        ), //i
    .port_i_3_0 (keyAdd_port_state_out_7_3_0[2:0]        ), //i
    .port_i_3_1 (keyAdd_port_state_out_7_3_1[2:0]        ), //i
    .port_i_3_2 (keyAdd_port_state_out_7_3_2[2:0]        ), //i
    .port_i_3_3 (keyAdd_port_state_out_7_3_3[2:0]        ), //i
    .port_i_3_4 (keyAdd_port_state_out_7_3_4[2:0]        ), //i
    .port_i_3_5 (keyAdd_port_state_out_7_3_5[2:0]        ), //i
    .port_i_3_6 (keyAdd_port_state_out_7_3_6[2:0]        ), //i
    .port_i_3_7 (keyAdd_port_state_out_7_3_7[2:0]        ), //i
    .port_o_0_0 (sbox_AES_BoyarPeralta_23_port_o_0_0[2:0]), //o
    .port_o_0_1 (sbox_AES_BoyarPeralta_23_port_o_0_1[2:0]), //o
    .port_o_0_2 (sbox_AES_BoyarPeralta_23_port_o_0_2[2:0]), //o
    .port_o_0_3 (sbox_AES_BoyarPeralta_23_port_o_0_3[2:0]), //o
    .port_o_0_4 (sbox_AES_BoyarPeralta_23_port_o_0_4[2:0]), //o
    .port_o_0_5 (sbox_AES_BoyarPeralta_23_port_o_0_5[2:0]), //o
    .port_o_0_6 (sbox_AES_BoyarPeralta_23_port_o_0_6[2:0]), //o
    .port_o_0_7 (sbox_AES_BoyarPeralta_23_port_o_0_7[2:0]), //o
    .port_o_1_0 (sbox_AES_BoyarPeralta_23_port_o_1_0[2:0]), //o
    .port_o_1_1 (sbox_AES_BoyarPeralta_23_port_o_1_1[2:0]), //o
    .port_o_1_2 (sbox_AES_BoyarPeralta_23_port_o_1_2[2:0]), //o
    .port_o_1_3 (sbox_AES_BoyarPeralta_23_port_o_1_3[2:0]), //o
    .port_o_1_4 (sbox_AES_BoyarPeralta_23_port_o_1_4[2:0]), //o
    .port_o_1_5 (sbox_AES_BoyarPeralta_23_port_o_1_5[2:0]), //o
    .port_o_1_6 (sbox_AES_BoyarPeralta_23_port_o_1_6[2:0]), //o
    .port_o_1_7 (sbox_AES_BoyarPeralta_23_port_o_1_7[2:0]), //o
    .port_o_2_0 (sbox_AES_BoyarPeralta_23_port_o_2_0[2:0]), //o
    .port_o_2_1 (sbox_AES_BoyarPeralta_23_port_o_2_1[2:0]), //o
    .port_o_2_2 (sbox_AES_BoyarPeralta_23_port_o_2_2[2:0]), //o
    .port_o_2_3 (sbox_AES_BoyarPeralta_23_port_o_2_3[2:0]), //o
    .port_o_2_4 (sbox_AES_BoyarPeralta_23_port_o_2_4[2:0]), //o
    .port_o_2_5 (sbox_AES_BoyarPeralta_23_port_o_2_5[2:0]), //o
    .port_o_2_6 (sbox_AES_BoyarPeralta_23_port_o_2_6[2:0]), //o
    .port_o_2_7 (sbox_AES_BoyarPeralta_23_port_o_2_7[2:0]), //o
    .port_o_3_0 (sbox_AES_BoyarPeralta_23_port_o_3_0[2:0]), //o
    .port_o_3_1 (sbox_AES_BoyarPeralta_23_port_o_3_1[2:0]), //o
    .port_o_3_2 (sbox_AES_BoyarPeralta_23_port_o_3_2[2:0]), //o
    .port_o_3_3 (sbox_AES_BoyarPeralta_23_port_o_3_3[2:0]), //o
    .port_o_3_4 (sbox_AES_BoyarPeralta_23_port_o_3_4[2:0]), //o
    .port_o_3_5 (sbox_AES_BoyarPeralta_23_port_o_3_5[2:0]), //o
    .port_o_3_6 (sbox_AES_BoyarPeralta_23_port_o_3_6[2:0]), //o
    .port_o_3_7 (sbox_AES_BoyarPeralta_23_port_o_3_7[2:0]), //o
    .clk        (clk                                     ), //i
    .reset      (reset                                   )  //i
  );
  Sbox_AES_BoyarPeralta sbox_AES_BoyarPeralta_24 (
    .port_i_0_0 (keyAdd_port_state_out_8_0_0[2:0]        ), //i
    .port_i_0_1 (keyAdd_port_state_out_8_0_1[2:0]        ), //i
    .port_i_0_2 (keyAdd_port_state_out_8_0_2[2:0]        ), //i
    .port_i_0_3 (keyAdd_port_state_out_8_0_3[2:0]        ), //i
    .port_i_0_4 (keyAdd_port_state_out_8_0_4[2:0]        ), //i
    .port_i_0_5 (keyAdd_port_state_out_8_0_5[2:0]        ), //i
    .port_i_0_6 (keyAdd_port_state_out_8_0_6[2:0]        ), //i
    .port_i_0_7 (keyAdd_port_state_out_8_0_7[2:0]        ), //i
    .port_i_1_0 (keyAdd_port_state_out_8_1_0[2:0]        ), //i
    .port_i_1_1 (keyAdd_port_state_out_8_1_1[2:0]        ), //i
    .port_i_1_2 (keyAdd_port_state_out_8_1_2[2:0]        ), //i
    .port_i_1_3 (keyAdd_port_state_out_8_1_3[2:0]        ), //i
    .port_i_1_4 (keyAdd_port_state_out_8_1_4[2:0]        ), //i
    .port_i_1_5 (keyAdd_port_state_out_8_1_5[2:0]        ), //i
    .port_i_1_6 (keyAdd_port_state_out_8_1_6[2:0]        ), //i
    .port_i_1_7 (keyAdd_port_state_out_8_1_7[2:0]        ), //i
    .port_i_2_0 (keyAdd_port_state_out_8_2_0[2:0]        ), //i
    .port_i_2_1 (keyAdd_port_state_out_8_2_1[2:0]        ), //i
    .port_i_2_2 (keyAdd_port_state_out_8_2_2[2:0]        ), //i
    .port_i_2_3 (keyAdd_port_state_out_8_2_3[2:0]        ), //i
    .port_i_2_4 (keyAdd_port_state_out_8_2_4[2:0]        ), //i
    .port_i_2_5 (keyAdd_port_state_out_8_2_5[2:0]        ), //i
    .port_i_2_6 (keyAdd_port_state_out_8_2_6[2:0]        ), //i
    .port_i_2_7 (keyAdd_port_state_out_8_2_7[2:0]        ), //i
    .port_i_3_0 (keyAdd_port_state_out_8_3_0[2:0]        ), //i
    .port_i_3_1 (keyAdd_port_state_out_8_3_1[2:0]        ), //i
    .port_i_3_2 (keyAdd_port_state_out_8_3_2[2:0]        ), //i
    .port_i_3_3 (keyAdd_port_state_out_8_3_3[2:0]        ), //i
    .port_i_3_4 (keyAdd_port_state_out_8_3_4[2:0]        ), //i
    .port_i_3_5 (keyAdd_port_state_out_8_3_5[2:0]        ), //i
    .port_i_3_6 (keyAdd_port_state_out_8_3_6[2:0]        ), //i
    .port_i_3_7 (keyAdd_port_state_out_8_3_7[2:0]        ), //i
    .port_o_0_0 (sbox_AES_BoyarPeralta_24_port_o_0_0[2:0]), //o
    .port_o_0_1 (sbox_AES_BoyarPeralta_24_port_o_0_1[2:0]), //o
    .port_o_0_2 (sbox_AES_BoyarPeralta_24_port_o_0_2[2:0]), //o
    .port_o_0_3 (sbox_AES_BoyarPeralta_24_port_o_0_3[2:0]), //o
    .port_o_0_4 (sbox_AES_BoyarPeralta_24_port_o_0_4[2:0]), //o
    .port_o_0_5 (sbox_AES_BoyarPeralta_24_port_o_0_5[2:0]), //o
    .port_o_0_6 (sbox_AES_BoyarPeralta_24_port_o_0_6[2:0]), //o
    .port_o_0_7 (sbox_AES_BoyarPeralta_24_port_o_0_7[2:0]), //o
    .port_o_1_0 (sbox_AES_BoyarPeralta_24_port_o_1_0[2:0]), //o
    .port_o_1_1 (sbox_AES_BoyarPeralta_24_port_o_1_1[2:0]), //o
    .port_o_1_2 (sbox_AES_BoyarPeralta_24_port_o_1_2[2:0]), //o
    .port_o_1_3 (sbox_AES_BoyarPeralta_24_port_o_1_3[2:0]), //o
    .port_o_1_4 (sbox_AES_BoyarPeralta_24_port_o_1_4[2:0]), //o
    .port_o_1_5 (sbox_AES_BoyarPeralta_24_port_o_1_5[2:0]), //o
    .port_o_1_6 (sbox_AES_BoyarPeralta_24_port_o_1_6[2:0]), //o
    .port_o_1_7 (sbox_AES_BoyarPeralta_24_port_o_1_7[2:0]), //o
    .port_o_2_0 (sbox_AES_BoyarPeralta_24_port_o_2_0[2:0]), //o
    .port_o_2_1 (sbox_AES_BoyarPeralta_24_port_o_2_1[2:0]), //o
    .port_o_2_2 (sbox_AES_BoyarPeralta_24_port_o_2_2[2:0]), //o
    .port_o_2_3 (sbox_AES_BoyarPeralta_24_port_o_2_3[2:0]), //o
    .port_o_2_4 (sbox_AES_BoyarPeralta_24_port_o_2_4[2:0]), //o
    .port_o_2_5 (sbox_AES_BoyarPeralta_24_port_o_2_5[2:0]), //o
    .port_o_2_6 (sbox_AES_BoyarPeralta_24_port_o_2_6[2:0]), //o
    .port_o_2_7 (sbox_AES_BoyarPeralta_24_port_o_2_7[2:0]), //o
    .port_o_3_0 (sbox_AES_BoyarPeralta_24_port_o_3_0[2:0]), //o
    .port_o_3_1 (sbox_AES_BoyarPeralta_24_port_o_3_1[2:0]), //o
    .port_o_3_2 (sbox_AES_BoyarPeralta_24_port_o_3_2[2:0]), //o
    .port_o_3_3 (sbox_AES_BoyarPeralta_24_port_o_3_3[2:0]), //o
    .port_o_3_4 (sbox_AES_BoyarPeralta_24_port_o_3_4[2:0]), //o
    .port_o_3_5 (sbox_AES_BoyarPeralta_24_port_o_3_5[2:0]), //o
    .port_o_3_6 (sbox_AES_BoyarPeralta_24_port_o_3_6[2:0]), //o
    .port_o_3_7 (sbox_AES_BoyarPeralta_24_port_o_3_7[2:0]), //o
    .clk        (clk                                     ), //i
    .reset      (reset                                   )  //i
  );
  Sbox_AES_BoyarPeralta sbox_AES_BoyarPeralta_25 (
    .port_i_0_0 (keyAdd_port_state_out_9_0_0[2:0]        ), //i
    .port_i_0_1 (keyAdd_port_state_out_9_0_1[2:0]        ), //i
    .port_i_0_2 (keyAdd_port_state_out_9_0_2[2:0]        ), //i
    .port_i_0_3 (keyAdd_port_state_out_9_0_3[2:0]        ), //i
    .port_i_0_4 (keyAdd_port_state_out_9_0_4[2:0]        ), //i
    .port_i_0_5 (keyAdd_port_state_out_9_0_5[2:0]        ), //i
    .port_i_0_6 (keyAdd_port_state_out_9_0_6[2:0]        ), //i
    .port_i_0_7 (keyAdd_port_state_out_9_0_7[2:0]        ), //i
    .port_i_1_0 (keyAdd_port_state_out_9_1_0[2:0]        ), //i
    .port_i_1_1 (keyAdd_port_state_out_9_1_1[2:0]        ), //i
    .port_i_1_2 (keyAdd_port_state_out_9_1_2[2:0]        ), //i
    .port_i_1_3 (keyAdd_port_state_out_9_1_3[2:0]        ), //i
    .port_i_1_4 (keyAdd_port_state_out_9_1_4[2:0]        ), //i
    .port_i_1_5 (keyAdd_port_state_out_9_1_5[2:0]        ), //i
    .port_i_1_6 (keyAdd_port_state_out_9_1_6[2:0]        ), //i
    .port_i_1_7 (keyAdd_port_state_out_9_1_7[2:0]        ), //i
    .port_i_2_0 (keyAdd_port_state_out_9_2_0[2:0]        ), //i
    .port_i_2_1 (keyAdd_port_state_out_9_2_1[2:0]        ), //i
    .port_i_2_2 (keyAdd_port_state_out_9_2_2[2:0]        ), //i
    .port_i_2_3 (keyAdd_port_state_out_9_2_3[2:0]        ), //i
    .port_i_2_4 (keyAdd_port_state_out_9_2_4[2:0]        ), //i
    .port_i_2_5 (keyAdd_port_state_out_9_2_5[2:0]        ), //i
    .port_i_2_6 (keyAdd_port_state_out_9_2_6[2:0]        ), //i
    .port_i_2_7 (keyAdd_port_state_out_9_2_7[2:0]        ), //i
    .port_i_3_0 (keyAdd_port_state_out_9_3_0[2:0]        ), //i
    .port_i_3_1 (keyAdd_port_state_out_9_3_1[2:0]        ), //i
    .port_i_3_2 (keyAdd_port_state_out_9_3_2[2:0]        ), //i
    .port_i_3_3 (keyAdd_port_state_out_9_3_3[2:0]        ), //i
    .port_i_3_4 (keyAdd_port_state_out_9_3_4[2:0]        ), //i
    .port_i_3_5 (keyAdd_port_state_out_9_3_5[2:0]        ), //i
    .port_i_3_6 (keyAdd_port_state_out_9_3_6[2:0]        ), //i
    .port_i_3_7 (keyAdd_port_state_out_9_3_7[2:0]        ), //i
    .port_o_0_0 (sbox_AES_BoyarPeralta_25_port_o_0_0[2:0]), //o
    .port_o_0_1 (sbox_AES_BoyarPeralta_25_port_o_0_1[2:0]), //o
    .port_o_0_2 (sbox_AES_BoyarPeralta_25_port_o_0_2[2:0]), //o
    .port_o_0_3 (sbox_AES_BoyarPeralta_25_port_o_0_3[2:0]), //o
    .port_o_0_4 (sbox_AES_BoyarPeralta_25_port_o_0_4[2:0]), //o
    .port_o_0_5 (sbox_AES_BoyarPeralta_25_port_o_0_5[2:0]), //o
    .port_o_0_6 (sbox_AES_BoyarPeralta_25_port_o_0_6[2:0]), //o
    .port_o_0_7 (sbox_AES_BoyarPeralta_25_port_o_0_7[2:0]), //o
    .port_o_1_0 (sbox_AES_BoyarPeralta_25_port_o_1_0[2:0]), //o
    .port_o_1_1 (sbox_AES_BoyarPeralta_25_port_o_1_1[2:0]), //o
    .port_o_1_2 (sbox_AES_BoyarPeralta_25_port_o_1_2[2:0]), //o
    .port_o_1_3 (sbox_AES_BoyarPeralta_25_port_o_1_3[2:0]), //o
    .port_o_1_4 (sbox_AES_BoyarPeralta_25_port_o_1_4[2:0]), //o
    .port_o_1_5 (sbox_AES_BoyarPeralta_25_port_o_1_5[2:0]), //o
    .port_o_1_6 (sbox_AES_BoyarPeralta_25_port_o_1_6[2:0]), //o
    .port_o_1_7 (sbox_AES_BoyarPeralta_25_port_o_1_7[2:0]), //o
    .port_o_2_0 (sbox_AES_BoyarPeralta_25_port_o_2_0[2:0]), //o
    .port_o_2_1 (sbox_AES_BoyarPeralta_25_port_o_2_1[2:0]), //o
    .port_o_2_2 (sbox_AES_BoyarPeralta_25_port_o_2_2[2:0]), //o
    .port_o_2_3 (sbox_AES_BoyarPeralta_25_port_o_2_3[2:0]), //o
    .port_o_2_4 (sbox_AES_BoyarPeralta_25_port_o_2_4[2:0]), //o
    .port_o_2_5 (sbox_AES_BoyarPeralta_25_port_o_2_5[2:0]), //o
    .port_o_2_6 (sbox_AES_BoyarPeralta_25_port_o_2_6[2:0]), //o
    .port_o_2_7 (sbox_AES_BoyarPeralta_25_port_o_2_7[2:0]), //o
    .port_o_3_0 (sbox_AES_BoyarPeralta_25_port_o_3_0[2:0]), //o
    .port_o_3_1 (sbox_AES_BoyarPeralta_25_port_o_3_1[2:0]), //o
    .port_o_3_2 (sbox_AES_BoyarPeralta_25_port_o_3_2[2:0]), //o
    .port_o_3_3 (sbox_AES_BoyarPeralta_25_port_o_3_3[2:0]), //o
    .port_o_3_4 (sbox_AES_BoyarPeralta_25_port_o_3_4[2:0]), //o
    .port_o_3_5 (sbox_AES_BoyarPeralta_25_port_o_3_5[2:0]), //o
    .port_o_3_6 (sbox_AES_BoyarPeralta_25_port_o_3_6[2:0]), //o
    .port_o_3_7 (sbox_AES_BoyarPeralta_25_port_o_3_7[2:0]), //o
    .clk        (clk                                     ), //i
    .reset      (reset                                   )  //i
  );
  Sbox_AES_BoyarPeralta sbox_AES_BoyarPeralta_26 (
    .port_i_0_0 (keyAdd_port_state_out_10_0_0[2:0]       ), //i
    .port_i_0_1 (keyAdd_port_state_out_10_0_1[2:0]       ), //i
    .port_i_0_2 (keyAdd_port_state_out_10_0_2[2:0]       ), //i
    .port_i_0_3 (keyAdd_port_state_out_10_0_3[2:0]       ), //i
    .port_i_0_4 (keyAdd_port_state_out_10_0_4[2:0]       ), //i
    .port_i_0_5 (keyAdd_port_state_out_10_0_5[2:0]       ), //i
    .port_i_0_6 (keyAdd_port_state_out_10_0_6[2:0]       ), //i
    .port_i_0_7 (keyAdd_port_state_out_10_0_7[2:0]       ), //i
    .port_i_1_0 (keyAdd_port_state_out_10_1_0[2:0]       ), //i
    .port_i_1_1 (keyAdd_port_state_out_10_1_1[2:0]       ), //i
    .port_i_1_2 (keyAdd_port_state_out_10_1_2[2:0]       ), //i
    .port_i_1_3 (keyAdd_port_state_out_10_1_3[2:0]       ), //i
    .port_i_1_4 (keyAdd_port_state_out_10_1_4[2:0]       ), //i
    .port_i_1_5 (keyAdd_port_state_out_10_1_5[2:0]       ), //i
    .port_i_1_6 (keyAdd_port_state_out_10_1_6[2:0]       ), //i
    .port_i_1_7 (keyAdd_port_state_out_10_1_7[2:0]       ), //i
    .port_i_2_0 (keyAdd_port_state_out_10_2_0[2:0]       ), //i
    .port_i_2_1 (keyAdd_port_state_out_10_2_1[2:0]       ), //i
    .port_i_2_2 (keyAdd_port_state_out_10_2_2[2:0]       ), //i
    .port_i_2_3 (keyAdd_port_state_out_10_2_3[2:0]       ), //i
    .port_i_2_4 (keyAdd_port_state_out_10_2_4[2:0]       ), //i
    .port_i_2_5 (keyAdd_port_state_out_10_2_5[2:0]       ), //i
    .port_i_2_6 (keyAdd_port_state_out_10_2_6[2:0]       ), //i
    .port_i_2_7 (keyAdd_port_state_out_10_2_7[2:0]       ), //i
    .port_i_3_0 (keyAdd_port_state_out_10_3_0[2:0]       ), //i
    .port_i_3_1 (keyAdd_port_state_out_10_3_1[2:0]       ), //i
    .port_i_3_2 (keyAdd_port_state_out_10_3_2[2:0]       ), //i
    .port_i_3_3 (keyAdd_port_state_out_10_3_3[2:0]       ), //i
    .port_i_3_4 (keyAdd_port_state_out_10_3_4[2:0]       ), //i
    .port_i_3_5 (keyAdd_port_state_out_10_3_5[2:0]       ), //i
    .port_i_3_6 (keyAdd_port_state_out_10_3_6[2:0]       ), //i
    .port_i_3_7 (keyAdd_port_state_out_10_3_7[2:0]       ), //i
    .port_o_0_0 (sbox_AES_BoyarPeralta_26_port_o_0_0[2:0]), //o
    .port_o_0_1 (sbox_AES_BoyarPeralta_26_port_o_0_1[2:0]), //o
    .port_o_0_2 (sbox_AES_BoyarPeralta_26_port_o_0_2[2:0]), //o
    .port_o_0_3 (sbox_AES_BoyarPeralta_26_port_o_0_3[2:0]), //o
    .port_o_0_4 (sbox_AES_BoyarPeralta_26_port_o_0_4[2:0]), //o
    .port_o_0_5 (sbox_AES_BoyarPeralta_26_port_o_0_5[2:0]), //o
    .port_o_0_6 (sbox_AES_BoyarPeralta_26_port_o_0_6[2:0]), //o
    .port_o_0_7 (sbox_AES_BoyarPeralta_26_port_o_0_7[2:0]), //o
    .port_o_1_0 (sbox_AES_BoyarPeralta_26_port_o_1_0[2:0]), //o
    .port_o_1_1 (sbox_AES_BoyarPeralta_26_port_o_1_1[2:0]), //o
    .port_o_1_2 (sbox_AES_BoyarPeralta_26_port_o_1_2[2:0]), //o
    .port_o_1_3 (sbox_AES_BoyarPeralta_26_port_o_1_3[2:0]), //o
    .port_o_1_4 (sbox_AES_BoyarPeralta_26_port_o_1_4[2:0]), //o
    .port_o_1_5 (sbox_AES_BoyarPeralta_26_port_o_1_5[2:0]), //o
    .port_o_1_6 (sbox_AES_BoyarPeralta_26_port_o_1_6[2:0]), //o
    .port_o_1_7 (sbox_AES_BoyarPeralta_26_port_o_1_7[2:0]), //o
    .port_o_2_0 (sbox_AES_BoyarPeralta_26_port_o_2_0[2:0]), //o
    .port_o_2_1 (sbox_AES_BoyarPeralta_26_port_o_2_1[2:0]), //o
    .port_o_2_2 (sbox_AES_BoyarPeralta_26_port_o_2_2[2:0]), //o
    .port_o_2_3 (sbox_AES_BoyarPeralta_26_port_o_2_3[2:0]), //o
    .port_o_2_4 (sbox_AES_BoyarPeralta_26_port_o_2_4[2:0]), //o
    .port_o_2_5 (sbox_AES_BoyarPeralta_26_port_o_2_5[2:0]), //o
    .port_o_2_6 (sbox_AES_BoyarPeralta_26_port_o_2_6[2:0]), //o
    .port_o_2_7 (sbox_AES_BoyarPeralta_26_port_o_2_7[2:0]), //o
    .port_o_3_0 (sbox_AES_BoyarPeralta_26_port_o_3_0[2:0]), //o
    .port_o_3_1 (sbox_AES_BoyarPeralta_26_port_o_3_1[2:0]), //o
    .port_o_3_2 (sbox_AES_BoyarPeralta_26_port_o_3_2[2:0]), //o
    .port_o_3_3 (sbox_AES_BoyarPeralta_26_port_o_3_3[2:0]), //o
    .port_o_3_4 (sbox_AES_BoyarPeralta_26_port_o_3_4[2:0]), //o
    .port_o_3_5 (sbox_AES_BoyarPeralta_26_port_o_3_5[2:0]), //o
    .port_o_3_6 (sbox_AES_BoyarPeralta_26_port_o_3_6[2:0]), //o
    .port_o_3_7 (sbox_AES_BoyarPeralta_26_port_o_3_7[2:0]), //o
    .clk        (clk                                     ), //i
    .reset      (reset                                   )  //i
  );
  Sbox_AES_BoyarPeralta sbox_AES_BoyarPeralta_27 (
    .port_i_0_0 (keyAdd_port_state_out_11_0_0[2:0]       ), //i
    .port_i_0_1 (keyAdd_port_state_out_11_0_1[2:0]       ), //i
    .port_i_0_2 (keyAdd_port_state_out_11_0_2[2:0]       ), //i
    .port_i_0_3 (keyAdd_port_state_out_11_0_3[2:0]       ), //i
    .port_i_0_4 (keyAdd_port_state_out_11_0_4[2:0]       ), //i
    .port_i_0_5 (keyAdd_port_state_out_11_0_5[2:0]       ), //i
    .port_i_0_6 (keyAdd_port_state_out_11_0_6[2:0]       ), //i
    .port_i_0_7 (keyAdd_port_state_out_11_0_7[2:0]       ), //i
    .port_i_1_0 (keyAdd_port_state_out_11_1_0[2:0]       ), //i
    .port_i_1_1 (keyAdd_port_state_out_11_1_1[2:0]       ), //i
    .port_i_1_2 (keyAdd_port_state_out_11_1_2[2:0]       ), //i
    .port_i_1_3 (keyAdd_port_state_out_11_1_3[2:0]       ), //i
    .port_i_1_4 (keyAdd_port_state_out_11_1_4[2:0]       ), //i
    .port_i_1_5 (keyAdd_port_state_out_11_1_5[2:0]       ), //i
    .port_i_1_6 (keyAdd_port_state_out_11_1_6[2:0]       ), //i
    .port_i_1_7 (keyAdd_port_state_out_11_1_7[2:0]       ), //i
    .port_i_2_0 (keyAdd_port_state_out_11_2_0[2:0]       ), //i
    .port_i_2_1 (keyAdd_port_state_out_11_2_1[2:0]       ), //i
    .port_i_2_2 (keyAdd_port_state_out_11_2_2[2:0]       ), //i
    .port_i_2_3 (keyAdd_port_state_out_11_2_3[2:0]       ), //i
    .port_i_2_4 (keyAdd_port_state_out_11_2_4[2:0]       ), //i
    .port_i_2_5 (keyAdd_port_state_out_11_2_5[2:0]       ), //i
    .port_i_2_6 (keyAdd_port_state_out_11_2_6[2:0]       ), //i
    .port_i_2_7 (keyAdd_port_state_out_11_2_7[2:0]       ), //i
    .port_i_3_0 (keyAdd_port_state_out_11_3_0[2:0]       ), //i
    .port_i_3_1 (keyAdd_port_state_out_11_3_1[2:0]       ), //i
    .port_i_3_2 (keyAdd_port_state_out_11_3_2[2:0]       ), //i
    .port_i_3_3 (keyAdd_port_state_out_11_3_3[2:0]       ), //i
    .port_i_3_4 (keyAdd_port_state_out_11_3_4[2:0]       ), //i
    .port_i_3_5 (keyAdd_port_state_out_11_3_5[2:0]       ), //i
    .port_i_3_6 (keyAdd_port_state_out_11_3_6[2:0]       ), //i
    .port_i_3_7 (keyAdd_port_state_out_11_3_7[2:0]       ), //i
    .port_o_0_0 (sbox_AES_BoyarPeralta_27_port_o_0_0[2:0]), //o
    .port_o_0_1 (sbox_AES_BoyarPeralta_27_port_o_0_1[2:0]), //o
    .port_o_0_2 (sbox_AES_BoyarPeralta_27_port_o_0_2[2:0]), //o
    .port_o_0_3 (sbox_AES_BoyarPeralta_27_port_o_0_3[2:0]), //o
    .port_o_0_4 (sbox_AES_BoyarPeralta_27_port_o_0_4[2:0]), //o
    .port_o_0_5 (sbox_AES_BoyarPeralta_27_port_o_0_5[2:0]), //o
    .port_o_0_6 (sbox_AES_BoyarPeralta_27_port_o_0_6[2:0]), //o
    .port_o_0_7 (sbox_AES_BoyarPeralta_27_port_o_0_7[2:0]), //o
    .port_o_1_0 (sbox_AES_BoyarPeralta_27_port_o_1_0[2:0]), //o
    .port_o_1_1 (sbox_AES_BoyarPeralta_27_port_o_1_1[2:0]), //o
    .port_o_1_2 (sbox_AES_BoyarPeralta_27_port_o_1_2[2:0]), //o
    .port_o_1_3 (sbox_AES_BoyarPeralta_27_port_o_1_3[2:0]), //o
    .port_o_1_4 (sbox_AES_BoyarPeralta_27_port_o_1_4[2:0]), //o
    .port_o_1_5 (sbox_AES_BoyarPeralta_27_port_o_1_5[2:0]), //o
    .port_o_1_6 (sbox_AES_BoyarPeralta_27_port_o_1_6[2:0]), //o
    .port_o_1_7 (sbox_AES_BoyarPeralta_27_port_o_1_7[2:0]), //o
    .port_o_2_0 (sbox_AES_BoyarPeralta_27_port_o_2_0[2:0]), //o
    .port_o_2_1 (sbox_AES_BoyarPeralta_27_port_o_2_1[2:0]), //o
    .port_o_2_2 (sbox_AES_BoyarPeralta_27_port_o_2_2[2:0]), //o
    .port_o_2_3 (sbox_AES_BoyarPeralta_27_port_o_2_3[2:0]), //o
    .port_o_2_4 (sbox_AES_BoyarPeralta_27_port_o_2_4[2:0]), //o
    .port_o_2_5 (sbox_AES_BoyarPeralta_27_port_o_2_5[2:0]), //o
    .port_o_2_6 (sbox_AES_BoyarPeralta_27_port_o_2_6[2:0]), //o
    .port_o_2_7 (sbox_AES_BoyarPeralta_27_port_o_2_7[2:0]), //o
    .port_o_3_0 (sbox_AES_BoyarPeralta_27_port_o_3_0[2:0]), //o
    .port_o_3_1 (sbox_AES_BoyarPeralta_27_port_o_3_1[2:0]), //o
    .port_o_3_2 (sbox_AES_BoyarPeralta_27_port_o_3_2[2:0]), //o
    .port_o_3_3 (sbox_AES_BoyarPeralta_27_port_o_3_3[2:0]), //o
    .port_o_3_4 (sbox_AES_BoyarPeralta_27_port_o_3_4[2:0]), //o
    .port_o_3_5 (sbox_AES_BoyarPeralta_27_port_o_3_5[2:0]), //o
    .port_o_3_6 (sbox_AES_BoyarPeralta_27_port_o_3_6[2:0]), //o
    .port_o_3_7 (sbox_AES_BoyarPeralta_27_port_o_3_7[2:0]), //o
    .clk        (clk                                     ), //i
    .reset      (reset                                   )  //i
  );
  Sbox_AES_BoyarPeralta sbox_AES_BoyarPeralta_28 (
    .port_i_0_0 (keyAdd_port_state_out_12_0_0[2:0]       ), //i
    .port_i_0_1 (keyAdd_port_state_out_12_0_1[2:0]       ), //i
    .port_i_0_2 (keyAdd_port_state_out_12_0_2[2:0]       ), //i
    .port_i_0_3 (keyAdd_port_state_out_12_0_3[2:0]       ), //i
    .port_i_0_4 (keyAdd_port_state_out_12_0_4[2:0]       ), //i
    .port_i_0_5 (keyAdd_port_state_out_12_0_5[2:0]       ), //i
    .port_i_0_6 (keyAdd_port_state_out_12_0_6[2:0]       ), //i
    .port_i_0_7 (keyAdd_port_state_out_12_0_7[2:0]       ), //i
    .port_i_1_0 (keyAdd_port_state_out_12_1_0[2:0]       ), //i
    .port_i_1_1 (keyAdd_port_state_out_12_1_1[2:0]       ), //i
    .port_i_1_2 (keyAdd_port_state_out_12_1_2[2:0]       ), //i
    .port_i_1_3 (keyAdd_port_state_out_12_1_3[2:0]       ), //i
    .port_i_1_4 (keyAdd_port_state_out_12_1_4[2:0]       ), //i
    .port_i_1_5 (keyAdd_port_state_out_12_1_5[2:0]       ), //i
    .port_i_1_6 (keyAdd_port_state_out_12_1_6[2:0]       ), //i
    .port_i_1_7 (keyAdd_port_state_out_12_1_7[2:0]       ), //i
    .port_i_2_0 (keyAdd_port_state_out_12_2_0[2:0]       ), //i
    .port_i_2_1 (keyAdd_port_state_out_12_2_1[2:0]       ), //i
    .port_i_2_2 (keyAdd_port_state_out_12_2_2[2:0]       ), //i
    .port_i_2_3 (keyAdd_port_state_out_12_2_3[2:0]       ), //i
    .port_i_2_4 (keyAdd_port_state_out_12_2_4[2:0]       ), //i
    .port_i_2_5 (keyAdd_port_state_out_12_2_5[2:0]       ), //i
    .port_i_2_6 (keyAdd_port_state_out_12_2_6[2:0]       ), //i
    .port_i_2_7 (keyAdd_port_state_out_12_2_7[2:0]       ), //i
    .port_i_3_0 (keyAdd_port_state_out_12_3_0[2:0]       ), //i
    .port_i_3_1 (keyAdd_port_state_out_12_3_1[2:0]       ), //i
    .port_i_3_2 (keyAdd_port_state_out_12_3_2[2:0]       ), //i
    .port_i_3_3 (keyAdd_port_state_out_12_3_3[2:0]       ), //i
    .port_i_3_4 (keyAdd_port_state_out_12_3_4[2:0]       ), //i
    .port_i_3_5 (keyAdd_port_state_out_12_3_5[2:0]       ), //i
    .port_i_3_6 (keyAdd_port_state_out_12_3_6[2:0]       ), //i
    .port_i_3_7 (keyAdd_port_state_out_12_3_7[2:0]       ), //i
    .port_o_0_0 (sbox_AES_BoyarPeralta_28_port_o_0_0[2:0]), //o
    .port_o_0_1 (sbox_AES_BoyarPeralta_28_port_o_0_1[2:0]), //o
    .port_o_0_2 (sbox_AES_BoyarPeralta_28_port_o_0_2[2:0]), //o
    .port_o_0_3 (sbox_AES_BoyarPeralta_28_port_o_0_3[2:0]), //o
    .port_o_0_4 (sbox_AES_BoyarPeralta_28_port_o_0_4[2:0]), //o
    .port_o_0_5 (sbox_AES_BoyarPeralta_28_port_o_0_5[2:0]), //o
    .port_o_0_6 (sbox_AES_BoyarPeralta_28_port_o_0_6[2:0]), //o
    .port_o_0_7 (sbox_AES_BoyarPeralta_28_port_o_0_7[2:0]), //o
    .port_o_1_0 (sbox_AES_BoyarPeralta_28_port_o_1_0[2:0]), //o
    .port_o_1_1 (sbox_AES_BoyarPeralta_28_port_o_1_1[2:0]), //o
    .port_o_1_2 (sbox_AES_BoyarPeralta_28_port_o_1_2[2:0]), //o
    .port_o_1_3 (sbox_AES_BoyarPeralta_28_port_o_1_3[2:0]), //o
    .port_o_1_4 (sbox_AES_BoyarPeralta_28_port_o_1_4[2:0]), //o
    .port_o_1_5 (sbox_AES_BoyarPeralta_28_port_o_1_5[2:0]), //o
    .port_o_1_6 (sbox_AES_BoyarPeralta_28_port_o_1_6[2:0]), //o
    .port_o_1_7 (sbox_AES_BoyarPeralta_28_port_o_1_7[2:0]), //o
    .port_o_2_0 (sbox_AES_BoyarPeralta_28_port_o_2_0[2:0]), //o
    .port_o_2_1 (sbox_AES_BoyarPeralta_28_port_o_2_1[2:0]), //o
    .port_o_2_2 (sbox_AES_BoyarPeralta_28_port_o_2_2[2:0]), //o
    .port_o_2_3 (sbox_AES_BoyarPeralta_28_port_o_2_3[2:0]), //o
    .port_o_2_4 (sbox_AES_BoyarPeralta_28_port_o_2_4[2:0]), //o
    .port_o_2_5 (sbox_AES_BoyarPeralta_28_port_o_2_5[2:0]), //o
    .port_o_2_6 (sbox_AES_BoyarPeralta_28_port_o_2_6[2:0]), //o
    .port_o_2_7 (sbox_AES_BoyarPeralta_28_port_o_2_7[2:0]), //o
    .port_o_3_0 (sbox_AES_BoyarPeralta_28_port_o_3_0[2:0]), //o
    .port_o_3_1 (sbox_AES_BoyarPeralta_28_port_o_3_1[2:0]), //o
    .port_o_3_2 (sbox_AES_BoyarPeralta_28_port_o_3_2[2:0]), //o
    .port_o_3_3 (sbox_AES_BoyarPeralta_28_port_o_3_3[2:0]), //o
    .port_o_3_4 (sbox_AES_BoyarPeralta_28_port_o_3_4[2:0]), //o
    .port_o_3_5 (sbox_AES_BoyarPeralta_28_port_o_3_5[2:0]), //o
    .port_o_3_6 (sbox_AES_BoyarPeralta_28_port_o_3_6[2:0]), //o
    .port_o_3_7 (sbox_AES_BoyarPeralta_28_port_o_3_7[2:0]), //o
    .clk        (clk                                     ), //i
    .reset      (reset                                   )  //i
  );
  Sbox_AES_BoyarPeralta sbox_AES_BoyarPeralta_29 (
    .port_i_0_0 (keyAdd_port_state_out_13_0_0[2:0]       ), //i
    .port_i_0_1 (keyAdd_port_state_out_13_0_1[2:0]       ), //i
    .port_i_0_2 (keyAdd_port_state_out_13_0_2[2:0]       ), //i
    .port_i_0_3 (keyAdd_port_state_out_13_0_3[2:0]       ), //i
    .port_i_0_4 (keyAdd_port_state_out_13_0_4[2:0]       ), //i
    .port_i_0_5 (keyAdd_port_state_out_13_0_5[2:0]       ), //i
    .port_i_0_6 (keyAdd_port_state_out_13_0_6[2:0]       ), //i
    .port_i_0_7 (keyAdd_port_state_out_13_0_7[2:0]       ), //i
    .port_i_1_0 (keyAdd_port_state_out_13_1_0[2:0]       ), //i
    .port_i_1_1 (keyAdd_port_state_out_13_1_1[2:0]       ), //i
    .port_i_1_2 (keyAdd_port_state_out_13_1_2[2:0]       ), //i
    .port_i_1_3 (keyAdd_port_state_out_13_1_3[2:0]       ), //i
    .port_i_1_4 (keyAdd_port_state_out_13_1_4[2:0]       ), //i
    .port_i_1_5 (keyAdd_port_state_out_13_1_5[2:0]       ), //i
    .port_i_1_6 (keyAdd_port_state_out_13_1_6[2:0]       ), //i
    .port_i_1_7 (keyAdd_port_state_out_13_1_7[2:0]       ), //i
    .port_i_2_0 (keyAdd_port_state_out_13_2_0[2:0]       ), //i
    .port_i_2_1 (keyAdd_port_state_out_13_2_1[2:0]       ), //i
    .port_i_2_2 (keyAdd_port_state_out_13_2_2[2:0]       ), //i
    .port_i_2_3 (keyAdd_port_state_out_13_2_3[2:0]       ), //i
    .port_i_2_4 (keyAdd_port_state_out_13_2_4[2:0]       ), //i
    .port_i_2_5 (keyAdd_port_state_out_13_2_5[2:0]       ), //i
    .port_i_2_6 (keyAdd_port_state_out_13_2_6[2:0]       ), //i
    .port_i_2_7 (keyAdd_port_state_out_13_2_7[2:0]       ), //i
    .port_i_3_0 (keyAdd_port_state_out_13_3_0[2:0]       ), //i
    .port_i_3_1 (keyAdd_port_state_out_13_3_1[2:0]       ), //i
    .port_i_3_2 (keyAdd_port_state_out_13_3_2[2:0]       ), //i
    .port_i_3_3 (keyAdd_port_state_out_13_3_3[2:0]       ), //i
    .port_i_3_4 (keyAdd_port_state_out_13_3_4[2:0]       ), //i
    .port_i_3_5 (keyAdd_port_state_out_13_3_5[2:0]       ), //i
    .port_i_3_6 (keyAdd_port_state_out_13_3_6[2:0]       ), //i
    .port_i_3_7 (keyAdd_port_state_out_13_3_7[2:0]       ), //i
    .port_o_0_0 (sbox_AES_BoyarPeralta_29_port_o_0_0[2:0]), //o
    .port_o_0_1 (sbox_AES_BoyarPeralta_29_port_o_0_1[2:0]), //o
    .port_o_0_2 (sbox_AES_BoyarPeralta_29_port_o_0_2[2:0]), //o
    .port_o_0_3 (sbox_AES_BoyarPeralta_29_port_o_0_3[2:0]), //o
    .port_o_0_4 (sbox_AES_BoyarPeralta_29_port_o_0_4[2:0]), //o
    .port_o_0_5 (sbox_AES_BoyarPeralta_29_port_o_0_5[2:0]), //o
    .port_o_0_6 (sbox_AES_BoyarPeralta_29_port_o_0_6[2:0]), //o
    .port_o_0_7 (sbox_AES_BoyarPeralta_29_port_o_0_7[2:0]), //o
    .port_o_1_0 (sbox_AES_BoyarPeralta_29_port_o_1_0[2:0]), //o
    .port_o_1_1 (sbox_AES_BoyarPeralta_29_port_o_1_1[2:0]), //o
    .port_o_1_2 (sbox_AES_BoyarPeralta_29_port_o_1_2[2:0]), //o
    .port_o_1_3 (sbox_AES_BoyarPeralta_29_port_o_1_3[2:0]), //o
    .port_o_1_4 (sbox_AES_BoyarPeralta_29_port_o_1_4[2:0]), //o
    .port_o_1_5 (sbox_AES_BoyarPeralta_29_port_o_1_5[2:0]), //o
    .port_o_1_6 (sbox_AES_BoyarPeralta_29_port_o_1_6[2:0]), //o
    .port_o_1_7 (sbox_AES_BoyarPeralta_29_port_o_1_7[2:0]), //o
    .port_o_2_0 (sbox_AES_BoyarPeralta_29_port_o_2_0[2:0]), //o
    .port_o_2_1 (sbox_AES_BoyarPeralta_29_port_o_2_1[2:0]), //o
    .port_o_2_2 (sbox_AES_BoyarPeralta_29_port_o_2_2[2:0]), //o
    .port_o_2_3 (sbox_AES_BoyarPeralta_29_port_o_2_3[2:0]), //o
    .port_o_2_4 (sbox_AES_BoyarPeralta_29_port_o_2_4[2:0]), //o
    .port_o_2_5 (sbox_AES_BoyarPeralta_29_port_o_2_5[2:0]), //o
    .port_o_2_6 (sbox_AES_BoyarPeralta_29_port_o_2_6[2:0]), //o
    .port_o_2_7 (sbox_AES_BoyarPeralta_29_port_o_2_7[2:0]), //o
    .port_o_3_0 (sbox_AES_BoyarPeralta_29_port_o_3_0[2:0]), //o
    .port_o_3_1 (sbox_AES_BoyarPeralta_29_port_o_3_1[2:0]), //o
    .port_o_3_2 (sbox_AES_BoyarPeralta_29_port_o_3_2[2:0]), //o
    .port_o_3_3 (sbox_AES_BoyarPeralta_29_port_o_3_3[2:0]), //o
    .port_o_3_4 (sbox_AES_BoyarPeralta_29_port_o_3_4[2:0]), //o
    .port_o_3_5 (sbox_AES_BoyarPeralta_29_port_o_3_5[2:0]), //o
    .port_o_3_6 (sbox_AES_BoyarPeralta_29_port_o_3_6[2:0]), //o
    .port_o_3_7 (sbox_AES_BoyarPeralta_29_port_o_3_7[2:0]), //o
    .clk        (clk                                     ), //i
    .reset      (reset                                   )  //i
  );
  Sbox_AES_BoyarPeralta sbox_AES_BoyarPeralta_30 (
    .port_i_0_0 (keyAdd_port_state_out_14_0_0[2:0]       ), //i
    .port_i_0_1 (keyAdd_port_state_out_14_0_1[2:0]       ), //i
    .port_i_0_2 (keyAdd_port_state_out_14_0_2[2:0]       ), //i
    .port_i_0_3 (keyAdd_port_state_out_14_0_3[2:0]       ), //i
    .port_i_0_4 (keyAdd_port_state_out_14_0_4[2:0]       ), //i
    .port_i_0_5 (keyAdd_port_state_out_14_0_5[2:0]       ), //i
    .port_i_0_6 (keyAdd_port_state_out_14_0_6[2:0]       ), //i
    .port_i_0_7 (keyAdd_port_state_out_14_0_7[2:0]       ), //i
    .port_i_1_0 (keyAdd_port_state_out_14_1_0[2:0]       ), //i
    .port_i_1_1 (keyAdd_port_state_out_14_1_1[2:0]       ), //i
    .port_i_1_2 (keyAdd_port_state_out_14_1_2[2:0]       ), //i
    .port_i_1_3 (keyAdd_port_state_out_14_1_3[2:0]       ), //i
    .port_i_1_4 (keyAdd_port_state_out_14_1_4[2:0]       ), //i
    .port_i_1_5 (keyAdd_port_state_out_14_1_5[2:0]       ), //i
    .port_i_1_6 (keyAdd_port_state_out_14_1_6[2:0]       ), //i
    .port_i_1_7 (keyAdd_port_state_out_14_1_7[2:0]       ), //i
    .port_i_2_0 (keyAdd_port_state_out_14_2_0[2:0]       ), //i
    .port_i_2_1 (keyAdd_port_state_out_14_2_1[2:0]       ), //i
    .port_i_2_2 (keyAdd_port_state_out_14_2_2[2:0]       ), //i
    .port_i_2_3 (keyAdd_port_state_out_14_2_3[2:0]       ), //i
    .port_i_2_4 (keyAdd_port_state_out_14_2_4[2:0]       ), //i
    .port_i_2_5 (keyAdd_port_state_out_14_2_5[2:0]       ), //i
    .port_i_2_6 (keyAdd_port_state_out_14_2_6[2:0]       ), //i
    .port_i_2_7 (keyAdd_port_state_out_14_2_7[2:0]       ), //i
    .port_i_3_0 (keyAdd_port_state_out_14_3_0[2:0]       ), //i
    .port_i_3_1 (keyAdd_port_state_out_14_3_1[2:0]       ), //i
    .port_i_3_2 (keyAdd_port_state_out_14_3_2[2:0]       ), //i
    .port_i_3_3 (keyAdd_port_state_out_14_3_3[2:0]       ), //i
    .port_i_3_4 (keyAdd_port_state_out_14_3_4[2:0]       ), //i
    .port_i_3_5 (keyAdd_port_state_out_14_3_5[2:0]       ), //i
    .port_i_3_6 (keyAdd_port_state_out_14_3_6[2:0]       ), //i
    .port_i_3_7 (keyAdd_port_state_out_14_3_7[2:0]       ), //i
    .port_o_0_0 (sbox_AES_BoyarPeralta_30_port_o_0_0[2:0]), //o
    .port_o_0_1 (sbox_AES_BoyarPeralta_30_port_o_0_1[2:0]), //o
    .port_o_0_2 (sbox_AES_BoyarPeralta_30_port_o_0_2[2:0]), //o
    .port_o_0_3 (sbox_AES_BoyarPeralta_30_port_o_0_3[2:0]), //o
    .port_o_0_4 (sbox_AES_BoyarPeralta_30_port_o_0_4[2:0]), //o
    .port_o_0_5 (sbox_AES_BoyarPeralta_30_port_o_0_5[2:0]), //o
    .port_o_0_6 (sbox_AES_BoyarPeralta_30_port_o_0_6[2:0]), //o
    .port_o_0_7 (sbox_AES_BoyarPeralta_30_port_o_0_7[2:0]), //o
    .port_o_1_0 (sbox_AES_BoyarPeralta_30_port_o_1_0[2:0]), //o
    .port_o_1_1 (sbox_AES_BoyarPeralta_30_port_o_1_1[2:0]), //o
    .port_o_1_2 (sbox_AES_BoyarPeralta_30_port_o_1_2[2:0]), //o
    .port_o_1_3 (sbox_AES_BoyarPeralta_30_port_o_1_3[2:0]), //o
    .port_o_1_4 (sbox_AES_BoyarPeralta_30_port_o_1_4[2:0]), //o
    .port_o_1_5 (sbox_AES_BoyarPeralta_30_port_o_1_5[2:0]), //o
    .port_o_1_6 (sbox_AES_BoyarPeralta_30_port_o_1_6[2:0]), //o
    .port_o_1_7 (sbox_AES_BoyarPeralta_30_port_o_1_7[2:0]), //o
    .port_o_2_0 (sbox_AES_BoyarPeralta_30_port_o_2_0[2:0]), //o
    .port_o_2_1 (sbox_AES_BoyarPeralta_30_port_o_2_1[2:0]), //o
    .port_o_2_2 (sbox_AES_BoyarPeralta_30_port_o_2_2[2:0]), //o
    .port_o_2_3 (sbox_AES_BoyarPeralta_30_port_o_2_3[2:0]), //o
    .port_o_2_4 (sbox_AES_BoyarPeralta_30_port_o_2_4[2:0]), //o
    .port_o_2_5 (sbox_AES_BoyarPeralta_30_port_o_2_5[2:0]), //o
    .port_o_2_6 (sbox_AES_BoyarPeralta_30_port_o_2_6[2:0]), //o
    .port_o_2_7 (sbox_AES_BoyarPeralta_30_port_o_2_7[2:0]), //o
    .port_o_3_0 (sbox_AES_BoyarPeralta_30_port_o_3_0[2:0]), //o
    .port_o_3_1 (sbox_AES_BoyarPeralta_30_port_o_3_1[2:0]), //o
    .port_o_3_2 (sbox_AES_BoyarPeralta_30_port_o_3_2[2:0]), //o
    .port_o_3_3 (sbox_AES_BoyarPeralta_30_port_o_3_3[2:0]), //o
    .port_o_3_4 (sbox_AES_BoyarPeralta_30_port_o_3_4[2:0]), //o
    .port_o_3_5 (sbox_AES_BoyarPeralta_30_port_o_3_5[2:0]), //o
    .port_o_3_6 (sbox_AES_BoyarPeralta_30_port_o_3_6[2:0]), //o
    .port_o_3_7 (sbox_AES_BoyarPeralta_30_port_o_3_7[2:0]), //o
    .clk        (clk                                     ), //i
    .reset      (reset                                   )  //i
  );
  Sbox_AES_BoyarPeralta sbox_AES_BoyarPeralta_31 (
    .port_i_0_0 (keyAdd_port_state_out_15_0_0[2:0]       ), //i
    .port_i_0_1 (keyAdd_port_state_out_15_0_1[2:0]       ), //i
    .port_i_0_2 (keyAdd_port_state_out_15_0_2[2:0]       ), //i
    .port_i_0_3 (keyAdd_port_state_out_15_0_3[2:0]       ), //i
    .port_i_0_4 (keyAdd_port_state_out_15_0_4[2:0]       ), //i
    .port_i_0_5 (keyAdd_port_state_out_15_0_5[2:0]       ), //i
    .port_i_0_6 (keyAdd_port_state_out_15_0_6[2:0]       ), //i
    .port_i_0_7 (keyAdd_port_state_out_15_0_7[2:0]       ), //i
    .port_i_1_0 (keyAdd_port_state_out_15_1_0[2:0]       ), //i
    .port_i_1_1 (keyAdd_port_state_out_15_1_1[2:0]       ), //i
    .port_i_1_2 (keyAdd_port_state_out_15_1_2[2:0]       ), //i
    .port_i_1_3 (keyAdd_port_state_out_15_1_3[2:0]       ), //i
    .port_i_1_4 (keyAdd_port_state_out_15_1_4[2:0]       ), //i
    .port_i_1_5 (keyAdd_port_state_out_15_1_5[2:0]       ), //i
    .port_i_1_6 (keyAdd_port_state_out_15_1_6[2:0]       ), //i
    .port_i_1_7 (keyAdd_port_state_out_15_1_7[2:0]       ), //i
    .port_i_2_0 (keyAdd_port_state_out_15_2_0[2:0]       ), //i
    .port_i_2_1 (keyAdd_port_state_out_15_2_1[2:0]       ), //i
    .port_i_2_2 (keyAdd_port_state_out_15_2_2[2:0]       ), //i
    .port_i_2_3 (keyAdd_port_state_out_15_2_3[2:0]       ), //i
    .port_i_2_4 (keyAdd_port_state_out_15_2_4[2:0]       ), //i
    .port_i_2_5 (keyAdd_port_state_out_15_2_5[2:0]       ), //i
    .port_i_2_6 (keyAdd_port_state_out_15_2_6[2:0]       ), //i
    .port_i_2_7 (keyAdd_port_state_out_15_2_7[2:0]       ), //i
    .port_i_3_0 (keyAdd_port_state_out_15_3_0[2:0]       ), //i
    .port_i_3_1 (keyAdd_port_state_out_15_3_1[2:0]       ), //i
    .port_i_3_2 (keyAdd_port_state_out_15_3_2[2:0]       ), //i
    .port_i_3_3 (keyAdd_port_state_out_15_3_3[2:0]       ), //i
    .port_i_3_4 (keyAdd_port_state_out_15_3_4[2:0]       ), //i
    .port_i_3_5 (keyAdd_port_state_out_15_3_5[2:0]       ), //i
    .port_i_3_6 (keyAdd_port_state_out_15_3_6[2:0]       ), //i
    .port_i_3_7 (keyAdd_port_state_out_15_3_7[2:0]       ), //i
    .port_o_0_0 (sbox_AES_BoyarPeralta_31_port_o_0_0[2:0]), //o
    .port_o_0_1 (sbox_AES_BoyarPeralta_31_port_o_0_1[2:0]), //o
    .port_o_0_2 (sbox_AES_BoyarPeralta_31_port_o_0_2[2:0]), //o
    .port_o_0_3 (sbox_AES_BoyarPeralta_31_port_o_0_3[2:0]), //o
    .port_o_0_4 (sbox_AES_BoyarPeralta_31_port_o_0_4[2:0]), //o
    .port_o_0_5 (sbox_AES_BoyarPeralta_31_port_o_0_5[2:0]), //o
    .port_o_0_6 (sbox_AES_BoyarPeralta_31_port_o_0_6[2:0]), //o
    .port_o_0_7 (sbox_AES_BoyarPeralta_31_port_o_0_7[2:0]), //o
    .port_o_1_0 (sbox_AES_BoyarPeralta_31_port_o_1_0[2:0]), //o
    .port_o_1_1 (sbox_AES_BoyarPeralta_31_port_o_1_1[2:0]), //o
    .port_o_1_2 (sbox_AES_BoyarPeralta_31_port_o_1_2[2:0]), //o
    .port_o_1_3 (sbox_AES_BoyarPeralta_31_port_o_1_3[2:0]), //o
    .port_o_1_4 (sbox_AES_BoyarPeralta_31_port_o_1_4[2:0]), //o
    .port_o_1_5 (sbox_AES_BoyarPeralta_31_port_o_1_5[2:0]), //o
    .port_o_1_6 (sbox_AES_BoyarPeralta_31_port_o_1_6[2:0]), //o
    .port_o_1_7 (sbox_AES_BoyarPeralta_31_port_o_1_7[2:0]), //o
    .port_o_2_0 (sbox_AES_BoyarPeralta_31_port_o_2_0[2:0]), //o
    .port_o_2_1 (sbox_AES_BoyarPeralta_31_port_o_2_1[2:0]), //o
    .port_o_2_2 (sbox_AES_BoyarPeralta_31_port_o_2_2[2:0]), //o
    .port_o_2_3 (sbox_AES_BoyarPeralta_31_port_o_2_3[2:0]), //o
    .port_o_2_4 (sbox_AES_BoyarPeralta_31_port_o_2_4[2:0]), //o
    .port_o_2_5 (sbox_AES_BoyarPeralta_31_port_o_2_5[2:0]), //o
    .port_o_2_6 (sbox_AES_BoyarPeralta_31_port_o_2_6[2:0]), //o
    .port_o_2_7 (sbox_AES_BoyarPeralta_31_port_o_2_7[2:0]), //o
    .port_o_3_0 (sbox_AES_BoyarPeralta_31_port_o_3_0[2:0]), //o
    .port_o_3_1 (sbox_AES_BoyarPeralta_31_port_o_3_1[2:0]), //o
    .port_o_3_2 (sbox_AES_BoyarPeralta_31_port_o_3_2[2:0]), //o
    .port_o_3_3 (sbox_AES_BoyarPeralta_31_port_o_3_3[2:0]), //o
    .port_o_3_4 (sbox_AES_BoyarPeralta_31_port_o_3_4[2:0]), //o
    .port_o_3_5 (sbox_AES_BoyarPeralta_31_port_o_3_5[2:0]), //o
    .port_o_3_6 (sbox_AES_BoyarPeralta_31_port_o_3_6[2:0]), //o
    .port_o_3_7 (sbox_AES_BoyarPeralta_31_port_o_3_7[2:0]), //o
    .clk        (clk                                     ), //i
    .reset      (reset                                   )  //i
  );
  AES_ShiftRows shiftRows (
    .port_state_in_0_0_0   (subBytes_out_0_0_0[2:0]             ), //i
    .port_state_in_0_0_1   (subBytes_out_0_0_1[2:0]             ), //i
    .port_state_in_0_0_2   (subBytes_out_0_0_2[2:0]             ), //i
    .port_state_in_0_0_3   (subBytes_out_0_0_3[2:0]             ), //i
    .port_state_in_0_0_4   (subBytes_out_0_0_4[2:0]             ), //i
    .port_state_in_0_0_5   (subBytes_out_0_0_5[2:0]             ), //i
    .port_state_in_0_0_6   (subBytes_out_0_0_6[2:0]             ), //i
    .port_state_in_0_0_7   (subBytes_out_0_0_7[2:0]             ), //i
    .port_state_in_0_1_0   (subBytes_out_0_1_0[2:0]             ), //i
    .port_state_in_0_1_1   (subBytes_out_0_1_1[2:0]             ), //i
    .port_state_in_0_1_2   (subBytes_out_0_1_2[2:0]             ), //i
    .port_state_in_0_1_3   (subBytes_out_0_1_3[2:0]             ), //i
    .port_state_in_0_1_4   (subBytes_out_0_1_4[2:0]             ), //i
    .port_state_in_0_1_5   (subBytes_out_0_1_5[2:0]             ), //i
    .port_state_in_0_1_6   (subBytes_out_0_1_6[2:0]             ), //i
    .port_state_in_0_1_7   (subBytes_out_0_1_7[2:0]             ), //i
    .port_state_in_0_2_0   (subBytes_out_0_2_0[2:0]             ), //i
    .port_state_in_0_2_1   (subBytes_out_0_2_1[2:0]             ), //i
    .port_state_in_0_2_2   (subBytes_out_0_2_2[2:0]             ), //i
    .port_state_in_0_2_3   (subBytes_out_0_2_3[2:0]             ), //i
    .port_state_in_0_2_4   (subBytes_out_0_2_4[2:0]             ), //i
    .port_state_in_0_2_5   (subBytes_out_0_2_5[2:0]             ), //i
    .port_state_in_0_2_6   (subBytes_out_0_2_6[2:0]             ), //i
    .port_state_in_0_2_7   (subBytes_out_0_2_7[2:0]             ), //i
    .port_state_in_0_3_0   (subBytes_out_0_3_0[2:0]             ), //i
    .port_state_in_0_3_1   (subBytes_out_0_3_1[2:0]             ), //i
    .port_state_in_0_3_2   (subBytes_out_0_3_2[2:0]             ), //i
    .port_state_in_0_3_3   (subBytes_out_0_3_3[2:0]             ), //i
    .port_state_in_0_3_4   (subBytes_out_0_3_4[2:0]             ), //i
    .port_state_in_0_3_5   (subBytes_out_0_3_5[2:0]             ), //i
    .port_state_in_0_3_6   (subBytes_out_0_3_6[2:0]             ), //i
    .port_state_in_0_3_7   (subBytes_out_0_3_7[2:0]             ), //i
    .port_state_in_1_0_0   (subBytes_out_1_0_0[2:0]             ), //i
    .port_state_in_1_0_1   (subBytes_out_1_0_1[2:0]             ), //i
    .port_state_in_1_0_2   (subBytes_out_1_0_2[2:0]             ), //i
    .port_state_in_1_0_3   (subBytes_out_1_0_3[2:0]             ), //i
    .port_state_in_1_0_4   (subBytes_out_1_0_4[2:0]             ), //i
    .port_state_in_1_0_5   (subBytes_out_1_0_5[2:0]             ), //i
    .port_state_in_1_0_6   (subBytes_out_1_0_6[2:0]             ), //i
    .port_state_in_1_0_7   (subBytes_out_1_0_7[2:0]             ), //i
    .port_state_in_1_1_0   (subBytes_out_1_1_0[2:0]             ), //i
    .port_state_in_1_1_1   (subBytes_out_1_1_1[2:0]             ), //i
    .port_state_in_1_1_2   (subBytes_out_1_1_2[2:0]             ), //i
    .port_state_in_1_1_3   (subBytes_out_1_1_3[2:0]             ), //i
    .port_state_in_1_1_4   (subBytes_out_1_1_4[2:0]             ), //i
    .port_state_in_1_1_5   (subBytes_out_1_1_5[2:0]             ), //i
    .port_state_in_1_1_6   (subBytes_out_1_1_6[2:0]             ), //i
    .port_state_in_1_1_7   (subBytes_out_1_1_7[2:0]             ), //i
    .port_state_in_1_2_0   (subBytes_out_1_2_0[2:0]             ), //i
    .port_state_in_1_2_1   (subBytes_out_1_2_1[2:0]             ), //i
    .port_state_in_1_2_2   (subBytes_out_1_2_2[2:0]             ), //i
    .port_state_in_1_2_3   (subBytes_out_1_2_3[2:0]             ), //i
    .port_state_in_1_2_4   (subBytes_out_1_2_4[2:0]             ), //i
    .port_state_in_1_2_5   (subBytes_out_1_2_5[2:0]             ), //i
    .port_state_in_1_2_6   (subBytes_out_1_2_6[2:0]             ), //i
    .port_state_in_1_2_7   (subBytes_out_1_2_7[2:0]             ), //i
    .port_state_in_1_3_0   (subBytes_out_1_3_0[2:0]             ), //i
    .port_state_in_1_3_1   (subBytes_out_1_3_1[2:0]             ), //i
    .port_state_in_1_3_2   (subBytes_out_1_3_2[2:0]             ), //i
    .port_state_in_1_3_3   (subBytes_out_1_3_3[2:0]             ), //i
    .port_state_in_1_3_4   (subBytes_out_1_3_4[2:0]             ), //i
    .port_state_in_1_3_5   (subBytes_out_1_3_5[2:0]             ), //i
    .port_state_in_1_3_6   (subBytes_out_1_3_6[2:0]             ), //i
    .port_state_in_1_3_7   (subBytes_out_1_3_7[2:0]             ), //i
    .port_state_in_2_0_0   (subBytes_out_2_0_0[2:0]             ), //i
    .port_state_in_2_0_1   (subBytes_out_2_0_1[2:0]             ), //i
    .port_state_in_2_0_2   (subBytes_out_2_0_2[2:0]             ), //i
    .port_state_in_2_0_3   (subBytes_out_2_0_3[2:0]             ), //i
    .port_state_in_2_0_4   (subBytes_out_2_0_4[2:0]             ), //i
    .port_state_in_2_0_5   (subBytes_out_2_0_5[2:0]             ), //i
    .port_state_in_2_0_6   (subBytes_out_2_0_6[2:0]             ), //i
    .port_state_in_2_0_7   (subBytes_out_2_0_7[2:0]             ), //i
    .port_state_in_2_1_0   (subBytes_out_2_1_0[2:0]             ), //i
    .port_state_in_2_1_1   (subBytes_out_2_1_1[2:0]             ), //i
    .port_state_in_2_1_2   (subBytes_out_2_1_2[2:0]             ), //i
    .port_state_in_2_1_3   (subBytes_out_2_1_3[2:0]             ), //i
    .port_state_in_2_1_4   (subBytes_out_2_1_4[2:0]             ), //i
    .port_state_in_2_1_5   (subBytes_out_2_1_5[2:0]             ), //i
    .port_state_in_2_1_6   (subBytes_out_2_1_6[2:0]             ), //i
    .port_state_in_2_1_7   (subBytes_out_2_1_7[2:0]             ), //i
    .port_state_in_2_2_0   (subBytes_out_2_2_0[2:0]             ), //i
    .port_state_in_2_2_1   (subBytes_out_2_2_1[2:0]             ), //i
    .port_state_in_2_2_2   (subBytes_out_2_2_2[2:0]             ), //i
    .port_state_in_2_2_3   (subBytes_out_2_2_3[2:0]             ), //i
    .port_state_in_2_2_4   (subBytes_out_2_2_4[2:0]             ), //i
    .port_state_in_2_2_5   (subBytes_out_2_2_5[2:0]             ), //i
    .port_state_in_2_2_6   (subBytes_out_2_2_6[2:0]             ), //i
    .port_state_in_2_2_7   (subBytes_out_2_2_7[2:0]             ), //i
    .port_state_in_2_3_0   (subBytes_out_2_3_0[2:0]             ), //i
    .port_state_in_2_3_1   (subBytes_out_2_3_1[2:0]             ), //i
    .port_state_in_2_3_2   (subBytes_out_2_3_2[2:0]             ), //i
    .port_state_in_2_3_3   (subBytes_out_2_3_3[2:0]             ), //i
    .port_state_in_2_3_4   (subBytes_out_2_3_4[2:0]             ), //i
    .port_state_in_2_3_5   (subBytes_out_2_3_5[2:0]             ), //i
    .port_state_in_2_3_6   (subBytes_out_2_3_6[2:0]             ), //i
    .port_state_in_2_3_7   (subBytes_out_2_3_7[2:0]             ), //i
    .port_state_in_3_0_0   (subBytes_out_3_0_0[2:0]             ), //i
    .port_state_in_3_0_1   (subBytes_out_3_0_1[2:0]             ), //i
    .port_state_in_3_0_2   (subBytes_out_3_0_2[2:0]             ), //i
    .port_state_in_3_0_3   (subBytes_out_3_0_3[2:0]             ), //i
    .port_state_in_3_0_4   (subBytes_out_3_0_4[2:0]             ), //i
    .port_state_in_3_0_5   (subBytes_out_3_0_5[2:0]             ), //i
    .port_state_in_3_0_6   (subBytes_out_3_0_6[2:0]             ), //i
    .port_state_in_3_0_7   (subBytes_out_3_0_7[2:0]             ), //i
    .port_state_in_3_1_0   (subBytes_out_3_1_0[2:0]             ), //i
    .port_state_in_3_1_1   (subBytes_out_3_1_1[2:0]             ), //i
    .port_state_in_3_1_2   (subBytes_out_3_1_2[2:0]             ), //i
    .port_state_in_3_1_3   (subBytes_out_3_1_3[2:0]             ), //i
    .port_state_in_3_1_4   (subBytes_out_3_1_4[2:0]             ), //i
    .port_state_in_3_1_5   (subBytes_out_3_1_5[2:0]             ), //i
    .port_state_in_3_1_6   (subBytes_out_3_1_6[2:0]             ), //i
    .port_state_in_3_1_7   (subBytes_out_3_1_7[2:0]             ), //i
    .port_state_in_3_2_0   (subBytes_out_3_2_0[2:0]             ), //i
    .port_state_in_3_2_1   (subBytes_out_3_2_1[2:0]             ), //i
    .port_state_in_3_2_2   (subBytes_out_3_2_2[2:0]             ), //i
    .port_state_in_3_2_3   (subBytes_out_3_2_3[2:0]             ), //i
    .port_state_in_3_2_4   (subBytes_out_3_2_4[2:0]             ), //i
    .port_state_in_3_2_5   (subBytes_out_3_2_5[2:0]             ), //i
    .port_state_in_3_2_6   (subBytes_out_3_2_6[2:0]             ), //i
    .port_state_in_3_2_7   (subBytes_out_3_2_7[2:0]             ), //i
    .port_state_in_3_3_0   (subBytes_out_3_3_0[2:0]             ), //i
    .port_state_in_3_3_1   (subBytes_out_3_3_1[2:0]             ), //i
    .port_state_in_3_3_2   (subBytes_out_3_3_2[2:0]             ), //i
    .port_state_in_3_3_3   (subBytes_out_3_3_3[2:0]             ), //i
    .port_state_in_3_3_4   (subBytes_out_3_3_4[2:0]             ), //i
    .port_state_in_3_3_5   (subBytes_out_3_3_5[2:0]             ), //i
    .port_state_in_3_3_6   (subBytes_out_3_3_6[2:0]             ), //i
    .port_state_in_3_3_7   (subBytes_out_3_3_7[2:0]             ), //i
    .port_state_in_4_0_0   (subBytes_out_4_0_0[2:0]             ), //i
    .port_state_in_4_0_1   (subBytes_out_4_0_1[2:0]             ), //i
    .port_state_in_4_0_2   (subBytes_out_4_0_2[2:0]             ), //i
    .port_state_in_4_0_3   (subBytes_out_4_0_3[2:0]             ), //i
    .port_state_in_4_0_4   (subBytes_out_4_0_4[2:0]             ), //i
    .port_state_in_4_0_5   (subBytes_out_4_0_5[2:0]             ), //i
    .port_state_in_4_0_6   (subBytes_out_4_0_6[2:0]             ), //i
    .port_state_in_4_0_7   (subBytes_out_4_0_7[2:0]             ), //i
    .port_state_in_4_1_0   (subBytes_out_4_1_0[2:0]             ), //i
    .port_state_in_4_1_1   (subBytes_out_4_1_1[2:0]             ), //i
    .port_state_in_4_1_2   (subBytes_out_4_1_2[2:0]             ), //i
    .port_state_in_4_1_3   (subBytes_out_4_1_3[2:0]             ), //i
    .port_state_in_4_1_4   (subBytes_out_4_1_4[2:0]             ), //i
    .port_state_in_4_1_5   (subBytes_out_4_1_5[2:0]             ), //i
    .port_state_in_4_1_6   (subBytes_out_4_1_6[2:0]             ), //i
    .port_state_in_4_1_7   (subBytes_out_4_1_7[2:0]             ), //i
    .port_state_in_4_2_0   (subBytes_out_4_2_0[2:0]             ), //i
    .port_state_in_4_2_1   (subBytes_out_4_2_1[2:0]             ), //i
    .port_state_in_4_2_2   (subBytes_out_4_2_2[2:0]             ), //i
    .port_state_in_4_2_3   (subBytes_out_4_2_3[2:0]             ), //i
    .port_state_in_4_2_4   (subBytes_out_4_2_4[2:0]             ), //i
    .port_state_in_4_2_5   (subBytes_out_4_2_5[2:0]             ), //i
    .port_state_in_4_2_6   (subBytes_out_4_2_6[2:0]             ), //i
    .port_state_in_4_2_7   (subBytes_out_4_2_7[2:0]             ), //i
    .port_state_in_4_3_0   (subBytes_out_4_3_0[2:0]             ), //i
    .port_state_in_4_3_1   (subBytes_out_4_3_1[2:0]             ), //i
    .port_state_in_4_3_2   (subBytes_out_4_3_2[2:0]             ), //i
    .port_state_in_4_3_3   (subBytes_out_4_3_3[2:0]             ), //i
    .port_state_in_4_3_4   (subBytes_out_4_3_4[2:0]             ), //i
    .port_state_in_4_3_5   (subBytes_out_4_3_5[2:0]             ), //i
    .port_state_in_4_3_6   (subBytes_out_4_3_6[2:0]             ), //i
    .port_state_in_4_3_7   (subBytes_out_4_3_7[2:0]             ), //i
    .port_state_in_5_0_0   (subBytes_out_5_0_0[2:0]             ), //i
    .port_state_in_5_0_1   (subBytes_out_5_0_1[2:0]             ), //i
    .port_state_in_5_0_2   (subBytes_out_5_0_2[2:0]             ), //i
    .port_state_in_5_0_3   (subBytes_out_5_0_3[2:0]             ), //i
    .port_state_in_5_0_4   (subBytes_out_5_0_4[2:0]             ), //i
    .port_state_in_5_0_5   (subBytes_out_5_0_5[2:0]             ), //i
    .port_state_in_5_0_6   (subBytes_out_5_0_6[2:0]             ), //i
    .port_state_in_5_0_7   (subBytes_out_5_0_7[2:0]             ), //i
    .port_state_in_5_1_0   (subBytes_out_5_1_0[2:0]             ), //i
    .port_state_in_5_1_1   (subBytes_out_5_1_1[2:0]             ), //i
    .port_state_in_5_1_2   (subBytes_out_5_1_2[2:0]             ), //i
    .port_state_in_5_1_3   (subBytes_out_5_1_3[2:0]             ), //i
    .port_state_in_5_1_4   (subBytes_out_5_1_4[2:0]             ), //i
    .port_state_in_5_1_5   (subBytes_out_5_1_5[2:0]             ), //i
    .port_state_in_5_1_6   (subBytes_out_5_1_6[2:0]             ), //i
    .port_state_in_5_1_7   (subBytes_out_5_1_7[2:0]             ), //i
    .port_state_in_5_2_0   (subBytes_out_5_2_0[2:0]             ), //i
    .port_state_in_5_2_1   (subBytes_out_5_2_1[2:0]             ), //i
    .port_state_in_5_2_2   (subBytes_out_5_2_2[2:0]             ), //i
    .port_state_in_5_2_3   (subBytes_out_5_2_3[2:0]             ), //i
    .port_state_in_5_2_4   (subBytes_out_5_2_4[2:0]             ), //i
    .port_state_in_5_2_5   (subBytes_out_5_2_5[2:0]             ), //i
    .port_state_in_5_2_6   (subBytes_out_5_2_6[2:0]             ), //i
    .port_state_in_5_2_7   (subBytes_out_5_2_7[2:0]             ), //i
    .port_state_in_5_3_0   (subBytes_out_5_3_0[2:0]             ), //i
    .port_state_in_5_3_1   (subBytes_out_5_3_1[2:0]             ), //i
    .port_state_in_5_3_2   (subBytes_out_5_3_2[2:0]             ), //i
    .port_state_in_5_3_3   (subBytes_out_5_3_3[2:0]             ), //i
    .port_state_in_5_3_4   (subBytes_out_5_3_4[2:0]             ), //i
    .port_state_in_5_3_5   (subBytes_out_5_3_5[2:0]             ), //i
    .port_state_in_5_3_6   (subBytes_out_5_3_6[2:0]             ), //i
    .port_state_in_5_3_7   (subBytes_out_5_3_7[2:0]             ), //i
    .port_state_in_6_0_0   (subBytes_out_6_0_0[2:0]             ), //i
    .port_state_in_6_0_1   (subBytes_out_6_0_1[2:0]             ), //i
    .port_state_in_6_0_2   (subBytes_out_6_0_2[2:0]             ), //i
    .port_state_in_6_0_3   (subBytes_out_6_0_3[2:0]             ), //i
    .port_state_in_6_0_4   (subBytes_out_6_0_4[2:0]             ), //i
    .port_state_in_6_0_5   (subBytes_out_6_0_5[2:0]             ), //i
    .port_state_in_6_0_6   (subBytes_out_6_0_6[2:0]             ), //i
    .port_state_in_6_0_7   (subBytes_out_6_0_7[2:0]             ), //i
    .port_state_in_6_1_0   (subBytes_out_6_1_0[2:0]             ), //i
    .port_state_in_6_1_1   (subBytes_out_6_1_1[2:0]             ), //i
    .port_state_in_6_1_2   (subBytes_out_6_1_2[2:0]             ), //i
    .port_state_in_6_1_3   (subBytes_out_6_1_3[2:0]             ), //i
    .port_state_in_6_1_4   (subBytes_out_6_1_4[2:0]             ), //i
    .port_state_in_6_1_5   (subBytes_out_6_1_5[2:0]             ), //i
    .port_state_in_6_1_6   (subBytes_out_6_1_6[2:0]             ), //i
    .port_state_in_6_1_7   (subBytes_out_6_1_7[2:0]             ), //i
    .port_state_in_6_2_0   (subBytes_out_6_2_0[2:0]             ), //i
    .port_state_in_6_2_1   (subBytes_out_6_2_1[2:0]             ), //i
    .port_state_in_6_2_2   (subBytes_out_6_2_2[2:0]             ), //i
    .port_state_in_6_2_3   (subBytes_out_6_2_3[2:0]             ), //i
    .port_state_in_6_2_4   (subBytes_out_6_2_4[2:0]             ), //i
    .port_state_in_6_2_5   (subBytes_out_6_2_5[2:0]             ), //i
    .port_state_in_6_2_6   (subBytes_out_6_2_6[2:0]             ), //i
    .port_state_in_6_2_7   (subBytes_out_6_2_7[2:0]             ), //i
    .port_state_in_6_3_0   (subBytes_out_6_3_0[2:0]             ), //i
    .port_state_in_6_3_1   (subBytes_out_6_3_1[2:0]             ), //i
    .port_state_in_6_3_2   (subBytes_out_6_3_2[2:0]             ), //i
    .port_state_in_6_3_3   (subBytes_out_6_3_3[2:0]             ), //i
    .port_state_in_6_3_4   (subBytes_out_6_3_4[2:0]             ), //i
    .port_state_in_6_3_5   (subBytes_out_6_3_5[2:0]             ), //i
    .port_state_in_6_3_6   (subBytes_out_6_3_6[2:0]             ), //i
    .port_state_in_6_3_7   (subBytes_out_6_3_7[2:0]             ), //i
    .port_state_in_7_0_0   (subBytes_out_7_0_0[2:0]             ), //i
    .port_state_in_7_0_1   (subBytes_out_7_0_1[2:0]             ), //i
    .port_state_in_7_0_2   (subBytes_out_7_0_2[2:0]             ), //i
    .port_state_in_7_0_3   (subBytes_out_7_0_3[2:0]             ), //i
    .port_state_in_7_0_4   (subBytes_out_7_0_4[2:0]             ), //i
    .port_state_in_7_0_5   (subBytes_out_7_0_5[2:0]             ), //i
    .port_state_in_7_0_6   (subBytes_out_7_0_6[2:0]             ), //i
    .port_state_in_7_0_7   (subBytes_out_7_0_7[2:0]             ), //i
    .port_state_in_7_1_0   (subBytes_out_7_1_0[2:0]             ), //i
    .port_state_in_7_1_1   (subBytes_out_7_1_1[2:0]             ), //i
    .port_state_in_7_1_2   (subBytes_out_7_1_2[2:0]             ), //i
    .port_state_in_7_1_3   (subBytes_out_7_1_3[2:0]             ), //i
    .port_state_in_7_1_4   (subBytes_out_7_1_4[2:0]             ), //i
    .port_state_in_7_1_5   (subBytes_out_7_1_5[2:0]             ), //i
    .port_state_in_7_1_6   (subBytes_out_7_1_6[2:0]             ), //i
    .port_state_in_7_1_7   (subBytes_out_7_1_7[2:0]             ), //i
    .port_state_in_7_2_0   (subBytes_out_7_2_0[2:0]             ), //i
    .port_state_in_7_2_1   (subBytes_out_7_2_1[2:0]             ), //i
    .port_state_in_7_2_2   (subBytes_out_7_2_2[2:0]             ), //i
    .port_state_in_7_2_3   (subBytes_out_7_2_3[2:0]             ), //i
    .port_state_in_7_2_4   (subBytes_out_7_2_4[2:0]             ), //i
    .port_state_in_7_2_5   (subBytes_out_7_2_5[2:0]             ), //i
    .port_state_in_7_2_6   (subBytes_out_7_2_6[2:0]             ), //i
    .port_state_in_7_2_7   (subBytes_out_7_2_7[2:0]             ), //i
    .port_state_in_7_3_0   (subBytes_out_7_3_0[2:0]             ), //i
    .port_state_in_7_3_1   (subBytes_out_7_3_1[2:0]             ), //i
    .port_state_in_7_3_2   (subBytes_out_7_3_2[2:0]             ), //i
    .port_state_in_7_3_3   (subBytes_out_7_3_3[2:0]             ), //i
    .port_state_in_7_3_4   (subBytes_out_7_3_4[2:0]             ), //i
    .port_state_in_7_3_5   (subBytes_out_7_3_5[2:0]             ), //i
    .port_state_in_7_3_6   (subBytes_out_7_3_6[2:0]             ), //i
    .port_state_in_7_3_7   (subBytes_out_7_3_7[2:0]             ), //i
    .port_state_in_8_0_0   (subBytes_out_8_0_0[2:0]             ), //i
    .port_state_in_8_0_1   (subBytes_out_8_0_1[2:0]             ), //i
    .port_state_in_8_0_2   (subBytes_out_8_0_2[2:0]             ), //i
    .port_state_in_8_0_3   (subBytes_out_8_0_3[2:0]             ), //i
    .port_state_in_8_0_4   (subBytes_out_8_0_4[2:0]             ), //i
    .port_state_in_8_0_5   (subBytes_out_8_0_5[2:0]             ), //i
    .port_state_in_8_0_6   (subBytes_out_8_0_6[2:0]             ), //i
    .port_state_in_8_0_7   (subBytes_out_8_0_7[2:0]             ), //i
    .port_state_in_8_1_0   (subBytes_out_8_1_0[2:0]             ), //i
    .port_state_in_8_1_1   (subBytes_out_8_1_1[2:0]             ), //i
    .port_state_in_8_1_2   (subBytes_out_8_1_2[2:0]             ), //i
    .port_state_in_8_1_3   (subBytes_out_8_1_3[2:0]             ), //i
    .port_state_in_8_1_4   (subBytes_out_8_1_4[2:0]             ), //i
    .port_state_in_8_1_5   (subBytes_out_8_1_5[2:0]             ), //i
    .port_state_in_8_1_6   (subBytes_out_8_1_6[2:0]             ), //i
    .port_state_in_8_1_7   (subBytes_out_8_1_7[2:0]             ), //i
    .port_state_in_8_2_0   (subBytes_out_8_2_0[2:0]             ), //i
    .port_state_in_8_2_1   (subBytes_out_8_2_1[2:0]             ), //i
    .port_state_in_8_2_2   (subBytes_out_8_2_2[2:0]             ), //i
    .port_state_in_8_2_3   (subBytes_out_8_2_3[2:0]             ), //i
    .port_state_in_8_2_4   (subBytes_out_8_2_4[2:0]             ), //i
    .port_state_in_8_2_5   (subBytes_out_8_2_5[2:0]             ), //i
    .port_state_in_8_2_6   (subBytes_out_8_2_6[2:0]             ), //i
    .port_state_in_8_2_7   (subBytes_out_8_2_7[2:0]             ), //i
    .port_state_in_8_3_0   (subBytes_out_8_3_0[2:0]             ), //i
    .port_state_in_8_3_1   (subBytes_out_8_3_1[2:0]             ), //i
    .port_state_in_8_3_2   (subBytes_out_8_3_2[2:0]             ), //i
    .port_state_in_8_3_3   (subBytes_out_8_3_3[2:0]             ), //i
    .port_state_in_8_3_4   (subBytes_out_8_3_4[2:0]             ), //i
    .port_state_in_8_3_5   (subBytes_out_8_3_5[2:0]             ), //i
    .port_state_in_8_3_6   (subBytes_out_8_3_6[2:0]             ), //i
    .port_state_in_8_3_7   (subBytes_out_8_3_7[2:0]             ), //i
    .port_state_in_9_0_0   (subBytes_out_9_0_0[2:0]             ), //i
    .port_state_in_9_0_1   (subBytes_out_9_0_1[2:0]             ), //i
    .port_state_in_9_0_2   (subBytes_out_9_0_2[2:0]             ), //i
    .port_state_in_9_0_3   (subBytes_out_9_0_3[2:0]             ), //i
    .port_state_in_9_0_4   (subBytes_out_9_0_4[2:0]             ), //i
    .port_state_in_9_0_5   (subBytes_out_9_0_5[2:0]             ), //i
    .port_state_in_9_0_6   (subBytes_out_9_0_6[2:0]             ), //i
    .port_state_in_9_0_7   (subBytes_out_9_0_7[2:0]             ), //i
    .port_state_in_9_1_0   (subBytes_out_9_1_0[2:0]             ), //i
    .port_state_in_9_1_1   (subBytes_out_9_1_1[2:0]             ), //i
    .port_state_in_9_1_2   (subBytes_out_9_1_2[2:0]             ), //i
    .port_state_in_9_1_3   (subBytes_out_9_1_3[2:0]             ), //i
    .port_state_in_9_1_4   (subBytes_out_9_1_4[2:0]             ), //i
    .port_state_in_9_1_5   (subBytes_out_9_1_5[2:0]             ), //i
    .port_state_in_9_1_6   (subBytes_out_9_1_6[2:0]             ), //i
    .port_state_in_9_1_7   (subBytes_out_9_1_7[2:0]             ), //i
    .port_state_in_9_2_0   (subBytes_out_9_2_0[2:0]             ), //i
    .port_state_in_9_2_1   (subBytes_out_9_2_1[2:0]             ), //i
    .port_state_in_9_2_2   (subBytes_out_9_2_2[2:0]             ), //i
    .port_state_in_9_2_3   (subBytes_out_9_2_3[2:0]             ), //i
    .port_state_in_9_2_4   (subBytes_out_9_2_4[2:0]             ), //i
    .port_state_in_9_2_5   (subBytes_out_9_2_5[2:0]             ), //i
    .port_state_in_9_2_6   (subBytes_out_9_2_6[2:0]             ), //i
    .port_state_in_9_2_7   (subBytes_out_9_2_7[2:0]             ), //i
    .port_state_in_9_3_0   (subBytes_out_9_3_0[2:0]             ), //i
    .port_state_in_9_3_1   (subBytes_out_9_3_1[2:0]             ), //i
    .port_state_in_9_3_2   (subBytes_out_9_3_2[2:0]             ), //i
    .port_state_in_9_3_3   (subBytes_out_9_3_3[2:0]             ), //i
    .port_state_in_9_3_4   (subBytes_out_9_3_4[2:0]             ), //i
    .port_state_in_9_3_5   (subBytes_out_9_3_5[2:0]             ), //i
    .port_state_in_9_3_6   (subBytes_out_9_3_6[2:0]             ), //i
    .port_state_in_9_3_7   (subBytes_out_9_3_7[2:0]             ), //i
    .port_state_in_10_0_0  (subBytes_out_10_0_0[2:0]            ), //i
    .port_state_in_10_0_1  (subBytes_out_10_0_1[2:0]            ), //i
    .port_state_in_10_0_2  (subBytes_out_10_0_2[2:0]            ), //i
    .port_state_in_10_0_3  (subBytes_out_10_0_3[2:0]            ), //i
    .port_state_in_10_0_4  (subBytes_out_10_0_4[2:0]            ), //i
    .port_state_in_10_0_5  (subBytes_out_10_0_5[2:0]            ), //i
    .port_state_in_10_0_6  (subBytes_out_10_0_6[2:0]            ), //i
    .port_state_in_10_0_7  (subBytes_out_10_0_7[2:0]            ), //i
    .port_state_in_10_1_0  (subBytes_out_10_1_0[2:0]            ), //i
    .port_state_in_10_1_1  (subBytes_out_10_1_1[2:0]            ), //i
    .port_state_in_10_1_2  (subBytes_out_10_1_2[2:0]            ), //i
    .port_state_in_10_1_3  (subBytes_out_10_1_3[2:0]            ), //i
    .port_state_in_10_1_4  (subBytes_out_10_1_4[2:0]            ), //i
    .port_state_in_10_1_5  (subBytes_out_10_1_5[2:0]            ), //i
    .port_state_in_10_1_6  (subBytes_out_10_1_6[2:0]            ), //i
    .port_state_in_10_1_7  (subBytes_out_10_1_7[2:0]            ), //i
    .port_state_in_10_2_0  (subBytes_out_10_2_0[2:0]            ), //i
    .port_state_in_10_2_1  (subBytes_out_10_2_1[2:0]            ), //i
    .port_state_in_10_2_2  (subBytes_out_10_2_2[2:0]            ), //i
    .port_state_in_10_2_3  (subBytes_out_10_2_3[2:0]            ), //i
    .port_state_in_10_2_4  (subBytes_out_10_2_4[2:0]            ), //i
    .port_state_in_10_2_5  (subBytes_out_10_2_5[2:0]            ), //i
    .port_state_in_10_2_6  (subBytes_out_10_2_6[2:0]            ), //i
    .port_state_in_10_2_7  (subBytes_out_10_2_7[2:0]            ), //i
    .port_state_in_10_3_0  (subBytes_out_10_3_0[2:0]            ), //i
    .port_state_in_10_3_1  (subBytes_out_10_3_1[2:0]            ), //i
    .port_state_in_10_3_2  (subBytes_out_10_3_2[2:0]            ), //i
    .port_state_in_10_3_3  (subBytes_out_10_3_3[2:0]            ), //i
    .port_state_in_10_3_4  (subBytes_out_10_3_4[2:0]            ), //i
    .port_state_in_10_3_5  (subBytes_out_10_3_5[2:0]            ), //i
    .port_state_in_10_3_6  (subBytes_out_10_3_6[2:0]            ), //i
    .port_state_in_10_3_7  (subBytes_out_10_3_7[2:0]            ), //i
    .port_state_in_11_0_0  (subBytes_out_11_0_0[2:0]            ), //i
    .port_state_in_11_0_1  (subBytes_out_11_0_1[2:0]            ), //i
    .port_state_in_11_0_2  (subBytes_out_11_0_2[2:0]            ), //i
    .port_state_in_11_0_3  (subBytes_out_11_0_3[2:0]            ), //i
    .port_state_in_11_0_4  (subBytes_out_11_0_4[2:0]            ), //i
    .port_state_in_11_0_5  (subBytes_out_11_0_5[2:0]            ), //i
    .port_state_in_11_0_6  (subBytes_out_11_0_6[2:0]            ), //i
    .port_state_in_11_0_7  (subBytes_out_11_0_7[2:0]            ), //i
    .port_state_in_11_1_0  (subBytes_out_11_1_0[2:0]            ), //i
    .port_state_in_11_1_1  (subBytes_out_11_1_1[2:0]            ), //i
    .port_state_in_11_1_2  (subBytes_out_11_1_2[2:0]            ), //i
    .port_state_in_11_1_3  (subBytes_out_11_1_3[2:0]            ), //i
    .port_state_in_11_1_4  (subBytes_out_11_1_4[2:0]            ), //i
    .port_state_in_11_1_5  (subBytes_out_11_1_5[2:0]            ), //i
    .port_state_in_11_1_6  (subBytes_out_11_1_6[2:0]            ), //i
    .port_state_in_11_1_7  (subBytes_out_11_1_7[2:0]            ), //i
    .port_state_in_11_2_0  (subBytes_out_11_2_0[2:0]            ), //i
    .port_state_in_11_2_1  (subBytes_out_11_2_1[2:0]            ), //i
    .port_state_in_11_2_2  (subBytes_out_11_2_2[2:0]            ), //i
    .port_state_in_11_2_3  (subBytes_out_11_2_3[2:0]            ), //i
    .port_state_in_11_2_4  (subBytes_out_11_2_4[2:0]            ), //i
    .port_state_in_11_2_5  (subBytes_out_11_2_5[2:0]            ), //i
    .port_state_in_11_2_6  (subBytes_out_11_2_6[2:0]            ), //i
    .port_state_in_11_2_7  (subBytes_out_11_2_7[2:0]            ), //i
    .port_state_in_11_3_0  (subBytes_out_11_3_0[2:0]            ), //i
    .port_state_in_11_3_1  (subBytes_out_11_3_1[2:0]            ), //i
    .port_state_in_11_3_2  (subBytes_out_11_3_2[2:0]            ), //i
    .port_state_in_11_3_3  (subBytes_out_11_3_3[2:0]            ), //i
    .port_state_in_11_3_4  (subBytes_out_11_3_4[2:0]            ), //i
    .port_state_in_11_3_5  (subBytes_out_11_3_5[2:0]            ), //i
    .port_state_in_11_3_6  (subBytes_out_11_3_6[2:0]            ), //i
    .port_state_in_11_3_7  (subBytes_out_11_3_7[2:0]            ), //i
    .port_state_in_12_0_0  (subBytes_out_12_0_0[2:0]            ), //i
    .port_state_in_12_0_1  (subBytes_out_12_0_1[2:0]            ), //i
    .port_state_in_12_0_2  (subBytes_out_12_0_2[2:0]            ), //i
    .port_state_in_12_0_3  (subBytes_out_12_0_3[2:0]            ), //i
    .port_state_in_12_0_4  (subBytes_out_12_0_4[2:0]            ), //i
    .port_state_in_12_0_5  (subBytes_out_12_0_5[2:0]            ), //i
    .port_state_in_12_0_6  (subBytes_out_12_0_6[2:0]            ), //i
    .port_state_in_12_0_7  (subBytes_out_12_0_7[2:0]            ), //i
    .port_state_in_12_1_0  (subBytes_out_12_1_0[2:0]            ), //i
    .port_state_in_12_1_1  (subBytes_out_12_1_1[2:0]            ), //i
    .port_state_in_12_1_2  (subBytes_out_12_1_2[2:0]            ), //i
    .port_state_in_12_1_3  (subBytes_out_12_1_3[2:0]            ), //i
    .port_state_in_12_1_4  (subBytes_out_12_1_4[2:0]            ), //i
    .port_state_in_12_1_5  (subBytes_out_12_1_5[2:0]            ), //i
    .port_state_in_12_1_6  (subBytes_out_12_1_6[2:0]            ), //i
    .port_state_in_12_1_7  (subBytes_out_12_1_7[2:0]            ), //i
    .port_state_in_12_2_0  (subBytes_out_12_2_0[2:0]            ), //i
    .port_state_in_12_2_1  (subBytes_out_12_2_1[2:0]            ), //i
    .port_state_in_12_2_2  (subBytes_out_12_2_2[2:0]            ), //i
    .port_state_in_12_2_3  (subBytes_out_12_2_3[2:0]            ), //i
    .port_state_in_12_2_4  (subBytes_out_12_2_4[2:0]            ), //i
    .port_state_in_12_2_5  (subBytes_out_12_2_5[2:0]            ), //i
    .port_state_in_12_2_6  (subBytes_out_12_2_6[2:0]            ), //i
    .port_state_in_12_2_7  (subBytes_out_12_2_7[2:0]            ), //i
    .port_state_in_12_3_0  (subBytes_out_12_3_0[2:0]            ), //i
    .port_state_in_12_3_1  (subBytes_out_12_3_1[2:0]            ), //i
    .port_state_in_12_3_2  (subBytes_out_12_3_2[2:0]            ), //i
    .port_state_in_12_3_3  (subBytes_out_12_3_3[2:0]            ), //i
    .port_state_in_12_3_4  (subBytes_out_12_3_4[2:0]            ), //i
    .port_state_in_12_3_5  (subBytes_out_12_3_5[2:0]            ), //i
    .port_state_in_12_3_6  (subBytes_out_12_3_6[2:0]            ), //i
    .port_state_in_12_3_7  (subBytes_out_12_3_7[2:0]            ), //i
    .port_state_in_13_0_0  (subBytes_out_13_0_0[2:0]            ), //i
    .port_state_in_13_0_1  (subBytes_out_13_0_1[2:0]            ), //i
    .port_state_in_13_0_2  (subBytes_out_13_0_2[2:0]            ), //i
    .port_state_in_13_0_3  (subBytes_out_13_0_3[2:0]            ), //i
    .port_state_in_13_0_4  (subBytes_out_13_0_4[2:0]            ), //i
    .port_state_in_13_0_5  (subBytes_out_13_0_5[2:0]            ), //i
    .port_state_in_13_0_6  (subBytes_out_13_0_6[2:0]            ), //i
    .port_state_in_13_0_7  (subBytes_out_13_0_7[2:0]            ), //i
    .port_state_in_13_1_0  (subBytes_out_13_1_0[2:0]            ), //i
    .port_state_in_13_1_1  (subBytes_out_13_1_1[2:0]            ), //i
    .port_state_in_13_1_2  (subBytes_out_13_1_2[2:0]            ), //i
    .port_state_in_13_1_3  (subBytes_out_13_1_3[2:0]            ), //i
    .port_state_in_13_1_4  (subBytes_out_13_1_4[2:0]            ), //i
    .port_state_in_13_1_5  (subBytes_out_13_1_5[2:0]            ), //i
    .port_state_in_13_1_6  (subBytes_out_13_1_6[2:0]            ), //i
    .port_state_in_13_1_7  (subBytes_out_13_1_7[2:0]            ), //i
    .port_state_in_13_2_0  (subBytes_out_13_2_0[2:0]            ), //i
    .port_state_in_13_2_1  (subBytes_out_13_2_1[2:0]            ), //i
    .port_state_in_13_2_2  (subBytes_out_13_2_2[2:0]            ), //i
    .port_state_in_13_2_3  (subBytes_out_13_2_3[2:0]            ), //i
    .port_state_in_13_2_4  (subBytes_out_13_2_4[2:0]            ), //i
    .port_state_in_13_2_5  (subBytes_out_13_2_5[2:0]            ), //i
    .port_state_in_13_2_6  (subBytes_out_13_2_6[2:0]            ), //i
    .port_state_in_13_2_7  (subBytes_out_13_2_7[2:0]            ), //i
    .port_state_in_13_3_0  (subBytes_out_13_3_0[2:0]            ), //i
    .port_state_in_13_3_1  (subBytes_out_13_3_1[2:0]            ), //i
    .port_state_in_13_3_2  (subBytes_out_13_3_2[2:0]            ), //i
    .port_state_in_13_3_3  (subBytes_out_13_3_3[2:0]            ), //i
    .port_state_in_13_3_4  (subBytes_out_13_3_4[2:0]            ), //i
    .port_state_in_13_3_5  (subBytes_out_13_3_5[2:0]            ), //i
    .port_state_in_13_3_6  (subBytes_out_13_3_6[2:0]            ), //i
    .port_state_in_13_3_7  (subBytes_out_13_3_7[2:0]            ), //i
    .port_state_in_14_0_0  (subBytes_out_14_0_0[2:0]            ), //i
    .port_state_in_14_0_1  (subBytes_out_14_0_1[2:0]            ), //i
    .port_state_in_14_0_2  (subBytes_out_14_0_2[2:0]            ), //i
    .port_state_in_14_0_3  (subBytes_out_14_0_3[2:0]            ), //i
    .port_state_in_14_0_4  (subBytes_out_14_0_4[2:0]            ), //i
    .port_state_in_14_0_5  (subBytes_out_14_0_5[2:0]            ), //i
    .port_state_in_14_0_6  (subBytes_out_14_0_6[2:0]            ), //i
    .port_state_in_14_0_7  (subBytes_out_14_0_7[2:0]            ), //i
    .port_state_in_14_1_0  (subBytes_out_14_1_0[2:0]            ), //i
    .port_state_in_14_1_1  (subBytes_out_14_1_1[2:0]            ), //i
    .port_state_in_14_1_2  (subBytes_out_14_1_2[2:0]            ), //i
    .port_state_in_14_1_3  (subBytes_out_14_1_3[2:0]            ), //i
    .port_state_in_14_1_4  (subBytes_out_14_1_4[2:0]            ), //i
    .port_state_in_14_1_5  (subBytes_out_14_1_5[2:0]            ), //i
    .port_state_in_14_1_6  (subBytes_out_14_1_6[2:0]            ), //i
    .port_state_in_14_1_7  (subBytes_out_14_1_7[2:0]            ), //i
    .port_state_in_14_2_0  (subBytes_out_14_2_0[2:0]            ), //i
    .port_state_in_14_2_1  (subBytes_out_14_2_1[2:0]            ), //i
    .port_state_in_14_2_2  (subBytes_out_14_2_2[2:0]            ), //i
    .port_state_in_14_2_3  (subBytes_out_14_2_3[2:0]            ), //i
    .port_state_in_14_2_4  (subBytes_out_14_2_4[2:0]            ), //i
    .port_state_in_14_2_5  (subBytes_out_14_2_5[2:0]            ), //i
    .port_state_in_14_2_6  (subBytes_out_14_2_6[2:0]            ), //i
    .port_state_in_14_2_7  (subBytes_out_14_2_7[2:0]            ), //i
    .port_state_in_14_3_0  (subBytes_out_14_3_0[2:0]            ), //i
    .port_state_in_14_3_1  (subBytes_out_14_3_1[2:0]            ), //i
    .port_state_in_14_3_2  (subBytes_out_14_3_2[2:0]            ), //i
    .port_state_in_14_3_3  (subBytes_out_14_3_3[2:0]            ), //i
    .port_state_in_14_3_4  (subBytes_out_14_3_4[2:0]            ), //i
    .port_state_in_14_3_5  (subBytes_out_14_3_5[2:0]            ), //i
    .port_state_in_14_3_6  (subBytes_out_14_3_6[2:0]            ), //i
    .port_state_in_14_3_7  (subBytes_out_14_3_7[2:0]            ), //i
    .port_state_in_15_0_0  (subBytes_out_15_0_0[2:0]            ), //i
    .port_state_in_15_0_1  (subBytes_out_15_0_1[2:0]            ), //i
    .port_state_in_15_0_2  (subBytes_out_15_0_2[2:0]            ), //i
    .port_state_in_15_0_3  (subBytes_out_15_0_3[2:0]            ), //i
    .port_state_in_15_0_4  (subBytes_out_15_0_4[2:0]            ), //i
    .port_state_in_15_0_5  (subBytes_out_15_0_5[2:0]            ), //i
    .port_state_in_15_0_6  (subBytes_out_15_0_6[2:0]            ), //i
    .port_state_in_15_0_7  (subBytes_out_15_0_7[2:0]            ), //i
    .port_state_in_15_1_0  (subBytes_out_15_1_0[2:0]            ), //i
    .port_state_in_15_1_1  (subBytes_out_15_1_1[2:0]            ), //i
    .port_state_in_15_1_2  (subBytes_out_15_1_2[2:0]            ), //i
    .port_state_in_15_1_3  (subBytes_out_15_1_3[2:0]            ), //i
    .port_state_in_15_1_4  (subBytes_out_15_1_4[2:0]            ), //i
    .port_state_in_15_1_5  (subBytes_out_15_1_5[2:0]            ), //i
    .port_state_in_15_1_6  (subBytes_out_15_1_6[2:0]            ), //i
    .port_state_in_15_1_7  (subBytes_out_15_1_7[2:0]            ), //i
    .port_state_in_15_2_0  (subBytes_out_15_2_0[2:0]            ), //i
    .port_state_in_15_2_1  (subBytes_out_15_2_1[2:0]            ), //i
    .port_state_in_15_2_2  (subBytes_out_15_2_2[2:0]            ), //i
    .port_state_in_15_2_3  (subBytes_out_15_2_3[2:0]            ), //i
    .port_state_in_15_2_4  (subBytes_out_15_2_4[2:0]            ), //i
    .port_state_in_15_2_5  (subBytes_out_15_2_5[2:0]            ), //i
    .port_state_in_15_2_6  (subBytes_out_15_2_6[2:0]            ), //i
    .port_state_in_15_2_7  (subBytes_out_15_2_7[2:0]            ), //i
    .port_state_in_15_3_0  (subBytes_out_15_3_0[2:0]            ), //i
    .port_state_in_15_3_1  (subBytes_out_15_3_1[2:0]            ), //i
    .port_state_in_15_3_2  (subBytes_out_15_3_2[2:0]            ), //i
    .port_state_in_15_3_3  (subBytes_out_15_3_3[2:0]            ), //i
    .port_state_in_15_3_4  (subBytes_out_15_3_4[2:0]            ), //i
    .port_state_in_15_3_5  (subBytes_out_15_3_5[2:0]            ), //i
    .port_state_in_15_3_6  (subBytes_out_15_3_6[2:0]            ), //i
    .port_state_in_15_3_7  (subBytes_out_15_3_7[2:0]            ), //i
    .port_state_out_0_0_0  (shiftRows_port_state_out_0_0_0[2:0] ), //o
    .port_state_out_0_0_1  (shiftRows_port_state_out_0_0_1[2:0] ), //o
    .port_state_out_0_0_2  (shiftRows_port_state_out_0_0_2[2:0] ), //o
    .port_state_out_0_0_3  (shiftRows_port_state_out_0_0_3[2:0] ), //o
    .port_state_out_0_0_4  (shiftRows_port_state_out_0_0_4[2:0] ), //o
    .port_state_out_0_0_5  (shiftRows_port_state_out_0_0_5[2:0] ), //o
    .port_state_out_0_0_6  (shiftRows_port_state_out_0_0_6[2:0] ), //o
    .port_state_out_0_0_7  (shiftRows_port_state_out_0_0_7[2:0] ), //o
    .port_state_out_0_1_0  (shiftRows_port_state_out_0_1_0[2:0] ), //o
    .port_state_out_0_1_1  (shiftRows_port_state_out_0_1_1[2:0] ), //o
    .port_state_out_0_1_2  (shiftRows_port_state_out_0_1_2[2:0] ), //o
    .port_state_out_0_1_3  (shiftRows_port_state_out_0_1_3[2:0] ), //o
    .port_state_out_0_1_4  (shiftRows_port_state_out_0_1_4[2:0] ), //o
    .port_state_out_0_1_5  (shiftRows_port_state_out_0_1_5[2:0] ), //o
    .port_state_out_0_1_6  (shiftRows_port_state_out_0_1_6[2:0] ), //o
    .port_state_out_0_1_7  (shiftRows_port_state_out_0_1_7[2:0] ), //o
    .port_state_out_0_2_0  (shiftRows_port_state_out_0_2_0[2:0] ), //o
    .port_state_out_0_2_1  (shiftRows_port_state_out_0_2_1[2:0] ), //o
    .port_state_out_0_2_2  (shiftRows_port_state_out_0_2_2[2:0] ), //o
    .port_state_out_0_2_3  (shiftRows_port_state_out_0_2_3[2:0] ), //o
    .port_state_out_0_2_4  (shiftRows_port_state_out_0_2_4[2:0] ), //o
    .port_state_out_0_2_5  (shiftRows_port_state_out_0_2_5[2:0] ), //o
    .port_state_out_0_2_6  (shiftRows_port_state_out_0_2_6[2:0] ), //o
    .port_state_out_0_2_7  (shiftRows_port_state_out_0_2_7[2:0] ), //o
    .port_state_out_0_3_0  (shiftRows_port_state_out_0_3_0[2:0] ), //o
    .port_state_out_0_3_1  (shiftRows_port_state_out_0_3_1[2:0] ), //o
    .port_state_out_0_3_2  (shiftRows_port_state_out_0_3_2[2:0] ), //o
    .port_state_out_0_3_3  (shiftRows_port_state_out_0_3_3[2:0] ), //o
    .port_state_out_0_3_4  (shiftRows_port_state_out_0_3_4[2:0] ), //o
    .port_state_out_0_3_5  (shiftRows_port_state_out_0_3_5[2:0] ), //o
    .port_state_out_0_3_6  (shiftRows_port_state_out_0_3_6[2:0] ), //o
    .port_state_out_0_3_7  (shiftRows_port_state_out_0_3_7[2:0] ), //o
    .port_state_out_1_0_0  (shiftRows_port_state_out_1_0_0[2:0] ), //o
    .port_state_out_1_0_1  (shiftRows_port_state_out_1_0_1[2:0] ), //o
    .port_state_out_1_0_2  (shiftRows_port_state_out_1_0_2[2:0] ), //o
    .port_state_out_1_0_3  (shiftRows_port_state_out_1_0_3[2:0] ), //o
    .port_state_out_1_0_4  (shiftRows_port_state_out_1_0_4[2:0] ), //o
    .port_state_out_1_0_5  (shiftRows_port_state_out_1_0_5[2:0] ), //o
    .port_state_out_1_0_6  (shiftRows_port_state_out_1_0_6[2:0] ), //o
    .port_state_out_1_0_7  (shiftRows_port_state_out_1_0_7[2:0] ), //o
    .port_state_out_1_1_0  (shiftRows_port_state_out_1_1_0[2:0] ), //o
    .port_state_out_1_1_1  (shiftRows_port_state_out_1_1_1[2:0] ), //o
    .port_state_out_1_1_2  (shiftRows_port_state_out_1_1_2[2:0] ), //o
    .port_state_out_1_1_3  (shiftRows_port_state_out_1_1_3[2:0] ), //o
    .port_state_out_1_1_4  (shiftRows_port_state_out_1_1_4[2:0] ), //o
    .port_state_out_1_1_5  (shiftRows_port_state_out_1_1_5[2:0] ), //o
    .port_state_out_1_1_6  (shiftRows_port_state_out_1_1_6[2:0] ), //o
    .port_state_out_1_1_7  (shiftRows_port_state_out_1_1_7[2:0] ), //o
    .port_state_out_1_2_0  (shiftRows_port_state_out_1_2_0[2:0] ), //o
    .port_state_out_1_2_1  (shiftRows_port_state_out_1_2_1[2:0] ), //o
    .port_state_out_1_2_2  (shiftRows_port_state_out_1_2_2[2:0] ), //o
    .port_state_out_1_2_3  (shiftRows_port_state_out_1_2_3[2:0] ), //o
    .port_state_out_1_2_4  (shiftRows_port_state_out_1_2_4[2:0] ), //o
    .port_state_out_1_2_5  (shiftRows_port_state_out_1_2_5[2:0] ), //o
    .port_state_out_1_2_6  (shiftRows_port_state_out_1_2_6[2:0] ), //o
    .port_state_out_1_2_7  (shiftRows_port_state_out_1_2_7[2:0] ), //o
    .port_state_out_1_3_0  (shiftRows_port_state_out_1_3_0[2:0] ), //o
    .port_state_out_1_3_1  (shiftRows_port_state_out_1_3_1[2:0] ), //o
    .port_state_out_1_3_2  (shiftRows_port_state_out_1_3_2[2:0] ), //o
    .port_state_out_1_3_3  (shiftRows_port_state_out_1_3_3[2:0] ), //o
    .port_state_out_1_3_4  (shiftRows_port_state_out_1_3_4[2:0] ), //o
    .port_state_out_1_3_5  (shiftRows_port_state_out_1_3_5[2:0] ), //o
    .port_state_out_1_3_6  (shiftRows_port_state_out_1_3_6[2:0] ), //o
    .port_state_out_1_3_7  (shiftRows_port_state_out_1_3_7[2:0] ), //o
    .port_state_out_2_0_0  (shiftRows_port_state_out_2_0_0[2:0] ), //o
    .port_state_out_2_0_1  (shiftRows_port_state_out_2_0_1[2:0] ), //o
    .port_state_out_2_0_2  (shiftRows_port_state_out_2_0_2[2:0] ), //o
    .port_state_out_2_0_3  (shiftRows_port_state_out_2_0_3[2:0] ), //o
    .port_state_out_2_0_4  (shiftRows_port_state_out_2_0_4[2:0] ), //o
    .port_state_out_2_0_5  (shiftRows_port_state_out_2_0_5[2:0] ), //o
    .port_state_out_2_0_6  (shiftRows_port_state_out_2_0_6[2:0] ), //o
    .port_state_out_2_0_7  (shiftRows_port_state_out_2_0_7[2:0] ), //o
    .port_state_out_2_1_0  (shiftRows_port_state_out_2_1_0[2:0] ), //o
    .port_state_out_2_1_1  (shiftRows_port_state_out_2_1_1[2:0] ), //o
    .port_state_out_2_1_2  (shiftRows_port_state_out_2_1_2[2:0] ), //o
    .port_state_out_2_1_3  (shiftRows_port_state_out_2_1_3[2:0] ), //o
    .port_state_out_2_1_4  (shiftRows_port_state_out_2_1_4[2:0] ), //o
    .port_state_out_2_1_5  (shiftRows_port_state_out_2_1_5[2:0] ), //o
    .port_state_out_2_1_6  (shiftRows_port_state_out_2_1_6[2:0] ), //o
    .port_state_out_2_1_7  (shiftRows_port_state_out_2_1_7[2:0] ), //o
    .port_state_out_2_2_0  (shiftRows_port_state_out_2_2_0[2:0] ), //o
    .port_state_out_2_2_1  (shiftRows_port_state_out_2_2_1[2:0] ), //o
    .port_state_out_2_2_2  (shiftRows_port_state_out_2_2_2[2:0] ), //o
    .port_state_out_2_2_3  (shiftRows_port_state_out_2_2_3[2:0] ), //o
    .port_state_out_2_2_4  (shiftRows_port_state_out_2_2_4[2:0] ), //o
    .port_state_out_2_2_5  (shiftRows_port_state_out_2_2_5[2:0] ), //o
    .port_state_out_2_2_6  (shiftRows_port_state_out_2_2_6[2:0] ), //o
    .port_state_out_2_2_7  (shiftRows_port_state_out_2_2_7[2:0] ), //o
    .port_state_out_2_3_0  (shiftRows_port_state_out_2_3_0[2:0] ), //o
    .port_state_out_2_3_1  (shiftRows_port_state_out_2_3_1[2:0] ), //o
    .port_state_out_2_3_2  (shiftRows_port_state_out_2_3_2[2:0] ), //o
    .port_state_out_2_3_3  (shiftRows_port_state_out_2_3_3[2:0] ), //o
    .port_state_out_2_3_4  (shiftRows_port_state_out_2_3_4[2:0] ), //o
    .port_state_out_2_3_5  (shiftRows_port_state_out_2_3_5[2:0] ), //o
    .port_state_out_2_3_6  (shiftRows_port_state_out_2_3_6[2:0] ), //o
    .port_state_out_2_3_7  (shiftRows_port_state_out_2_3_7[2:0] ), //o
    .port_state_out_3_0_0  (shiftRows_port_state_out_3_0_0[2:0] ), //o
    .port_state_out_3_0_1  (shiftRows_port_state_out_3_0_1[2:0] ), //o
    .port_state_out_3_0_2  (shiftRows_port_state_out_3_0_2[2:0] ), //o
    .port_state_out_3_0_3  (shiftRows_port_state_out_3_0_3[2:0] ), //o
    .port_state_out_3_0_4  (shiftRows_port_state_out_3_0_4[2:0] ), //o
    .port_state_out_3_0_5  (shiftRows_port_state_out_3_0_5[2:0] ), //o
    .port_state_out_3_0_6  (shiftRows_port_state_out_3_0_6[2:0] ), //o
    .port_state_out_3_0_7  (shiftRows_port_state_out_3_0_7[2:0] ), //o
    .port_state_out_3_1_0  (shiftRows_port_state_out_3_1_0[2:0] ), //o
    .port_state_out_3_1_1  (shiftRows_port_state_out_3_1_1[2:0] ), //o
    .port_state_out_3_1_2  (shiftRows_port_state_out_3_1_2[2:0] ), //o
    .port_state_out_3_1_3  (shiftRows_port_state_out_3_1_3[2:0] ), //o
    .port_state_out_3_1_4  (shiftRows_port_state_out_3_1_4[2:0] ), //o
    .port_state_out_3_1_5  (shiftRows_port_state_out_3_1_5[2:0] ), //o
    .port_state_out_3_1_6  (shiftRows_port_state_out_3_1_6[2:0] ), //o
    .port_state_out_3_1_7  (shiftRows_port_state_out_3_1_7[2:0] ), //o
    .port_state_out_3_2_0  (shiftRows_port_state_out_3_2_0[2:0] ), //o
    .port_state_out_3_2_1  (shiftRows_port_state_out_3_2_1[2:0] ), //o
    .port_state_out_3_2_2  (shiftRows_port_state_out_3_2_2[2:0] ), //o
    .port_state_out_3_2_3  (shiftRows_port_state_out_3_2_3[2:0] ), //o
    .port_state_out_3_2_4  (shiftRows_port_state_out_3_2_4[2:0] ), //o
    .port_state_out_3_2_5  (shiftRows_port_state_out_3_2_5[2:0] ), //o
    .port_state_out_3_2_6  (shiftRows_port_state_out_3_2_6[2:0] ), //o
    .port_state_out_3_2_7  (shiftRows_port_state_out_3_2_7[2:0] ), //o
    .port_state_out_3_3_0  (shiftRows_port_state_out_3_3_0[2:0] ), //o
    .port_state_out_3_3_1  (shiftRows_port_state_out_3_3_1[2:0] ), //o
    .port_state_out_3_3_2  (shiftRows_port_state_out_3_3_2[2:0] ), //o
    .port_state_out_3_3_3  (shiftRows_port_state_out_3_3_3[2:0] ), //o
    .port_state_out_3_3_4  (shiftRows_port_state_out_3_3_4[2:0] ), //o
    .port_state_out_3_3_5  (shiftRows_port_state_out_3_3_5[2:0] ), //o
    .port_state_out_3_3_6  (shiftRows_port_state_out_3_3_6[2:0] ), //o
    .port_state_out_3_3_7  (shiftRows_port_state_out_3_3_7[2:0] ), //o
    .port_state_out_4_0_0  (shiftRows_port_state_out_4_0_0[2:0] ), //o
    .port_state_out_4_0_1  (shiftRows_port_state_out_4_0_1[2:0] ), //o
    .port_state_out_4_0_2  (shiftRows_port_state_out_4_0_2[2:0] ), //o
    .port_state_out_4_0_3  (shiftRows_port_state_out_4_0_3[2:0] ), //o
    .port_state_out_4_0_4  (shiftRows_port_state_out_4_0_4[2:0] ), //o
    .port_state_out_4_0_5  (shiftRows_port_state_out_4_0_5[2:0] ), //o
    .port_state_out_4_0_6  (shiftRows_port_state_out_4_0_6[2:0] ), //o
    .port_state_out_4_0_7  (shiftRows_port_state_out_4_0_7[2:0] ), //o
    .port_state_out_4_1_0  (shiftRows_port_state_out_4_1_0[2:0] ), //o
    .port_state_out_4_1_1  (shiftRows_port_state_out_4_1_1[2:0] ), //o
    .port_state_out_4_1_2  (shiftRows_port_state_out_4_1_2[2:0] ), //o
    .port_state_out_4_1_3  (shiftRows_port_state_out_4_1_3[2:0] ), //o
    .port_state_out_4_1_4  (shiftRows_port_state_out_4_1_4[2:0] ), //o
    .port_state_out_4_1_5  (shiftRows_port_state_out_4_1_5[2:0] ), //o
    .port_state_out_4_1_6  (shiftRows_port_state_out_4_1_6[2:0] ), //o
    .port_state_out_4_1_7  (shiftRows_port_state_out_4_1_7[2:0] ), //o
    .port_state_out_4_2_0  (shiftRows_port_state_out_4_2_0[2:0] ), //o
    .port_state_out_4_2_1  (shiftRows_port_state_out_4_2_1[2:0] ), //o
    .port_state_out_4_2_2  (shiftRows_port_state_out_4_2_2[2:0] ), //o
    .port_state_out_4_2_3  (shiftRows_port_state_out_4_2_3[2:0] ), //o
    .port_state_out_4_2_4  (shiftRows_port_state_out_4_2_4[2:0] ), //o
    .port_state_out_4_2_5  (shiftRows_port_state_out_4_2_5[2:0] ), //o
    .port_state_out_4_2_6  (shiftRows_port_state_out_4_2_6[2:0] ), //o
    .port_state_out_4_2_7  (shiftRows_port_state_out_4_2_7[2:0] ), //o
    .port_state_out_4_3_0  (shiftRows_port_state_out_4_3_0[2:0] ), //o
    .port_state_out_4_3_1  (shiftRows_port_state_out_4_3_1[2:0] ), //o
    .port_state_out_4_3_2  (shiftRows_port_state_out_4_3_2[2:0] ), //o
    .port_state_out_4_3_3  (shiftRows_port_state_out_4_3_3[2:0] ), //o
    .port_state_out_4_3_4  (shiftRows_port_state_out_4_3_4[2:0] ), //o
    .port_state_out_4_3_5  (shiftRows_port_state_out_4_3_5[2:0] ), //o
    .port_state_out_4_3_6  (shiftRows_port_state_out_4_3_6[2:0] ), //o
    .port_state_out_4_3_7  (shiftRows_port_state_out_4_3_7[2:0] ), //o
    .port_state_out_5_0_0  (shiftRows_port_state_out_5_0_0[2:0] ), //o
    .port_state_out_5_0_1  (shiftRows_port_state_out_5_0_1[2:0] ), //o
    .port_state_out_5_0_2  (shiftRows_port_state_out_5_0_2[2:0] ), //o
    .port_state_out_5_0_3  (shiftRows_port_state_out_5_0_3[2:0] ), //o
    .port_state_out_5_0_4  (shiftRows_port_state_out_5_0_4[2:0] ), //o
    .port_state_out_5_0_5  (shiftRows_port_state_out_5_0_5[2:0] ), //o
    .port_state_out_5_0_6  (shiftRows_port_state_out_5_0_6[2:0] ), //o
    .port_state_out_5_0_7  (shiftRows_port_state_out_5_0_7[2:0] ), //o
    .port_state_out_5_1_0  (shiftRows_port_state_out_5_1_0[2:0] ), //o
    .port_state_out_5_1_1  (shiftRows_port_state_out_5_1_1[2:0] ), //o
    .port_state_out_5_1_2  (shiftRows_port_state_out_5_1_2[2:0] ), //o
    .port_state_out_5_1_3  (shiftRows_port_state_out_5_1_3[2:0] ), //o
    .port_state_out_5_1_4  (shiftRows_port_state_out_5_1_4[2:0] ), //o
    .port_state_out_5_1_5  (shiftRows_port_state_out_5_1_5[2:0] ), //o
    .port_state_out_5_1_6  (shiftRows_port_state_out_5_1_6[2:0] ), //o
    .port_state_out_5_1_7  (shiftRows_port_state_out_5_1_7[2:0] ), //o
    .port_state_out_5_2_0  (shiftRows_port_state_out_5_2_0[2:0] ), //o
    .port_state_out_5_2_1  (shiftRows_port_state_out_5_2_1[2:0] ), //o
    .port_state_out_5_2_2  (shiftRows_port_state_out_5_2_2[2:0] ), //o
    .port_state_out_5_2_3  (shiftRows_port_state_out_5_2_3[2:0] ), //o
    .port_state_out_5_2_4  (shiftRows_port_state_out_5_2_4[2:0] ), //o
    .port_state_out_5_2_5  (shiftRows_port_state_out_5_2_5[2:0] ), //o
    .port_state_out_5_2_6  (shiftRows_port_state_out_5_2_6[2:0] ), //o
    .port_state_out_5_2_7  (shiftRows_port_state_out_5_2_7[2:0] ), //o
    .port_state_out_5_3_0  (shiftRows_port_state_out_5_3_0[2:0] ), //o
    .port_state_out_5_3_1  (shiftRows_port_state_out_5_3_1[2:0] ), //o
    .port_state_out_5_3_2  (shiftRows_port_state_out_5_3_2[2:0] ), //o
    .port_state_out_5_3_3  (shiftRows_port_state_out_5_3_3[2:0] ), //o
    .port_state_out_5_3_4  (shiftRows_port_state_out_5_3_4[2:0] ), //o
    .port_state_out_5_3_5  (shiftRows_port_state_out_5_3_5[2:0] ), //o
    .port_state_out_5_3_6  (shiftRows_port_state_out_5_3_6[2:0] ), //o
    .port_state_out_5_3_7  (shiftRows_port_state_out_5_3_7[2:0] ), //o
    .port_state_out_6_0_0  (shiftRows_port_state_out_6_0_0[2:0] ), //o
    .port_state_out_6_0_1  (shiftRows_port_state_out_6_0_1[2:0] ), //o
    .port_state_out_6_0_2  (shiftRows_port_state_out_6_0_2[2:0] ), //o
    .port_state_out_6_0_3  (shiftRows_port_state_out_6_0_3[2:0] ), //o
    .port_state_out_6_0_4  (shiftRows_port_state_out_6_0_4[2:0] ), //o
    .port_state_out_6_0_5  (shiftRows_port_state_out_6_0_5[2:0] ), //o
    .port_state_out_6_0_6  (shiftRows_port_state_out_6_0_6[2:0] ), //o
    .port_state_out_6_0_7  (shiftRows_port_state_out_6_0_7[2:0] ), //o
    .port_state_out_6_1_0  (shiftRows_port_state_out_6_1_0[2:0] ), //o
    .port_state_out_6_1_1  (shiftRows_port_state_out_6_1_1[2:0] ), //o
    .port_state_out_6_1_2  (shiftRows_port_state_out_6_1_2[2:0] ), //o
    .port_state_out_6_1_3  (shiftRows_port_state_out_6_1_3[2:0] ), //o
    .port_state_out_6_1_4  (shiftRows_port_state_out_6_1_4[2:0] ), //o
    .port_state_out_6_1_5  (shiftRows_port_state_out_6_1_5[2:0] ), //o
    .port_state_out_6_1_6  (shiftRows_port_state_out_6_1_6[2:0] ), //o
    .port_state_out_6_1_7  (shiftRows_port_state_out_6_1_7[2:0] ), //o
    .port_state_out_6_2_0  (shiftRows_port_state_out_6_2_0[2:0] ), //o
    .port_state_out_6_2_1  (shiftRows_port_state_out_6_2_1[2:0] ), //o
    .port_state_out_6_2_2  (shiftRows_port_state_out_6_2_2[2:0] ), //o
    .port_state_out_6_2_3  (shiftRows_port_state_out_6_2_3[2:0] ), //o
    .port_state_out_6_2_4  (shiftRows_port_state_out_6_2_4[2:0] ), //o
    .port_state_out_6_2_5  (shiftRows_port_state_out_6_2_5[2:0] ), //o
    .port_state_out_6_2_6  (shiftRows_port_state_out_6_2_6[2:0] ), //o
    .port_state_out_6_2_7  (shiftRows_port_state_out_6_2_7[2:0] ), //o
    .port_state_out_6_3_0  (shiftRows_port_state_out_6_3_0[2:0] ), //o
    .port_state_out_6_3_1  (shiftRows_port_state_out_6_3_1[2:0] ), //o
    .port_state_out_6_3_2  (shiftRows_port_state_out_6_3_2[2:0] ), //o
    .port_state_out_6_3_3  (shiftRows_port_state_out_6_3_3[2:0] ), //o
    .port_state_out_6_3_4  (shiftRows_port_state_out_6_3_4[2:0] ), //o
    .port_state_out_6_3_5  (shiftRows_port_state_out_6_3_5[2:0] ), //o
    .port_state_out_6_3_6  (shiftRows_port_state_out_6_3_6[2:0] ), //o
    .port_state_out_6_3_7  (shiftRows_port_state_out_6_3_7[2:0] ), //o
    .port_state_out_7_0_0  (shiftRows_port_state_out_7_0_0[2:0] ), //o
    .port_state_out_7_0_1  (shiftRows_port_state_out_7_0_1[2:0] ), //o
    .port_state_out_7_0_2  (shiftRows_port_state_out_7_0_2[2:0] ), //o
    .port_state_out_7_0_3  (shiftRows_port_state_out_7_0_3[2:0] ), //o
    .port_state_out_7_0_4  (shiftRows_port_state_out_7_0_4[2:0] ), //o
    .port_state_out_7_0_5  (shiftRows_port_state_out_7_0_5[2:0] ), //o
    .port_state_out_7_0_6  (shiftRows_port_state_out_7_0_6[2:0] ), //o
    .port_state_out_7_0_7  (shiftRows_port_state_out_7_0_7[2:0] ), //o
    .port_state_out_7_1_0  (shiftRows_port_state_out_7_1_0[2:0] ), //o
    .port_state_out_7_1_1  (shiftRows_port_state_out_7_1_1[2:0] ), //o
    .port_state_out_7_1_2  (shiftRows_port_state_out_7_1_2[2:0] ), //o
    .port_state_out_7_1_3  (shiftRows_port_state_out_7_1_3[2:0] ), //o
    .port_state_out_7_1_4  (shiftRows_port_state_out_7_1_4[2:0] ), //o
    .port_state_out_7_1_5  (shiftRows_port_state_out_7_1_5[2:0] ), //o
    .port_state_out_7_1_6  (shiftRows_port_state_out_7_1_6[2:0] ), //o
    .port_state_out_7_1_7  (shiftRows_port_state_out_7_1_7[2:0] ), //o
    .port_state_out_7_2_0  (shiftRows_port_state_out_7_2_0[2:0] ), //o
    .port_state_out_7_2_1  (shiftRows_port_state_out_7_2_1[2:0] ), //o
    .port_state_out_7_2_2  (shiftRows_port_state_out_7_2_2[2:0] ), //o
    .port_state_out_7_2_3  (shiftRows_port_state_out_7_2_3[2:0] ), //o
    .port_state_out_7_2_4  (shiftRows_port_state_out_7_2_4[2:0] ), //o
    .port_state_out_7_2_5  (shiftRows_port_state_out_7_2_5[2:0] ), //o
    .port_state_out_7_2_6  (shiftRows_port_state_out_7_2_6[2:0] ), //o
    .port_state_out_7_2_7  (shiftRows_port_state_out_7_2_7[2:0] ), //o
    .port_state_out_7_3_0  (shiftRows_port_state_out_7_3_0[2:0] ), //o
    .port_state_out_7_3_1  (shiftRows_port_state_out_7_3_1[2:0] ), //o
    .port_state_out_7_3_2  (shiftRows_port_state_out_7_3_2[2:0] ), //o
    .port_state_out_7_3_3  (shiftRows_port_state_out_7_3_3[2:0] ), //o
    .port_state_out_7_3_4  (shiftRows_port_state_out_7_3_4[2:0] ), //o
    .port_state_out_7_3_5  (shiftRows_port_state_out_7_3_5[2:0] ), //o
    .port_state_out_7_3_6  (shiftRows_port_state_out_7_3_6[2:0] ), //o
    .port_state_out_7_3_7  (shiftRows_port_state_out_7_3_7[2:0] ), //o
    .port_state_out_8_0_0  (shiftRows_port_state_out_8_0_0[2:0] ), //o
    .port_state_out_8_0_1  (shiftRows_port_state_out_8_0_1[2:0] ), //o
    .port_state_out_8_0_2  (shiftRows_port_state_out_8_0_2[2:0] ), //o
    .port_state_out_8_0_3  (shiftRows_port_state_out_8_0_3[2:0] ), //o
    .port_state_out_8_0_4  (shiftRows_port_state_out_8_0_4[2:0] ), //o
    .port_state_out_8_0_5  (shiftRows_port_state_out_8_0_5[2:0] ), //o
    .port_state_out_8_0_6  (shiftRows_port_state_out_8_0_6[2:0] ), //o
    .port_state_out_8_0_7  (shiftRows_port_state_out_8_0_7[2:0] ), //o
    .port_state_out_8_1_0  (shiftRows_port_state_out_8_1_0[2:0] ), //o
    .port_state_out_8_1_1  (shiftRows_port_state_out_8_1_1[2:0] ), //o
    .port_state_out_8_1_2  (shiftRows_port_state_out_8_1_2[2:0] ), //o
    .port_state_out_8_1_3  (shiftRows_port_state_out_8_1_3[2:0] ), //o
    .port_state_out_8_1_4  (shiftRows_port_state_out_8_1_4[2:0] ), //o
    .port_state_out_8_1_5  (shiftRows_port_state_out_8_1_5[2:0] ), //o
    .port_state_out_8_1_6  (shiftRows_port_state_out_8_1_6[2:0] ), //o
    .port_state_out_8_1_7  (shiftRows_port_state_out_8_1_7[2:0] ), //o
    .port_state_out_8_2_0  (shiftRows_port_state_out_8_2_0[2:0] ), //o
    .port_state_out_8_2_1  (shiftRows_port_state_out_8_2_1[2:0] ), //o
    .port_state_out_8_2_2  (shiftRows_port_state_out_8_2_2[2:0] ), //o
    .port_state_out_8_2_3  (shiftRows_port_state_out_8_2_3[2:0] ), //o
    .port_state_out_8_2_4  (shiftRows_port_state_out_8_2_4[2:0] ), //o
    .port_state_out_8_2_5  (shiftRows_port_state_out_8_2_5[2:0] ), //o
    .port_state_out_8_2_6  (shiftRows_port_state_out_8_2_6[2:0] ), //o
    .port_state_out_8_2_7  (shiftRows_port_state_out_8_2_7[2:0] ), //o
    .port_state_out_8_3_0  (shiftRows_port_state_out_8_3_0[2:0] ), //o
    .port_state_out_8_3_1  (shiftRows_port_state_out_8_3_1[2:0] ), //o
    .port_state_out_8_3_2  (shiftRows_port_state_out_8_3_2[2:0] ), //o
    .port_state_out_8_3_3  (shiftRows_port_state_out_8_3_3[2:0] ), //o
    .port_state_out_8_3_4  (shiftRows_port_state_out_8_3_4[2:0] ), //o
    .port_state_out_8_3_5  (shiftRows_port_state_out_8_3_5[2:0] ), //o
    .port_state_out_8_3_6  (shiftRows_port_state_out_8_3_6[2:0] ), //o
    .port_state_out_8_3_7  (shiftRows_port_state_out_8_3_7[2:0] ), //o
    .port_state_out_9_0_0  (shiftRows_port_state_out_9_0_0[2:0] ), //o
    .port_state_out_9_0_1  (shiftRows_port_state_out_9_0_1[2:0] ), //o
    .port_state_out_9_0_2  (shiftRows_port_state_out_9_0_2[2:0] ), //o
    .port_state_out_9_0_3  (shiftRows_port_state_out_9_0_3[2:0] ), //o
    .port_state_out_9_0_4  (shiftRows_port_state_out_9_0_4[2:0] ), //o
    .port_state_out_9_0_5  (shiftRows_port_state_out_9_0_5[2:0] ), //o
    .port_state_out_9_0_6  (shiftRows_port_state_out_9_0_6[2:0] ), //o
    .port_state_out_9_0_7  (shiftRows_port_state_out_9_0_7[2:0] ), //o
    .port_state_out_9_1_0  (shiftRows_port_state_out_9_1_0[2:0] ), //o
    .port_state_out_9_1_1  (shiftRows_port_state_out_9_1_1[2:0] ), //o
    .port_state_out_9_1_2  (shiftRows_port_state_out_9_1_2[2:0] ), //o
    .port_state_out_9_1_3  (shiftRows_port_state_out_9_1_3[2:0] ), //o
    .port_state_out_9_1_4  (shiftRows_port_state_out_9_1_4[2:0] ), //o
    .port_state_out_9_1_5  (shiftRows_port_state_out_9_1_5[2:0] ), //o
    .port_state_out_9_1_6  (shiftRows_port_state_out_9_1_6[2:0] ), //o
    .port_state_out_9_1_7  (shiftRows_port_state_out_9_1_7[2:0] ), //o
    .port_state_out_9_2_0  (shiftRows_port_state_out_9_2_0[2:0] ), //o
    .port_state_out_9_2_1  (shiftRows_port_state_out_9_2_1[2:0] ), //o
    .port_state_out_9_2_2  (shiftRows_port_state_out_9_2_2[2:0] ), //o
    .port_state_out_9_2_3  (shiftRows_port_state_out_9_2_3[2:0] ), //o
    .port_state_out_9_2_4  (shiftRows_port_state_out_9_2_4[2:0] ), //o
    .port_state_out_9_2_5  (shiftRows_port_state_out_9_2_5[2:0] ), //o
    .port_state_out_9_2_6  (shiftRows_port_state_out_9_2_6[2:0] ), //o
    .port_state_out_9_2_7  (shiftRows_port_state_out_9_2_7[2:0] ), //o
    .port_state_out_9_3_0  (shiftRows_port_state_out_9_3_0[2:0] ), //o
    .port_state_out_9_3_1  (shiftRows_port_state_out_9_3_1[2:0] ), //o
    .port_state_out_9_3_2  (shiftRows_port_state_out_9_3_2[2:0] ), //o
    .port_state_out_9_3_3  (shiftRows_port_state_out_9_3_3[2:0] ), //o
    .port_state_out_9_3_4  (shiftRows_port_state_out_9_3_4[2:0] ), //o
    .port_state_out_9_3_5  (shiftRows_port_state_out_9_3_5[2:0] ), //o
    .port_state_out_9_3_6  (shiftRows_port_state_out_9_3_6[2:0] ), //o
    .port_state_out_9_3_7  (shiftRows_port_state_out_9_3_7[2:0] ), //o
    .port_state_out_10_0_0 (shiftRows_port_state_out_10_0_0[2:0]), //o
    .port_state_out_10_0_1 (shiftRows_port_state_out_10_0_1[2:0]), //o
    .port_state_out_10_0_2 (shiftRows_port_state_out_10_0_2[2:0]), //o
    .port_state_out_10_0_3 (shiftRows_port_state_out_10_0_3[2:0]), //o
    .port_state_out_10_0_4 (shiftRows_port_state_out_10_0_4[2:0]), //o
    .port_state_out_10_0_5 (shiftRows_port_state_out_10_0_5[2:0]), //o
    .port_state_out_10_0_6 (shiftRows_port_state_out_10_0_6[2:0]), //o
    .port_state_out_10_0_7 (shiftRows_port_state_out_10_0_7[2:0]), //o
    .port_state_out_10_1_0 (shiftRows_port_state_out_10_1_0[2:0]), //o
    .port_state_out_10_1_1 (shiftRows_port_state_out_10_1_1[2:0]), //o
    .port_state_out_10_1_2 (shiftRows_port_state_out_10_1_2[2:0]), //o
    .port_state_out_10_1_3 (shiftRows_port_state_out_10_1_3[2:0]), //o
    .port_state_out_10_1_4 (shiftRows_port_state_out_10_1_4[2:0]), //o
    .port_state_out_10_1_5 (shiftRows_port_state_out_10_1_5[2:0]), //o
    .port_state_out_10_1_6 (shiftRows_port_state_out_10_1_6[2:0]), //o
    .port_state_out_10_1_7 (shiftRows_port_state_out_10_1_7[2:0]), //o
    .port_state_out_10_2_0 (shiftRows_port_state_out_10_2_0[2:0]), //o
    .port_state_out_10_2_1 (shiftRows_port_state_out_10_2_1[2:0]), //o
    .port_state_out_10_2_2 (shiftRows_port_state_out_10_2_2[2:0]), //o
    .port_state_out_10_2_3 (shiftRows_port_state_out_10_2_3[2:0]), //o
    .port_state_out_10_2_4 (shiftRows_port_state_out_10_2_4[2:0]), //o
    .port_state_out_10_2_5 (shiftRows_port_state_out_10_2_5[2:0]), //o
    .port_state_out_10_2_6 (shiftRows_port_state_out_10_2_6[2:0]), //o
    .port_state_out_10_2_7 (shiftRows_port_state_out_10_2_7[2:0]), //o
    .port_state_out_10_3_0 (shiftRows_port_state_out_10_3_0[2:0]), //o
    .port_state_out_10_3_1 (shiftRows_port_state_out_10_3_1[2:0]), //o
    .port_state_out_10_3_2 (shiftRows_port_state_out_10_3_2[2:0]), //o
    .port_state_out_10_3_3 (shiftRows_port_state_out_10_3_3[2:0]), //o
    .port_state_out_10_3_4 (shiftRows_port_state_out_10_3_4[2:0]), //o
    .port_state_out_10_3_5 (shiftRows_port_state_out_10_3_5[2:0]), //o
    .port_state_out_10_3_6 (shiftRows_port_state_out_10_3_6[2:0]), //o
    .port_state_out_10_3_7 (shiftRows_port_state_out_10_3_7[2:0]), //o
    .port_state_out_11_0_0 (shiftRows_port_state_out_11_0_0[2:0]), //o
    .port_state_out_11_0_1 (shiftRows_port_state_out_11_0_1[2:0]), //o
    .port_state_out_11_0_2 (shiftRows_port_state_out_11_0_2[2:0]), //o
    .port_state_out_11_0_3 (shiftRows_port_state_out_11_0_3[2:0]), //o
    .port_state_out_11_0_4 (shiftRows_port_state_out_11_0_4[2:0]), //o
    .port_state_out_11_0_5 (shiftRows_port_state_out_11_0_5[2:0]), //o
    .port_state_out_11_0_6 (shiftRows_port_state_out_11_0_6[2:0]), //o
    .port_state_out_11_0_7 (shiftRows_port_state_out_11_0_7[2:0]), //o
    .port_state_out_11_1_0 (shiftRows_port_state_out_11_1_0[2:0]), //o
    .port_state_out_11_1_1 (shiftRows_port_state_out_11_1_1[2:0]), //o
    .port_state_out_11_1_2 (shiftRows_port_state_out_11_1_2[2:0]), //o
    .port_state_out_11_1_3 (shiftRows_port_state_out_11_1_3[2:0]), //o
    .port_state_out_11_1_4 (shiftRows_port_state_out_11_1_4[2:0]), //o
    .port_state_out_11_1_5 (shiftRows_port_state_out_11_1_5[2:0]), //o
    .port_state_out_11_1_6 (shiftRows_port_state_out_11_1_6[2:0]), //o
    .port_state_out_11_1_7 (shiftRows_port_state_out_11_1_7[2:0]), //o
    .port_state_out_11_2_0 (shiftRows_port_state_out_11_2_0[2:0]), //o
    .port_state_out_11_2_1 (shiftRows_port_state_out_11_2_1[2:0]), //o
    .port_state_out_11_2_2 (shiftRows_port_state_out_11_2_2[2:0]), //o
    .port_state_out_11_2_3 (shiftRows_port_state_out_11_2_3[2:0]), //o
    .port_state_out_11_2_4 (shiftRows_port_state_out_11_2_4[2:0]), //o
    .port_state_out_11_2_5 (shiftRows_port_state_out_11_2_5[2:0]), //o
    .port_state_out_11_2_6 (shiftRows_port_state_out_11_2_6[2:0]), //o
    .port_state_out_11_2_7 (shiftRows_port_state_out_11_2_7[2:0]), //o
    .port_state_out_11_3_0 (shiftRows_port_state_out_11_3_0[2:0]), //o
    .port_state_out_11_3_1 (shiftRows_port_state_out_11_3_1[2:0]), //o
    .port_state_out_11_3_2 (shiftRows_port_state_out_11_3_2[2:0]), //o
    .port_state_out_11_3_3 (shiftRows_port_state_out_11_3_3[2:0]), //o
    .port_state_out_11_3_4 (shiftRows_port_state_out_11_3_4[2:0]), //o
    .port_state_out_11_3_5 (shiftRows_port_state_out_11_3_5[2:0]), //o
    .port_state_out_11_3_6 (shiftRows_port_state_out_11_3_6[2:0]), //o
    .port_state_out_11_3_7 (shiftRows_port_state_out_11_3_7[2:0]), //o
    .port_state_out_12_0_0 (shiftRows_port_state_out_12_0_0[2:0]), //o
    .port_state_out_12_0_1 (shiftRows_port_state_out_12_0_1[2:0]), //o
    .port_state_out_12_0_2 (shiftRows_port_state_out_12_0_2[2:0]), //o
    .port_state_out_12_0_3 (shiftRows_port_state_out_12_0_3[2:0]), //o
    .port_state_out_12_0_4 (shiftRows_port_state_out_12_0_4[2:0]), //o
    .port_state_out_12_0_5 (shiftRows_port_state_out_12_0_5[2:0]), //o
    .port_state_out_12_0_6 (shiftRows_port_state_out_12_0_6[2:0]), //o
    .port_state_out_12_0_7 (shiftRows_port_state_out_12_0_7[2:0]), //o
    .port_state_out_12_1_0 (shiftRows_port_state_out_12_1_0[2:0]), //o
    .port_state_out_12_1_1 (shiftRows_port_state_out_12_1_1[2:0]), //o
    .port_state_out_12_1_2 (shiftRows_port_state_out_12_1_2[2:0]), //o
    .port_state_out_12_1_3 (shiftRows_port_state_out_12_1_3[2:0]), //o
    .port_state_out_12_1_4 (shiftRows_port_state_out_12_1_4[2:0]), //o
    .port_state_out_12_1_5 (shiftRows_port_state_out_12_1_5[2:0]), //o
    .port_state_out_12_1_6 (shiftRows_port_state_out_12_1_6[2:0]), //o
    .port_state_out_12_1_7 (shiftRows_port_state_out_12_1_7[2:0]), //o
    .port_state_out_12_2_0 (shiftRows_port_state_out_12_2_0[2:0]), //o
    .port_state_out_12_2_1 (shiftRows_port_state_out_12_2_1[2:0]), //o
    .port_state_out_12_2_2 (shiftRows_port_state_out_12_2_2[2:0]), //o
    .port_state_out_12_2_3 (shiftRows_port_state_out_12_2_3[2:0]), //o
    .port_state_out_12_2_4 (shiftRows_port_state_out_12_2_4[2:0]), //o
    .port_state_out_12_2_5 (shiftRows_port_state_out_12_2_5[2:0]), //o
    .port_state_out_12_2_6 (shiftRows_port_state_out_12_2_6[2:0]), //o
    .port_state_out_12_2_7 (shiftRows_port_state_out_12_2_7[2:0]), //o
    .port_state_out_12_3_0 (shiftRows_port_state_out_12_3_0[2:0]), //o
    .port_state_out_12_3_1 (shiftRows_port_state_out_12_3_1[2:0]), //o
    .port_state_out_12_3_2 (shiftRows_port_state_out_12_3_2[2:0]), //o
    .port_state_out_12_3_3 (shiftRows_port_state_out_12_3_3[2:0]), //o
    .port_state_out_12_3_4 (shiftRows_port_state_out_12_3_4[2:0]), //o
    .port_state_out_12_3_5 (shiftRows_port_state_out_12_3_5[2:0]), //o
    .port_state_out_12_3_6 (shiftRows_port_state_out_12_3_6[2:0]), //o
    .port_state_out_12_3_7 (shiftRows_port_state_out_12_3_7[2:0]), //o
    .port_state_out_13_0_0 (shiftRows_port_state_out_13_0_0[2:0]), //o
    .port_state_out_13_0_1 (shiftRows_port_state_out_13_0_1[2:0]), //o
    .port_state_out_13_0_2 (shiftRows_port_state_out_13_0_2[2:0]), //o
    .port_state_out_13_0_3 (shiftRows_port_state_out_13_0_3[2:0]), //o
    .port_state_out_13_0_4 (shiftRows_port_state_out_13_0_4[2:0]), //o
    .port_state_out_13_0_5 (shiftRows_port_state_out_13_0_5[2:0]), //o
    .port_state_out_13_0_6 (shiftRows_port_state_out_13_0_6[2:0]), //o
    .port_state_out_13_0_7 (shiftRows_port_state_out_13_0_7[2:0]), //o
    .port_state_out_13_1_0 (shiftRows_port_state_out_13_1_0[2:0]), //o
    .port_state_out_13_1_1 (shiftRows_port_state_out_13_1_1[2:0]), //o
    .port_state_out_13_1_2 (shiftRows_port_state_out_13_1_2[2:0]), //o
    .port_state_out_13_1_3 (shiftRows_port_state_out_13_1_3[2:0]), //o
    .port_state_out_13_1_4 (shiftRows_port_state_out_13_1_4[2:0]), //o
    .port_state_out_13_1_5 (shiftRows_port_state_out_13_1_5[2:0]), //o
    .port_state_out_13_1_6 (shiftRows_port_state_out_13_1_6[2:0]), //o
    .port_state_out_13_1_7 (shiftRows_port_state_out_13_1_7[2:0]), //o
    .port_state_out_13_2_0 (shiftRows_port_state_out_13_2_0[2:0]), //o
    .port_state_out_13_2_1 (shiftRows_port_state_out_13_2_1[2:0]), //o
    .port_state_out_13_2_2 (shiftRows_port_state_out_13_2_2[2:0]), //o
    .port_state_out_13_2_3 (shiftRows_port_state_out_13_2_3[2:0]), //o
    .port_state_out_13_2_4 (shiftRows_port_state_out_13_2_4[2:0]), //o
    .port_state_out_13_2_5 (shiftRows_port_state_out_13_2_5[2:0]), //o
    .port_state_out_13_2_6 (shiftRows_port_state_out_13_2_6[2:0]), //o
    .port_state_out_13_2_7 (shiftRows_port_state_out_13_2_7[2:0]), //o
    .port_state_out_13_3_0 (shiftRows_port_state_out_13_3_0[2:0]), //o
    .port_state_out_13_3_1 (shiftRows_port_state_out_13_3_1[2:0]), //o
    .port_state_out_13_3_2 (shiftRows_port_state_out_13_3_2[2:0]), //o
    .port_state_out_13_3_3 (shiftRows_port_state_out_13_3_3[2:0]), //o
    .port_state_out_13_3_4 (shiftRows_port_state_out_13_3_4[2:0]), //o
    .port_state_out_13_3_5 (shiftRows_port_state_out_13_3_5[2:0]), //o
    .port_state_out_13_3_6 (shiftRows_port_state_out_13_3_6[2:0]), //o
    .port_state_out_13_3_7 (shiftRows_port_state_out_13_3_7[2:0]), //o
    .port_state_out_14_0_0 (shiftRows_port_state_out_14_0_0[2:0]), //o
    .port_state_out_14_0_1 (shiftRows_port_state_out_14_0_1[2:0]), //o
    .port_state_out_14_0_2 (shiftRows_port_state_out_14_0_2[2:0]), //o
    .port_state_out_14_0_3 (shiftRows_port_state_out_14_0_3[2:0]), //o
    .port_state_out_14_0_4 (shiftRows_port_state_out_14_0_4[2:0]), //o
    .port_state_out_14_0_5 (shiftRows_port_state_out_14_0_5[2:0]), //o
    .port_state_out_14_0_6 (shiftRows_port_state_out_14_0_6[2:0]), //o
    .port_state_out_14_0_7 (shiftRows_port_state_out_14_0_7[2:0]), //o
    .port_state_out_14_1_0 (shiftRows_port_state_out_14_1_0[2:0]), //o
    .port_state_out_14_1_1 (shiftRows_port_state_out_14_1_1[2:0]), //o
    .port_state_out_14_1_2 (shiftRows_port_state_out_14_1_2[2:0]), //o
    .port_state_out_14_1_3 (shiftRows_port_state_out_14_1_3[2:0]), //o
    .port_state_out_14_1_4 (shiftRows_port_state_out_14_1_4[2:0]), //o
    .port_state_out_14_1_5 (shiftRows_port_state_out_14_1_5[2:0]), //o
    .port_state_out_14_1_6 (shiftRows_port_state_out_14_1_6[2:0]), //o
    .port_state_out_14_1_7 (shiftRows_port_state_out_14_1_7[2:0]), //o
    .port_state_out_14_2_0 (shiftRows_port_state_out_14_2_0[2:0]), //o
    .port_state_out_14_2_1 (shiftRows_port_state_out_14_2_1[2:0]), //o
    .port_state_out_14_2_2 (shiftRows_port_state_out_14_2_2[2:0]), //o
    .port_state_out_14_2_3 (shiftRows_port_state_out_14_2_3[2:0]), //o
    .port_state_out_14_2_4 (shiftRows_port_state_out_14_2_4[2:0]), //o
    .port_state_out_14_2_5 (shiftRows_port_state_out_14_2_5[2:0]), //o
    .port_state_out_14_2_6 (shiftRows_port_state_out_14_2_6[2:0]), //o
    .port_state_out_14_2_7 (shiftRows_port_state_out_14_2_7[2:0]), //o
    .port_state_out_14_3_0 (shiftRows_port_state_out_14_3_0[2:0]), //o
    .port_state_out_14_3_1 (shiftRows_port_state_out_14_3_1[2:0]), //o
    .port_state_out_14_3_2 (shiftRows_port_state_out_14_3_2[2:0]), //o
    .port_state_out_14_3_3 (shiftRows_port_state_out_14_3_3[2:0]), //o
    .port_state_out_14_3_4 (shiftRows_port_state_out_14_3_4[2:0]), //o
    .port_state_out_14_3_5 (shiftRows_port_state_out_14_3_5[2:0]), //o
    .port_state_out_14_3_6 (shiftRows_port_state_out_14_3_6[2:0]), //o
    .port_state_out_14_3_7 (shiftRows_port_state_out_14_3_7[2:0]), //o
    .port_state_out_15_0_0 (shiftRows_port_state_out_15_0_0[2:0]), //o
    .port_state_out_15_0_1 (shiftRows_port_state_out_15_0_1[2:0]), //o
    .port_state_out_15_0_2 (shiftRows_port_state_out_15_0_2[2:0]), //o
    .port_state_out_15_0_3 (shiftRows_port_state_out_15_0_3[2:0]), //o
    .port_state_out_15_0_4 (shiftRows_port_state_out_15_0_4[2:0]), //o
    .port_state_out_15_0_5 (shiftRows_port_state_out_15_0_5[2:0]), //o
    .port_state_out_15_0_6 (shiftRows_port_state_out_15_0_6[2:0]), //o
    .port_state_out_15_0_7 (shiftRows_port_state_out_15_0_7[2:0]), //o
    .port_state_out_15_1_0 (shiftRows_port_state_out_15_1_0[2:0]), //o
    .port_state_out_15_1_1 (shiftRows_port_state_out_15_1_1[2:0]), //o
    .port_state_out_15_1_2 (shiftRows_port_state_out_15_1_2[2:0]), //o
    .port_state_out_15_1_3 (shiftRows_port_state_out_15_1_3[2:0]), //o
    .port_state_out_15_1_4 (shiftRows_port_state_out_15_1_4[2:0]), //o
    .port_state_out_15_1_5 (shiftRows_port_state_out_15_1_5[2:0]), //o
    .port_state_out_15_1_6 (shiftRows_port_state_out_15_1_6[2:0]), //o
    .port_state_out_15_1_7 (shiftRows_port_state_out_15_1_7[2:0]), //o
    .port_state_out_15_2_0 (shiftRows_port_state_out_15_2_0[2:0]), //o
    .port_state_out_15_2_1 (shiftRows_port_state_out_15_2_1[2:0]), //o
    .port_state_out_15_2_2 (shiftRows_port_state_out_15_2_2[2:0]), //o
    .port_state_out_15_2_3 (shiftRows_port_state_out_15_2_3[2:0]), //o
    .port_state_out_15_2_4 (shiftRows_port_state_out_15_2_4[2:0]), //o
    .port_state_out_15_2_5 (shiftRows_port_state_out_15_2_5[2:0]), //o
    .port_state_out_15_2_6 (shiftRows_port_state_out_15_2_6[2:0]), //o
    .port_state_out_15_2_7 (shiftRows_port_state_out_15_2_7[2:0]), //o
    .port_state_out_15_3_0 (shiftRows_port_state_out_15_3_0[2:0]), //o
    .port_state_out_15_3_1 (shiftRows_port_state_out_15_3_1[2:0]), //o
    .port_state_out_15_3_2 (shiftRows_port_state_out_15_3_2[2:0]), //o
    .port_state_out_15_3_3 (shiftRows_port_state_out_15_3_3[2:0]), //o
    .port_state_out_15_3_4 (shiftRows_port_state_out_15_3_4[2:0]), //o
    .port_state_out_15_3_5 (shiftRows_port_state_out_15_3_5[2:0]), //o
    .port_state_out_15_3_6 (shiftRows_port_state_out_15_3_6[2:0]), //o
    .port_state_out_15_3_7 (shiftRows_port_state_out_15_3_7[2:0])  //o
  );
  Aes_MixColumn mixColumns (
    .port_state_in_0_0_0   (shiftRows_port_state_out_0_0_0[2:0]  ), //i
    .port_state_in_0_0_1   (shiftRows_port_state_out_0_0_1[2:0]  ), //i
    .port_state_in_0_0_2   (shiftRows_port_state_out_0_0_2[2:0]  ), //i
    .port_state_in_0_0_3   (shiftRows_port_state_out_0_0_3[2:0]  ), //i
    .port_state_in_0_0_4   (shiftRows_port_state_out_0_0_4[2:0]  ), //i
    .port_state_in_0_0_5   (shiftRows_port_state_out_0_0_5[2:0]  ), //i
    .port_state_in_0_0_6   (shiftRows_port_state_out_0_0_6[2:0]  ), //i
    .port_state_in_0_0_7   (shiftRows_port_state_out_0_0_7[2:0]  ), //i
    .port_state_in_0_1_0   (shiftRows_port_state_out_0_1_0[2:0]  ), //i
    .port_state_in_0_1_1   (shiftRows_port_state_out_0_1_1[2:0]  ), //i
    .port_state_in_0_1_2   (shiftRows_port_state_out_0_1_2[2:0]  ), //i
    .port_state_in_0_1_3   (shiftRows_port_state_out_0_1_3[2:0]  ), //i
    .port_state_in_0_1_4   (shiftRows_port_state_out_0_1_4[2:0]  ), //i
    .port_state_in_0_1_5   (shiftRows_port_state_out_0_1_5[2:0]  ), //i
    .port_state_in_0_1_6   (shiftRows_port_state_out_0_1_6[2:0]  ), //i
    .port_state_in_0_1_7   (shiftRows_port_state_out_0_1_7[2:0]  ), //i
    .port_state_in_0_2_0   (shiftRows_port_state_out_0_2_0[2:0]  ), //i
    .port_state_in_0_2_1   (shiftRows_port_state_out_0_2_1[2:0]  ), //i
    .port_state_in_0_2_2   (shiftRows_port_state_out_0_2_2[2:0]  ), //i
    .port_state_in_0_2_3   (shiftRows_port_state_out_0_2_3[2:0]  ), //i
    .port_state_in_0_2_4   (shiftRows_port_state_out_0_2_4[2:0]  ), //i
    .port_state_in_0_2_5   (shiftRows_port_state_out_0_2_5[2:0]  ), //i
    .port_state_in_0_2_6   (shiftRows_port_state_out_0_2_6[2:0]  ), //i
    .port_state_in_0_2_7   (shiftRows_port_state_out_0_2_7[2:0]  ), //i
    .port_state_in_0_3_0   (shiftRows_port_state_out_0_3_0[2:0]  ), //i
    .port_state_in_0_3_1   (shiftRows_port_state_out_0_3_1[2:0]  ), //i
    .port_state_in_0_3_2   (shiftRows_port_state_out_0_3_2[2:0]  ), //i
    .port_state_in_0_3_3   (shiftRows_port_state_out_0_3_3[2:0]  ), //i
    .port_state_in_0_3_4   (shiftRows_port_state_out_0_3_4[2:0]  ), //i
    .port_state_in_0_3_5   (shiftRows_port_state_out_0_3_5[2:0]  ), //i
    .port_state_in_0_3_6   (shiftRows_port_state_out_0_3_6[2:0]  ), //i
    .port_state_in_0_3_7   (shiftRows_port_state_out_0_3_7[2:0]  ), //i
    .port_state_in_1_0_0   (shiftRows_port_state_out_1_0_0[2:0]  ), //i
    .port_state_in_1_0_1   (shiftRows_port_state_out_1_0_1[2:0]  ), //i
    .port_state_in_1_0_2   (shiftRows_port_state_out_1_0_2[2:0]  ), //i
    .port_state_in_1_0_3   (shiftRows_port_state_out_1_0_3[2:0]  ), //i
    .port_state_in_1_0_4   (shiftRows_port_state_out_1_0_4[2:0]  ), //i
    .port_state_in_1_0_5   (shiftRows_port_state_out_1_0_5[2:0]  ), //i
    .port_state_in_1_0_6   (shiftRows_port_state_out_1_0_6[2:0]  ), //i
    .port_state_in_1_0_7   (shiftRows_port_state_out_1_0_7[2:0]  ), //i
    .port_state_in_1_1_0   (shiftRows_port_state_out_1_1_0[2:0]  ), //i
    .port_state_in_1_1_1   (shiftRows_port_state_out_1_1_1[2:0]  ), //i
    .port_state_in_1_1_2   (shiftRows_port_state_out_1_1_2[2:0]  ), //i
    .port_state_in_1_1_3   (shiftRows_port_state_out_1_1_3[2:0]  ), //i
    .port_state_in_1_1_4   (shiftRows_port_state_out_1_1_4[2:0]  ), //i
    .port_state_in_1_1_5   (shiftRows_port_state_out_1_1_5[2:0]  ), //i
    .port_state_in_1_1_6   (shiftRows_port_state_out_1_1_6[2:0]  ), //i
    .port_state_in_1_1_7   (shiftRows_port_state_out_1_1_7[2:0]  ), //i
    .port_state_in_1_2_0   (shiftRows_port_state_out_1_2_0[2:0]  ), //i
    .port_state_in_1_2_1   (shiftRows_port_state_out_1_2_1[2:0]  ), //i
    .port_state_in_1_2_2   (shiftRows_port_state_out_1_2_2[2:0]  ), //i
    .port_state_in_1_2_3   (shiftRows_port_state_out_1_2_3[2:0]  ), //i
    .port_state_in_1_2_4   (shiftRows_port_state_out_1_2_4[2:0]  ), //i
    .port_state_in_1_2_5   (shiftRows_port_state_out_1_2_5[2:0]  ), //i
    .port_state_in_1_2_6   (shiftRows_port_state_out_1_2_6[2:0]  ), //i
    .port_state_in_1_2_7   (shiftRows_port_state_out_1_2_7[2:0]  ), //i
    .port_state_in_1_3_0   (shiftRows_port_state_out_1_3_0[2:0]  ), //i
    .port_state_in_1_3_1   (shiftRows_port_state_out_1_3_1[2:0]  ), //i
    .port_state_in_1_3_2   (shiftRows_port_state_out_1_3_2[2:0]  ), //i
    .port_state_in_1_3_3   (shiftRows_port_state_out_1_3_3[2:0]  ), //i
    .port_state_in_1_3_4   (shiftRows_port_state_out_1_3_4[2:0]  ), //i
    .port_state_in_1_3_5   (shiftRows_port_state_out_1_3_5[2:0]  ), //i
    .port_state_in_1_3_6   (shiftRows_port_state_out_1_3_6[2:0]  ), //i
    .port_state_in_1_3_7   (shiftRows_port_state_out_1_3_7[2:0]  ), //i
    .port_state_in_2_0_0   (shiftRows_port_state_out_2_0_0[2:0]  ), //i
    .port_state_in_2_0_1   (shiftRows_port_state_out_2_0_1[2:0]  ), //i
    .port_state_in_2_0_2   (shiftRows_port_state_out_2_0_2[2:0]  ), //i
    .port_state_in_2_0_3   (shiftRows_port_state_out_2_0_3[2:0]  ), //i
    .port_state_in_2_0_4   (shiftRows_port_state_out_2_0_4[2:0]  ), //i
    .port_state_in_2_0_5   (shiftRows_port_state_out_2_0_5[2:0]  ), //i
    .port_state_in_2_0_6   (shiftRows_port_state_out_2_0_6[2:0]  ), //i
    .port_state_in_2_0_7   (shiftRows_port_state_out_2_0_7[2:0]  ), //i
    .port_state_in_2_1_0   (shiftRows_port_state_out_2_1_0[2:0]  ), //i
    .port_state_in_2_1_1   (shiftRows_port_state_out_2_1_1[2:0]  ), //i
    .port_state_in_2_1_2   (shiftRows_port_state_out_2_1_2[2:0]  ), //i
    .port_state_in_2_1_3   (shiftRows_port_state_out_2_1_3[2:0]  ), //i
    .port_state_in_2_1_4   (shiftRows_port_state_out_2_1_4[2:0]  ), //i
    .port_state_in_2_1_5   (shiftRows_port_state_out_2_1_5[2:0]  ), //i
    .port_state_in_2_1_6   (shiftRows_port_state_out_2_1_6[2:0]  ), //i
    .port_state_in_2_1_7   (shiftRows_port_state_out_2_1_7[2:0]  ), //i
    .port_state_in_2_2_0   (shiftRows_port_state_out_2_2_0[2:0]  ), //i
    .port_state_in_2_2_1   (shiftRows_port_state_out_2_2_1[2:0]  ), //i
    .port_state_in_2_2_2   (shiftRows_port_state_out_2_2_2[2:0]  ), //i
    .port_state_in_2_2_3   (shiftRows_port_state_out_2_2_3[2:0]  ), //i
    .port_state_in_2_2_4   (shiftRows_port_state_out_2_2_4[2:0]  ), //i
    .port_state_in_2_2_5   (shiftRows_port_state_out_2_2_5[2:0]  ), //i
    .port_state_in_2_2_6   (shiftRows_port_state_out_2_2_6[2:0]  ), //i
    .port_state_in_2_2_7   (shiftRows_port_state_out_2_2_7[2:0]  ), //i
    .port_state_in_2_3_0   (shiftRows_port_state_out_2_3_0[2:0]  ), //i
    .port_state_in_2_3_1   (shiftRows_port_state_out_2_3_1[2:0]  ), //i
    .port_state_in_2_3_2   (shiftRows_port_state_out_2_3_2[2:0]  ), //i
    .port_state_in_2_3_3   (shiftRows_port_state_out_2_3_3[2:0]  ), //i
    .port_state_in_2_3_4   (shiftRows_port_state_out_2_3_4[2:0]  ), //i
    .port_state_in_2_3_5   (shiftRows_port_state_out_2_3_5[2:0]  ), //i
    .port_state_in_2_3_6   (shiftRows_port_state_out_2_3_6[2:0]  ), //i
    .port_state_in_2_3_7   (shiftRows_port_state_out_2_3_7[2:0]  ), //i
    .port_state_in_3_0_0   (shiftRows_port_state_out_3_0_0[2:0]  ), //i
    .port_state_in_3_0_1   (shiftRows_port_state_out_3_0_1[2:0]  ), //i
    .port_state_in_3_0_2   (shiftRows_port_state_out_3_0_2[2:0]  ), //i
    .port_state_in_3_0_3   (shiftRows_port_state_out_3_0_3[2:0]  ), //i
    .port_state_in_3_0_4   (shiftRows_port_state_out_3_0_4[2:0]  ), //i
    .port_state_in_3_0_5   (shiftRows_port_state_out_3_0_5[2:0]  ), //i
    .port_state_in_3_0_6   (shiftRows_port_state_out_3_0_6[2:0]  ), //i
    .port_state_in_3_0_7   (shiftRows_port_state_out_3_0_7[2:0]  ), //i
    .port_state_in_3_1_0   (shiftRows_port_state_out_3_1_0[2:0]  ), //i
    .port_state_in_3_1_1   (shiftRows_port_state_out_3_1_1[2:0]  ), //i
    .port_state_in_3_1_2   (shiftRows_port_state_out_3_1_2[2:0]  ), //i
    .port_state_in_3_1_3   (shiftRows_port_state_out_3_1_3[2:0]  ), //i
    .port_state_in_3_1_4   (shiftRows_port_state_out_3_1_4[2:0]  ), //i
    .port_state_in_3_1_5   (shiftRows_port_state_out_3_1_5[2:0]  ), //i
    .port_state_in_3_1_6   (shiftRows_port_state_out_3_1_6[2:0]  ), //i
    .port_state_in_3_1_7   (shiftRows_port_state_out_3_1_7[2:0]  ), //i
    .port_state_in_3_2_0   (shiftRows_port_state_out_3_2_0[2:0]  ), //i
    .port_state_in_3_2_1   (shiftRows_port_state_out_3_2_1[2:0]  ), //i
    .port_state_in_3_2_2   (shiftRows_port_state_out_3_2_2[2:0]  ), //i
    .port_state_in_3_2_3   (shiftRows_port_state_out_3_2_3[2:0]  ), //i
    .port_state_in_3_2_4   (shiftRows_port_state_out_3_2_4[2:0]  ), //i
    .port_state_in_3_2_5   (shiftRows_port_state_out_3_2_5[2:0]  ), //i
    .port_state_in_3_2_6   (shiftRows_port_state_out_3_2_6[2:0]  ), //i
    .port_state_in_3_2_7   (shiftRows_port_state_out_3_2_7[2:0]  ), //i
    .port_state_in_3_3_0   (shiftRows_port_state_out_3_3_0[2:0]  ), //i
    .port_state_in_3_3_1   (shiftRows_port_state_out_3_3_1[2:0]  ), //i
    .port_state_in_3_3_2   (shiftRows_port_state_out_3_3_2[2:0]  ), //i
    .port_state_in_3_3_3   (shiftRows_port_state_out_3_3_3[2:0]  ), //i
    .port_state_in_3_3_4   (shiftRows_port_state_out_3_3_4[2:0]  ), //i
    .port_state_in_3_3_5   (shiftRows_port_state_out_3_3_5[2:0]  ), //i
    .port_state_in_3_3_6   (shiftRows_port_state_out_3_3_6[2:0]  ), //i
    .port_state_in_3_3_7   (shiftRows_port_state_out_3_3_7[2:0]  ), //i
    .port_state_in_4_0_0   (shiftRows_port_state_out_4_0_0[2:0]  ), //i
    .port_state_in_4_0_1   (shiftRows_port_state_out_4_0_1[2:0]  ), //i
    .port_state_in_4_0_2   (shiftRows_port_state_out_4_0_2[2:0]  ), //i
    .port_state_in_4_0_3   (shiftRows_port_state_out_4_0_3[2:0]  ), //i
    .port_state_in_4_0_4   (shiftRows_port_state_out_4_0_4[2:0]  ), //i
    .port_state_in_4_0_5   (shiftRows_port_state_out_4_0_5[2:0]  ), //i
    .port_state_in_4_0_6   (shiftRows_port_state_out_4_0_6[2:0]  ), //i
    .port_state_in_4_0_7   (shiftRows_port_state_out_4_0_7[2:0]  ), //i
    .port_state_in_4_1_0   (shiftRows_port_state_out_4_1_0[2:0]  ), //i
    .port_state_in_4_1_1   (shiftRows_port_state_out_4_1_1[2:0]  ), //i
    .port_state_in_4_1_2   (shiftRows_port_state_out_4_1_2[2:0]  ), //i
    .port_state_in_4_1_3   (shiftRows_port_state_out_4_1_3[2:0]  ), //i
    .port_state_in_4_1_4   (shiftRows_port_state_out_4_1_4[2:0]  ), //i
    .port_state_in_4_1_5   (shiftRows_port_state_out_4_1_5[2:0]  ), //i
    .port_state_in_4_1_6   (shiftRows_port_state_out_4_1_6[2:0]  ), //i
    .port_state_in_4_1_7   (shiftRows_port_state_out_4_1_7[2:0]  ), //i
    .port_state_in_4_2_0   (shiftRows_port_state_out_4_2_0[2:0]  ), //i
    .port_state_in_4_2_1   (shiftRows_port_state_out_4_2_1[2:0]  ), //i
    .port_state_in_4_2_2   (shiftRows_port_state_out_4_2_2[2:0]  ), //i
    .port_state_in_4_2_3   (shiftRows_port_state_out_4_2_3[2:0]  ), //i
    .port_state_in_4_2_4   (shiftRows_port_state_out_4_2_4[2:0]  ), //i
    .port_state_in_4_2_5   (shiftRows_port_state_out_4_2_5[2:0]  ), //i
    .port_state_in_4_2_6   (shiftRows_port_state_out_4_2_6[2:0]  ), //i
    .port_state_in_4_2_7   (shiftRows_port_state_out_4_2_7[2:0]  ), //i
    .port_state_in_4_3_0   (shiftRows_port_state_out_4_3_0[2:0]  ), //i
    .port_state_in_4_3_1   (shiftRows_port_state_out_4_3_1[2:0]  ), //i
    .port_state_in_4_3_2   (shiftRows_port_state_out_4_3_2[2:0]  ), //i
    .port_state_in_4_3_3   (shiftRows_port_state_out_4_3_3[2:0]  ), //i
    .port_state_in_4_3_4   (shiftRows_port_state_out_4_3_4[2:0]  ), //i
    .port_state_in_4_3_5   (shiftRows_port_state_out_4_3_5[2:0]  ), //i
    .port_state_in_4_3_6   (shiftRows_port_state_out_4_3_6[2:0]  ), //i
    .port_state_in_4_3_7   (shiftRows_port_state_out_4_3_7[2:0]  ), //i
    .port_state_in_5_0_0   (shiftRows_port_state_out_5_0_0[2:0]  ), //i
    .port_state_in_5_0_1   (shiftRows_port_state_out_5_0_1[2:0]  ), //i
    .port_state_in_5_0_2   (shiftRows_port_state_out_5_0_2[2:0]  ), //i
    .port_state_in_5_0_3   (shiftRows_port_state_out_5_0_3[2:0]  ), //i
    .port_state_in_5_0_4   (shiftRows_port_state_out_5_0_4[2:0]  ), //i
    .port_state_in_5_0_5   (shiftRows_port_state_out_5_0_5[2:0]  ), //i
    .port_state_in_5_0_6   (shiftRows_port_state_out_5_0_6[2:0]  ), //i
    .port_state_in_5_0_7   (shiftRows_port_state_out_5_0_7[2:0]  ), //i
    .port_state_in_5_1_0   (shiftRows_port_state_out_5_1_0[2:0]  ), //i
    .port_state_in_5_1_1   (shiftRows_port_state_out_5_1_1[2:0]  ), //i
    .port_state_in_5_1_2   (shiftRows_port_state_out_5_1_2[2:0]  ), //i
    .port_state_in_5_1_3   (shiftRows_port_state_out_5_1_3[2:0]  ), //i
    .port_state_in_5_1_4   (shiftRows_port_state_out_5_1_4[2:0]  ), //i
    .port_state_in_5_1_5   (shiftRows_port_state_out_5_1_5[2:0]  ), //i
    .port_state_in_5_1_6   (shiftRows_port_state_out_5_1_6[2:0]  ), //i
    .port_state_in_5_1_7   (shiftRows_port_state_out_5_1_7[2:0]  ), //i
    .port_state_in_5_2_0   (shiftRows_port_state_out_5_2_0[2:0]  ), //i
    .port_state_in_5_2_1   (shiftRows_port_state_out_5_2_1[2:0]  ), //i
    .port_state_in_5_2_2   (shiftRows_port_state_out_5_2_2[2:0]  ), //i
    .port_state_in_5_2_3   (shiftRows_port_state_out_5_2_3[2:0]  ), //i
    .port_state_in_5_2_4   (shiftRows_port_state_out_5_2_4[2:0]  ), //i
    .port_state_in_5_2_5   (shiftRows_port_state_out_5_2_5[2:0]  ), //i
    .port_state_in_5_2_6   (shiftRows_port_state_out_5_2_6[2:0]  ), //i
    .port_state_in_5_2_7   (shiftRows_port_state_out_5_2_7[2:0]  ), //i
    .port_state_in_5_3_0   (shiftRows_port_state_out_5_3_0[2:0]  ), //i
    .port_state_in_5_3_1   (shiftRows_port_state_out_5_3_1[2:0]  ), //i
    .port_state_in_5_3_2   (shiftRows_port_state_out_5_3_2[2:0]  ), //i
    .port_state_in_5_3_3   (shiftRows_port_state_out_5_3_3[2:0]  ), //i
    .port_state_in_5_3_4   (shiftRows_port_state_out_5_3_4[2:0]  ), //i
    .port_state_in_5_3_5   (shiftRows_port_state_out_5_3_5[2:0]  ), //i
    .port_state_in_5_3_6   (shiftRows_port_state_out_5_3_6[2:0]  ), //i
    .port_state_in_5_3_7   (shiftRows_port_state_out_5_3_7[2:0]  ), //i
    .port_state_in_6_0_0   (shiftRows_port_state_out_6_0_0[2:0]  ), //i
    .port_state_in_6_0_1   (shiftRows_port_state_out_6_0_1[2:0]  ), //i
    .port_state_in_6_0_2   (shiftRows_port_state_out_6_0_2[2:0]  ), //i
    .port_state_in_6_0_3   (shiftRows_port_state_out_6_0_3[2:0]  ), //i
    .port_state_in_6_0_4   (shiftRows_port_state_out_6_0_4[2:0]  ), //i
    .port_state_in_6_0_5   (shiftRows_port_state_out_6_0_5[2:0]  ), //i
    .port_state_in_6_0_6   (shiftRows_port_state_out_6_0_6[2:0]  ), //i
    .port_state_in_6_0_7   (shiftRows_port_state_out_6_0_7[2:0]  ), //i
    .port_state_in_6_1_0   (shiftRows_port_state_out_6_1_0[2:0]  ), //i
    .port_state_in_6_1_1   (shiftRows_port_state_out_6_1_1[2:0]  ), //i
    .port_state_in_6_1_2   (shiftRows_port_state_out_6_1_2[2:0]  ), //i
    .port_state_in_6_1_3   (shiftRows_port_state_out_6_1_3[2:0]  ), //i
    .port_state_in_6_1_4   (shiftRows_port_state_out_6_1_4[2:0]  ), //i
    .port_state_in_6_1_5   (shiftRows_port_state_out_6_1_5[2:0]  ), //i
    .port_state_in_6_1_6   (shiftRows_port_state_out_6_1_6[2:0]  ), //i
    .port_state_in_6_1_7   (shiftRows_port_state_out_6_1_7[2:0]  ), //i
    .port_state_in_6_2_0   (shiftRows_port_state_out_6_2_0[2:0]  ), //i
    .port_state_in_6_2_1   (shiftRows_port_state_out_6_2_1[2:0]  ), //i
    .port_state_in_6_2_2   (shiftRows_port_state_out_6_2_2[2:0]  ), //i
    .port_state_in_6_2_3   (shiftRows_port_state_out_6_2_3[2:0]  ), //i
    .port_state_in_6_2_4   (shiftRows_port_state_out_6_2_4[2:0]  ), //i
    .port_state_in_6_2_5   (shiftRows_port_state_out_6_2_5[2:0]  ), //i
    .port_state_in_6_2_6   (shiftRows_port_state_out_6_2_6[2:0]  ), //i
    .port_state_in_6_2_7   (shiftRows_port_state_out_6_2_7[2:0]  ), //i
    .port_state_in_6_3_0   (shiftRows_port_state_out_6_3_0[2:0]  ), //i
    .port_state_in_6_3_1   (shiftRows_port_state_out_6_3_1[2:0]  ), //i
    .port_state_in_6_3_2   (shiftRows_port_state_out_6_3_2[2:0]  ), //i
    .port_state_in_6_3_3   (shiftRows_port_state_out_6_3_3[2:0]  ), //i
    .port_state_in_6_3_4   (shiftRows_port_state_out_6_3_4[2:0]  ), //i
    .port_state_in_6_3_5   (shiftRows_port_state_out_6_3_5[2:0]  ), //i
    .port_state_in_6_3_6   (shiftRows_port_state_out_6_3_6[2:0]  ), //i
    .port_state_in_6_3_7   (shiftRows_port_state_out_6_3_7[2:0]  ), //i
    .port_state_in_7_0_0   (shiftRows_port_state_out_7_0_0[2:0]  ), //i
    .port_state_in_7_0_1   (shiftRows_port_state_out_7_0_1[2:0]  ), //i
    .port_state_in_7_0_2   (shiftRows_port_state_out_7_0_2[2:0]  ), //i
    .port_state_in_7_0_3   (shiftRows_port_state_out_7_0_3[2:0]  ), //i
    .port_state_in_7_0_4   (shiftRows_port_state_out_7_0_4[2:0]  ), //i
    .port_state_in_7_0_5   (shiftRows_port_state_out_7_0_5[2:0]  ), //i
    .port_state_in_7_0_6   (shiftRows_port_state_out_7_0_6[2:0]  ), //i
    .port_state_in_7_0_7   (shiftRows_port_state_out_7_0_7[2:0]  ), //i
    .port_state_in_7_1_0   (shiftRows_port_state_out_7_1_0[2:0]  ), //i
    .port_state_in_7_1_1   (shiftRows_port_state_out_7_1_1[2:0]  ), //i
    .port_state_in_7_1_2   (shiftRows_port_state_out_7_1_2[2:0]  ), //i
    .port_state_in_7_1_3   (shiftRows_port_state_out_7_1_3[2:0]  ), //i
    .port_state_in_7_1_4   (shiftRows_port_state_out_7_1_4[2:0]  ), //i
    .port_state_in_7_1_5   (shiftRows_port_state_out_7_1_5[2:0]  ), //i
    .port_state_in_7_1_6   (shiftRows_port_state_out_7_1_6[2:0]  ), //i
    .port_state_in_7_1_7   (shiftRows_port_state_out_7_1_7[2:0]  ), //i
    .port_state_in_7_2_0   (shiftRows_port_state_out_7_2_0[2:0]  ), //i
    .port_state_in_7_2_1   (shiftRows_port_state_out_7_2_1[2:0]  ), //i
    .port_state_in_7_2_2   (shiftRows_port_state_out_7_2_2[2:0]  ), //i
    .port_state_in_7_2_3   (shiftRows_port_state_out_7_2_3[2:0]  ), //i
    .port_state_in_7_2_4   (shiftRows_port_state_out_7_2_4[2:0]  ), //i
    .port_state_in_7_2_5   (shiftRows_port_state_out_7_2_5[2:0]  ), //i
    .port_state_in_7_2_6   (shiftRows_port_state_out_7_2_6[2:0]  ), //i
    .port_state_in_7_2_7   (shiftRows_port_state_out_7_2_7[2:0]  ), //i
    .port_state_in_7_3_0   (shiftRows_port_state_out_7_3_0[2:0]  ), //i
    .port_state_in_7_3_1   (shiftRows_port_state_out_7_3_1[2:0]  ), //i
    .port_state_in_7_3_2   (shiftRows_port_state_out_7_3_2[2:0]  ), //i
    .port_state_in_7_3_3   (shiftRows_port_state_out_7_3_3[2:0]  ), //i
    .port_state_in_7_3_4   (shiftRows_port_state_out_7_3_4[2:0]  ), //i
    .port_state_in_7_3_5   (shiftRows_port_state_out_7_3_5[2:0]  ), //i
    .port_state_in_7_3_6   (shiftRows_port_state_out_7_3_6[2:0]  ), //i
    .port_state_in_7_3_7   (shiftRows_port_state_out_7_3_7[2:0]  ), //i
    .port_state_in_8_0_0   (shiftRows_port_state_out_8_0_0[2:0]  ), //i
    .port_state_in_8_0_1   (shiftRows_port_state_out_8_0_1[2:0]  ), //i
    .port_state_in_8_0_2   (shiftRows_port_state_out_8_0_2[2:0]  ), //i
    .port_state_in_8_0_3   (shiftRows_port_state_out_8_0_3[2:0]  ), //i
    .port_state_in_8_0_4   (shiftRows_port_state_out_8_0_4[2:0]  ), //i
    .port_state_in_8_0_5   (shiftRows_port_state_out_8_0_5[2:0]  ), //i
    .port_state_in_8_0_6   (shiftRows_port_state_out_8_0_6[2:0]  ), //i
    .port_state_in_8_0_7   (shiftRows_port_state_out_8_0_7[2:0]  ), //i
    .port_state_in_8_1_0   (shiftRows_port_state_out_8_1_0[2:0]  ), //i
    .port_state_in_8_1_1   (shiftRows_port_state_out_8_1_1[2:0]  ), //i
    .port_state_in_8_1_2   (shiftRows_port_state_out_8_1_2[2:0]  ), //i
    .port_state_in_8_1_3   (shiftRows_port_state_out_8_1_3[2:0]  ), //i
    .port_state_in_8_1_4   (shiftRows_port_state_out_8_1_4[2:0]  ), //i
    .port_state_in_8_1_5   (shiftRows_port_state_out_8_1_5[2:0]  ), //i
    .port_state_in_8_1_6   (shiftRows_port_state_out_8_1_6[2:0]  ), //i
    .port_state_in_8_1_7   (shiftRows_port_state_out_8_1_7[2:0]  ), //i
    .port_state_in_8_2_0   (shiftRows_port_state_out_8_2_0[2:0]  ), //i
    .port_state_in_8_2_1   (shiftRows_port_state_out_8_2_1[2:0]  ), //i
    .port_state_in_8_2_2   (shiftRows_port_state_out_8_2_2[2:0]  ), //i
    .port_state_in_8_2_3   (shiftRows_port_state_out_8_2_3[2:0]  ), //i
    .port_state_in_8_2_4   (shiftRows_port_state_out_8_2_4[2:0]  ), //i
    .port_state_in_8_2_5   (shiftRows_port_state_out_8_2_5[2:0]  ), //i
    .port_state_in_8_2_6   (shiftRows_port_state_out_8_2_6[2:0]  ), //i
    .port_state_in_8_2_7   (shiftRows_port_state_out_8_2_7[2:0]  ), //i
    .port_state_in_8_3_0   (shiftRows_port_state_out_8_3_0[2:0]  ), //i
    .port_state_in_8_3_1   (shiftRows_port_state_out_8_3_1[2:0]  ), //i
    .port_state_in_8_3_2   (shiftRows_port_state_out_8_3_2[2:0]  ), //i
    .port_state_in_8_3_3   (shiftRows_port_state_out_8_3_3[2:0]  ), //i
    .port_state_in_8_3_4   (shiftRows_port_state_out_8_3_4[2:0]  ), //i
    .port_state_in_8_3_5   (shiftRows_port_state_out_8_3_5[2:0]  ), //i
    .port_state_in_8_3_6   (shiftRows_port_state_out_8_3_6[2:0]  ), //i
    .port_state_in_8_3_7   (shiftRows_port_state_out_8_3_7[2:0]  ), //i
    .port_state_in_9_0_0   (shiftRows_port_state_out_9_0_0[2:0]  ), //i
    .port_state_in_9_0_1   (shiftRows_port_state_out_9_0_1[2:0]  ), //i
    .port_state_in_9_0_2   (shiftRows_port_state_out_9_0_2[2:0]  ), //i
    .port_state_in_9_0_3   (shiftRows_port_state_out_9_0_3[2:0]  ), //i
    .port_state_in_9_0_4   (shiftRows_port_state_out_9_0_4[2:0]  ), //i
    .port_state_in_9_0_5   (shiftRows_port_state_out_9_0_5[2:0]  ), //i
    .port_state_in_9_0_6   (shiftRows_port_state_out_9_0_6[2:0]  ), //i
    .port_state_in_9_0_7   (shiftRows_port_state_out_9_0_7[2:0]  ), //i
    .port_state_in_9_1_0   (shiftRows_port_state_out_9_1_0[2:0]  ), //i
    .port_state_in_9_1_1   (shiftRows_port_state_out_9_1_1[2:0]  ), //i
    .port_state_in_9_1_2   (shiftRows_port_state_out_9_1_2[2:0]  ), //i
    .port_state_in_9_1_3   (shiftRows_port_state_out_9_1_3[2:0]  ), //i
    .port_state_in_9_1_4   (shiftRows_port_state_out_9_1_4[2:0]  ), //i
    .port_state_in_9_1_5   (shiftRows_port_state_out_9_1_5[2:0]  ), //i
    .port_state_in_9_1_6   (shiftRows_port_state_out_9_1_6[2:0]  ), //i
    .port_state_in_9_1_7   (shiftRows_port_state_out_9_1_7[2:0]  ), //i
    .port_state_in_9_2_0   (shiftRows_port_state_out_9_2_0[2:0]  ), //i
    .port_state_in_9_2_1   (shiftRows_port_state_out_9_2_1[2:0]  ), //i
    .port_state_in_9_2_2   (shiftRows_port_state_out_9_2_2[2:0]  ), //i
    .port_state_in_9_2_3   (shiftRows_port_state_out_9_2_3[2:0]  ), //i
    .port_state_in_9_2_4   (shiftRows_port_state_out_9_2_4[2:0]  ), //i
    .port_state_in_9_2_5   (shiftRows_port_state_out_9_2_5[2:0]  ), //i
    .port_state_in_9_2_6   (shiftRows_port_state_out_9_2_6[2:0]  ), //i
    .port_state_in_9_2_7   (shiftRows_port_state_out_9_2_7[2:0]  ), //i
    .port_state_in_9_3_0   (shiftRows_port_state_out_9_3_0[2:0]  ), //i
    .port_state_in_9_3_1   (shiftRows_port_state_out_9_3_1[2:0]  ), //i
    .port_state_in_9_3_2   (shiftRows_port_state_out_9_3_2[2:0]  ), //i
    .port_state_in_9_3_3   (shiftRows_port_state_out_9_3_3[2:0]  ), //i
    .port_state_in_9_3_4   (shiftRows_port_state_out_9_3_4[2:0]  ), //i
    .port_state_in_9_3_5   (shiftRows_port_state_out_9_3_5[2:0]  ), //i
    .port_state_in_9_3_6   (shiftRows_port_state_out_9_3_6[2:0]  ), //i
    .port_state_in_9_3_7   (shiftRows_port_state_out_9_3_7[2:0]  ), //i
    .port_state_in_10_0_0  (shiftRows_port_state_out_10_0_0[2:0] ), //i
    .port_state_in_10_0_1  (shiftRows_port_state_out_10_0_1[2:0] ), //i
    .port_state_in_10_0_2  (shiftRows_port_state_out_10_0_2[2:0] ), //i
    .port_state_in_10_0_3  (shiftRows_port_state_out_10_0_3[2:0] ), //i
    .port_state_in_10_0_4  (shiftRows_port_state_out_10_0_4[2:0] ), //i
    .port_state_in_10_0_5  (shiftRows_port_state_out_10_0_5[2:0] ), //i
    .port_state_in_10_0_6  (shiftRows_port_state_out_10_0_6[2:0] ), //i
    .port_state_in_10_0_7  (shiftRows_port_state_out_10_0_7[2:0] ), //i
    .port_state_in_10_1_0  (shiftRows_port_state_out_10_1_0[2:0] ), //i
    .port_state_in_10_1_1  (shiftRows_port_state_out_10_1_1[2:0] ), //i
    .port_state_in_10_1_2  (shiftRows_port_state_out_10_1_2[2:0] ), //i
    .port_state_in_10_1_3  (shiftRows_port_state_out_10_1_3[2:0] ), //i
    .port_state_in_10_1_4  (shiftRows_port_state_out_10_1_4[2:0] ), //i
    .port_state_in_10_1_5  (shiftRows_port_state_out_10_1_5[2:0] ), //i
    .port_state_in_10_1_6  (shiftRows_port_state_out_10_1_6[2:0] ), //i
    .port_state_in_10_1_7  (shiftRows_port_state_out_10_1_7[2:0] ), //i
    .port_state_in_10_2_0  (shiftRows_port_state_out_10_2_0[2:0] ), //i
    .port_state_in_10_2_1  (shiftRows_port_state_out_10_2_1[2:0] ), //i
    .port_state_in_10_2_2  (shiftRows_port_state_out_10_2_2[2:0] ), //i
    .port_state_in_10_2_3  (shiftRows_port_state_out_10_2_3[2:0] ), //i
    .port_state_in_10_2_4  (shiftRows_port_state_out_10_2_4[2:0] ), //i
    .port_state_in_10_2_5  (shiftRows_port_state_out_10_2_5[2:0] ), //i
    .port_state_in_10_2_6  (shiftRows_port_state_out_10_2_6[2:0] ), //i
    .port_state_in_10_2_7  (shiftRows_port_state_out_10_2_7[2:0] ), //i
    .port_state_in_10_3_0  (shiftRows_port_state_out_10_3_0[2:0] ), //i
    .port_state_in_10_3_1  (shiftRows_port_state_out_10_3_1[2:0] ), //i
    .port_state_in_10_3_2  (shiftRows_port_state_out_10_3_2[2:0] ), //i
    .port_state_in_10_3_3  (shiftRows_port_state_out_10_3_3[2:0] ), //i
    .port_state_in_10_3_4  (shiftRows_port_state_out_10_3_4[2:0] ), //i
    .port_state_in_10_3_5  (shiftRows_port_state_out_10_3_5[2:0] ), //i
    .port_state_in_10_3_6  (shiftRows_port_state_out_10_3_6[2:0] ), //i
    .port_state_in_10_3_7  (shiftRows_port_state_out_10_3_7[2:0] ), //i
    .port_state_in_11_0_0  (shiftRows_port_state_out_11_0_0[2:0] ), //i
    .port_state_in_11_0_1  (shiftRows_port_state_out_11_0_1[2:0] ), //i
    .port_state_in_11_0_2  (shiftRows_port_state_out_11_0_2[2:0] ), //i
    .port_state_in_11_0_3  (shiftRows_port_state_out_11_0_3[2:0] ), //i
    .port_state_in_11_0_4  (shiftRows_port_state_out_11_0_4[2:0] ), //i
    .port_state_in_11_0_5  (shiftRows_port_state_out_11_0_5[2:0] ), //i
    .port_state_in_11_0_6  (shiftRows_port_state_out_11_0_6[2:0] ), //i
    .port_state_in_11_0_7  (shiftRows_port_state_out_11_0_7[2:0] ), //i
    .port_state_in_11_1_0  (shiftRows_port_state_out_11_1_0[2:0] ), //i
    .port_state_in_11_1_1  (shiftRows_port_state_out_11_1_1[2:0] ), //i
    .port_state_in_11_1_2  (shiftRows_port_state_out_11_1_2[2:0] ), //i
    .port_state_in_11_1_3  (shiftRows_port_state_out_11_1_3[2:0] ), //i
    .port_state_in_11_1_4  (shiftRows_port_state_out_11_1_4[2:0] ), //i
    .port_state_in_11_1_5  (shiftRows_port_state_out_11_1_5[2:0] ), //i
    .port_state_in_11_1_6  (shiftRows_port_state_out_11_1_6[2:0] ), //i
    .port_state_in_11_1_7  (shiftRows_port_state_out_11_1_7[2:0] ), //i
    .port_state_in_11_2_0  (shiftRows_port_state_out_11_2_0[2:0] ), //i
    .port_state_in_11_2_1  (shiftRows_port_state_out_11_2_1[2:0] ), //i
    .port_state_in_11_2_2  (shiftRows_port_state_out_11_2_2[2:0] ), //i
    .port_state_in_11_2_3  (shiftRows_port_state_out_11_2_3[2:0] ), //i
    .port_state_in_11_2_4  (shiftRows_port_state_out_11_2_4[2:0] ), //i
    .port_state_in_11_2_5  (shiftRows_port_state_out_11_2_5[2:0] ), //i
    .port_state_in_11_2_6  (shiftRows_port_state_out_11_2_6[2:0] ), //i
    .port_state_in_11_2_7  (shiftRows_port_state_out_11_2_7[2:0] ), //i
    .port_state_in_11_3_0  (shiftRows_port_state_out_11_3_0[2:0] ), //i
    .port_state_in_11_3_1  (shiftRows_port_state_out_11_3_1[2:0] ), //i
    .port_state_in_11_3_2  (shiftRows_port_state_out_11_3_2[2:0] ), //i
    .port_state_in_11_3_3  (shiftRows_port_state_out_11_3_3[2:0] ), //i
    .port_state_in_11_3_4  (shiftRows_port_state_out_11_3_4[2:0] ), //i
    .port_state_in_11_3_5  (shiftRows_port_state_out_11_3_5[2:0] ), //i
    .port_state_in_11_3_6  (shiftRows_port_state_out_11_3_6[2:0] ), //i
    .port_state_in_11_3_7  (shiftRows_port_state_out_11_3_7[2:0] ), //i
    .port_state_in_12_0_0  (shiftRows_port_state_out_12_0_0[2:0] ), //i
    .port_state_in_12_0_1  (shiftRows_port_state_out_12_0_1[2:0] ), //i
    .port_state_in_12_0_2  (shiftRows_port_state_out_12_0_2[2:0] ), //i
    .port_state_in_12_0_3  (shiftRows_port_state_out_12_0_3[2:0] ), //i
    .port_state_in_12_0_4  (shiftRows_port_state_out_12_0_4[2:0] ), //i
    .port_state_in_12_0_5  (shiftRows_port_state_out_12_0_5[2:0] ), //i
    .port_state_in_12_0_6  (shiftRows_port_state_out_12_0_6[2:0] ), //i
    .port_state_in_12_0_7  (shiftRows_port_state_out_12_0_7[2:0] ), //i
    .port_state_in_12_1_0  (shiftRows_port_state_out_12_1_0[2:0] ), //i
    .port_state_in_12_1_1  (shiftRows_port_state_out_12_1_1[2:0] ), //i
    .port_state_in_12_1_2  (shiftRows_port_state_out_12_1_2[2:0] ), //i
    .port_state_in_12_1_3  (shiftRows_port_state_out_12_1_3[2:0] ), //i
    .port_state_in_12_1_4  (shiftRows_port_state_out_12_1_4[2:0] ), //i
    .port_state_in_12_1_5  (shiftRows_port_state_out_12_1_5[2:0] ), //i
    .port_state_in_12_1_6  (shiftRows_port_state_out_12_1_6[2:0] ), //i
    .port_state_in_12_1_7  (shiftRows_port_state_out_12_1_7[2:0] ), //i
    .port_state_in_12_2_0  (shiftRows_port_state_out_12_2_0[2:0] ), //i
    .port_state_in_12_2_1  (shiftRows_port_state_out_12_2_1[2:0] ), //i
    .port_state_in_12_2_2  (shiftRows_port_state_out_12_2_2[2:0] ), //i
    .port_state_in_12_2_3  (shiftRows_port_state_out_12_2_3[2:0] ), //i
    .port_state_in_12_2_4  (shiftRows_port_state_out_12_2_4[2:0] ), //i
    .port_state_in_12_2_5  (shiftRows_port_state_out_12_2_5[2:0] ), //i
    .port_state_in_12_2_6  (shiftRows_port_state_out_12_2_6[2:0] ), //i
    .port_state_in_12_2_7  (shiftRows_port_state_out_12_2_7[2:0] ), //i
    .port_state_in_12_3_0  (shiftRows_port_state_out_12_3_0[2:0] ), //i
    .port_state_in_12_3_1  (shiftRows_port_state_out_12_3_1[2:0] ), //i
    .port_state_in_12_3_2  (shiftRows_port_state_out_12_3_2[2:0] ), //i
    .port_state_in_12_3_3  (shiftRows_port_state_out_12_3_3[2:0] ), //i
    .port_state_in_12_3_4  (shiftRows_port_state_out_12_3_4[2:0] ), //i
    .port_state_in_12_3_5  (shiftRows_port_state_out_12_3_5[2:0] ), //i
    .port_state_in_12_3_6  (shiftRows_port_state_out_12_3_6[2:0] ), //i
    .port_state_in_12_3_7  (shiftRows_port_state_out_12_3_7[2:0] ), //i
    .port_state_in_13_0_0  (shiftRows_port_state_out_13_0_0[2:0] ), //i
    .port_state_in_13_0_1  (shiftRows_port_state_out_13_0_1[2:0] ), //i
    .port_state_in_13_0_2  (shiftRows_port_state_out_13_0_2[2:0] ), //i
    .port_state_in_13_0_3  (shiftRows_port_state_out_13_0_3[2:0] ), //i
    .port_state_in_13_0_4  (shiftRows_port_state_out_13_0_4[2:0] ), //i
    .port_state_in_13_0_5  (shiftRows_port_state_out_13_0_5[2:0] ), //i
    .port_state_in_13_0_6  (shiftRows_port_state_out_13_0_6[2:0] ), //i
    .port_state_in_13_0_7  (shiftRows_port_state_out_13_0_7[2:0] ), //i
    .port_state_in_13_1_0  (shiftRows_port_state_out_13_1_0[2:0] ), //i
    .port_state_in_13_1_1  (shiftRows_port_state_out_13_1_1[2:0] ), //i
    .port_state_in_13_1_2  (shiftRows_port_state_out_13_1_2[2:0] ), //i
    .port_state_in_13_1_3  (shiftRows_port_state_out_13_1_3[2:0] ), //i
    .port_state_in_13_1_4  (shiftRows_port_state_out_13_1_4[2:0] ), //i
    .port_state_in_13_1_5  (shiftRows_port_state_out_13_1_5[2:0] ), //i
    .port_state_in_13_1_6  (shiftRows_port_state_out_13_1_6[2:0] ), //i
    .port_state_in_13_1_7  (shiftRows_port_state_out_13_1_7[2:0] ), //i
    .port_state_in_13_2_0  (shiftRows_port_state_out_13_2_0[2:0] ), //i
    .port_state_in_13_2_1  (shiftRows_port_state_out_13_2_1[2:0] ), //i
    .port_state_in_13_2_2  (shiftRows_port_state_out_13_2_2[2:0] ), //i
    .port_state_in_13_2_3  (shiftRows_port_state_out_13_2_3[2:0] ), //i
    .port_state_in_13_2_4  (shiftRows_port_state_out_13_2_4[2:0] ), //i
    .port_state_in_13_2_5  (shiftRows_port_state_out_13_2_5[2:0] ), //i
    .port_state_in_13_2_6  (shiftRows_port_state_out_13_2_6[2:0] ), //i
    .port_state_in_13_2_7  (shiftRows_port_state_out_13_2_7[2:0] ), //i
    .port_state_in_13_3_0  (shiftRows_port_state_out_13_3_0[2:0] ), //i
    .port_state_in_13_3_1  (shiftRows_port_state_out_13_3_1[2:0] ), //i
    .port_state_in_13_3_2  (shiftRows_port_state_out_13_3_2[2:0] ), //i
    .port_state_in_13_3_3  (shiftRows_port_state_out_13_3_3[2:0] ), //i
    .port_state_in_13_3_4  (shiftRows_port_state_out_13_3_4[2:0] ), //i
    .port_state_in_13_3_5  (shiftRows_port_state_out_13_3_5[2:0] ), //i
    .port_state_in_13_3_6  (shiftRows_port_state_out_13_3_6[2:0] ), //i
    .port_state_in_13_3_7  (shiftRows_port_state_out_13_3_7[2:0] ), //i
    .port_state_in_14_0_0  (shiftRows_port_state_out_14_0_0[2:0] ), //i
    .port_state_in_14_0_1  (shiftRows_port_state_out_14_0_1[2:0] ), //i
    .port_state_in_14_0_2  (shiftRows_port_state_out_14_0_2[2:0] ), //i
    .port_state_in_14_0_3  (shiftRows_port_state_out_14_0_3[2:0] ), //i
    .port_state_in_14_0_4  (shiftRows_port_state_out_14_0_4[2:0] ), //i
    .port_state_in_14_0_5  (shiftRows_port_state_out_14_0_5[2:0] ), //i
    .port_state_in_14_0_6  (shiftRows_port_state_out_14_0_6[2:0] ), //i
    .port_state_in_14_0_7  (shiftRows_port_state_out_14_0_7[2:0] ), //i
    .port_state_in_14_1_0  (shiftRows_port_state_out_14_1_0[2:0] ), //i
    .port_state_in_14_1_1  (shiftRows_port_state_out_14_1_1[2:0] ), //i
    .port_state_in_14_1_2  (shiftRows_port_state_out_14_1_2[2:0] ), //i
    .port_state_in_14_1_3  (shiftRows_port_state_out_14_1_3[2:0] ), //i
    .port_state_in_14_1_4  (shiftRows_port_state_out_14_1_4[2:0] ), //i
    .port_state_in_14_1_5  (shiftRows_port_state_out_14_1_5[2:0] ), //i
    .port_state_in_14_1_6  (shiftRows_port_state_out_14_1_6[2:0] ), //i
    .port_state_in_14_1_7  (shiftRows_port_state_out_14_1_7[2:0] ), //i
    .port_state_in_14_2_0  (shiftRows_port_state_out_14_2_0[2:0] ), //i
    .port_state_in_14_2_1  (shiftRows_port_state_out_14_2_1[2:0] ), //i
    .port_state_in_14_2_2  (shiftRows_port_state_out_14_2_2[2:0] ), //i
    .port_state_in_14_2_3  (shiftRows_port_state_out_14_2_3[2:0] ), //i
    .port_state_in_14_2_4  (shiftRows_port_state_out_14_2_4[2:0] ), //i
    .port_state_in_14_2_5  (shiftRows_port_state_out_14_2_5[2:0] ), //i
    .port_state_in_14_2_6  (shiftRows_port_state_out_14_2_6[2:0] ), //i
    .port_state_in_14_2_7  (shiftRows_port_state_out_14_2_7[2:0] ), //i
    .port_state_in_14_3_0  (shiftRows_port_state_out_14_3_0[2:0] ), //i
    .port_state_in_14_3_1  (shiftRows_port_state_out_14_3_1[2:0] ), //i
    .port_state_in_14_3_2  (shiftRows_port_state_out_14_3_2[2:0] ), //i
    .port_state_in_14_3_3  (shiftRows_port_state_out_14_3_3[2:0] ), //i
    .port_state_in_14_3_4  (shiftRows_port_state_out_14_3_4[2:0] ), //i
    .port_state_in_14_3_5  (shiftRows_port_state_out_14_3_5[2:0] ), //i
    .port_state_in_14_3_6  (shiftRows_port_state_out_14_3_6[2:0] ), //i
    .port_state_in_14_3_7  (shiftRows_port_state_out_14_3_7[2:0] ), //i
    .port_state_in_15_0_0  (shiftRows_port_state_out_15_0_0[2:0] ), //i
    .port_state_in_15_0_1  (shiftRows_port_state_out_15_0_1[2:0] ), //i
    .port_state_in_15_0_2  (shiftRows_port_state_out_15_0_2[2:0] ), //i
    .port_state_in_15_0_3  (shiftRows_port_state_out_15_0_3[2:0] ), //i
    .port_state_in_15_0_4  (shiftRows_port_state_out_15_0_4[2:0] ), //i
    .port_state_in_15_0_5  (shiftRows_port_state_out_15_0_5[2:0] ), //i
    .port_state_in_15_0_6  (shiftRows_port_state_out_15_0_6[2:0] ), //i
    .port_state_in_15_0_7  (shiftRows_port_state_out_15_0_7[2:0] ), //i
    .port_state_in_15_1_0  (shiftRows_port_state_out_15_1_0[2:0] ), //i
    .port_state_in_15_1_1  (shiftRows_port_state_out_15_1_1[2:0] ), //i
    .port_state_in_15_1_2  (shiftRows_port_state_out_15_1_2[2:0] ), //i
    .port_state_in_15_1_3  (shiftRows_port_state_out_15_1_3[2:0] ), //i
    .port_state_in_15_1_4  (shiftRows_port_state_out_15_1_4[2:0] ), //i
    .port_state_in_15_1_5  (shiftRows_port_state_out_15_1_5[2:0] ), //i
    .port_state_in_15_1_6  (shiftRows_port_state_out_15_1_6[2:0] ), //i
    .port_state_in_15_1_7  (shiftRows_port_state_out_15_1_7[2:0] ), //i
    .port_state_in_15_2_0  (shiftRows_port_state_out_15_2_0[2:0] ), //i
    .port_state_in_15_2_1  (shiftRows_port_state_out_15_2_1[2:0] ), //i
    .port_state_in_15_2_2  (shiftRows_port_state_out_15_2_2[2:0] ), //i
    .port_state_in_15_2_3  (shiftRows_port_state_out_15_2_3[2:0] ), //i
    .port_state_in_15_2_4  (shiftRows_port_state_out_15_2_4[2:0] ), //i
    .port_state_in_15_2_5  (shiftRows_port_state_out_15_2_5[2:0] ), //i
    .port_state_in_15_2_6  (shiftRows_port_state_out_15_2_6[2:0] ), //i
    .port_state_in_15_2_7  (shiftRows_port_state_out_15_2_7[2:0] ), //i
    .port_state_in_15_3_0  (shiftRows_port_state_out_15_3_0[2:0] ), //i
    .port_state_in_15_3_1  (shiftRows_port_state_out_15_3_1[2:0] ), //i
    .port_state_in_15_3_2  (shiftRows_port_state_out_15_3_2[2:0] ), //i
    .port_state_in_15_3_3  (shiftRows_port_state_out_15_3_3[2:0] ), //i
    .port_state_in_15_3_4  (shiftRows_port_state_out_15_3_4[2:0] ), //i
    .port_state_in_15_3_5  (shiftRows_port_state_out_15_3_5[2:0] ), //i
    .port_state_in_15_3_6  (shiftRows_port_state_out_15_3_6[2:0] ), //i
    .port_state_in_15_3_7  (shiftRows_port_state_out_15_3_7[2:0] ), //i
    .port_state_out_0_0_0  (mixColumns_port_state_out_0_0_0[2:0] ), //o
    .port_state_out_0_0_1  (mixColumns_port_state_out_0_0_1[2:0] ), //o
    .port_state_out_0_0_2  (mixColumns_port_state_out_0_0_2[2:0] ), //o
    .port_state_out_0_0_3  (mixColumns_port_state_out_0_0_3[2:0] ), //o
    .port_state_out_0_0_4  (mixColumns_port_state_out_0_0_4[2:0] ), //o
    .port_state_out_0_0_5  (mixColumns_port_state_out_0_0_5[2:0] ), //o
    .port_state_out_0_0_6  (mixColumns_port_state_out_0_0_6[2:0] ), //o
    .port_state_out_0_0_7  (mixColumns_port_state_out_0_0_7[2:0] ), //o
    .port_state_out_0_1_0  (mixColumns_port_state_out_0_1_0[2:0] ), //o
    .port_state_out_0_1_1  (mixColumns_port_state_out_0_1_1[2:0] ), //o
    .port_state_out_0_1_2  (mixColumns_port_state_out_0_1_2[2:0] ), //o
    .port_state_out_0_1_3  (mixColumns_port_state_out_0_1_3[2:0] ), //o
    .port_state_out_0_1_4  (mixColumns_port_state_out_0_1_4[2:0] ), //o
    .port_state_out_0_1_5  (mixColumns_port_state_out_0_1_5[2:0] ), //o
    .port_state_out_0_1_6  (mixColumns_port_state_out_0_1_6[2:0] ), //o
    .port_state_out_0_1_7  (mixColumns_port_state_out_0_1_7[2:0] ), //o
    .port_state_out_0_2_0  (mixColumns_port_state_out_0_2_0[2:0] ), //o
    .port_state_out_0_2_1  (mixColumns_port_state_out_0_2_1[2:0] ), //o
    .port_state_out_0_2_2  (mixColumns_port_state_out_0_2_2[2:0] ), //o
    .port_state_out_0_2_3  (mixColumns_port_state_out_0_2_3[2:0] ), //o
    .port_state_out_0_2_4  (mixColumns_port_state_out_0_2_4[2:0] ), //o
    .port_state_out_0_2_5  (mixColumns_port_state_out_0_2_5[2:0] ), //o
    .port_state_out_0_2_6  (mixColumns_port_state_out_0_2_6[2:0] ), //o
    .port_state_out_0_2_7  (mixColumns_port_state_out_0_2_7[2:0] ), //o
    .port_state_out_0_3_0  (mixColumns_port_state_out_0_3_0[2:0] ), //o
    .port_state_out_0_3_1  (mixColumns_port_state_out_0_3_1[2:0] ), //o
    .port_state_out_0_3_2  (mixColumns_port_state_out_0_3_2[2:0] ), //o
    .port_state_out_0_3_3  (mixColumns_port_state_out_0_3_3[2:0] ), //o
    .port_state_out_0_3_4  (mixColumns_port_state_out_0_3_4[2:0] ), //o
    .port_state_out_0_3_5  (mixColumns_port_state_out_0_3_5[2:0] ), //o
    .port_state_out_0_3_6  (mixColumns_port_state_out_0_3_6[2:0] ), //o
    .port_state_out_0_3_7  (mixColumns_port_state_out_0_3_7[2:0] ), //o
    .port_state_out_1_0_0  (mixColumns_port_state_out_1_0_0[2:0] ), //o
    .port_state_out_1_0_1  (mixColumns_port_state_out_1_0_1[2:0] ), //o
    .port_state_out_1_0_2  (mixColumns_port_state_out_1_0_2[2:0] ), //o
    .port_state_out_1_0_3  (mixColumns_port_state_out_1_0_3[2:0] ), //o
    .port_state_out_1_0_4  (mixColumns_port_state_out_1_0_4[2:0] ), //o
    .port_state_out_1_0_5  (mixColumns_port_state_out_1_0_5[2:0] ), //o
    .port_state_out_1_0_6  (mixColumns_port_state_out_1_0_6[2:0] ), //o
    .port_state_out_1_0_7  (mixColumns_port_state_out_1_0_7[2:0] ), //o
    .port_state_out_1_1_0  (mixColumns_port_state_out_1_1_0[2:0] ), //o
    .port_state_out_1_1_1  (mixColumns_port_state_out_1_1_1[2:0] ), //o
    .port_state_out_1_1_2  (mixColumns_port_state_out_1_1_2[2:0] ), //o
    .port_state_out_1_1_3  (mixColumns_port_state_out_1_1_3[2:0] ), //o
    .port_state_out_1_1_4  (mixColumns_port_state_out_1_1_4[2:0] ), //o
    .port_state_out_1_1_5  (mixColumns_port_state_out_1_1_5[2:0] ), //o
    .port_state_out_1_1_6  (mixColumns_port_state_out_1_1_6[2:0] ), //o
    .port_state_out_1_1_7  (mixColumns_port_state_out_1_1_7[2:0] ), //o
    .port_state_out_1_2_0  (mixColumns_port_state_out_1_2_0[2:0] ), //o
    .port_state_out_1_2_1  (mixColumns_port_state_out_1_2_1[2:0] ), //o
    .port_state_out_1_2_2  (mixColumns_port_state_out_1_2_2[2:0] ), //o
    .port_state_out_1_2_3  (mixColumns_port_state_out_1_2_3[2:0] ), //o
    .port_state_out_1_2_4  (mixColumns_port_state_out_1_2_4[2:0] ), //o
    .port_state_out_1_2_5  (mixColumns_port_state_out_1_2_5[2:0] ), //o
    .port_state_out_1_2_6  (mixColumns_port_state_out_1_2_6[2:0] ), //o
    .port_state_out_1_2_7  (mixColumns_port_state_out_1_2_7[2:0] ), //o
    .port_state_out_1_3_0  (mixColumns_port_state_out_1_3_0[2:0] ), //o
    .port_state_out_1_3_1  (mixColumns_port_state_out_1_3_1[2:0] ), //o
    .port_state_out_1_3_2  (mixColumns_port_state_out_1_3_2[2:0] ), //o
    .port_state_out_1_3_3  (mixColumns_port_state_out_1_3_3[2:0] ), //o
    .port_state_out_1_3_4  (mixColumns_port_state_out_1_3_4[2:0] ), //o
    .port_state_out_1_3_5  (mixColumns_port_state_out_1_3_5[2:0] ), //o
    .port_state_out_1_3_6  (mixColumns_port_state_out_1_3_6[2:0] ), //o
    .port_state_out_1_3_7  (mixColumns_port_state_out_1_3_7[2:0] ), //o
    .port_state_out_2_0_0  (mixColumns_port_state_out_2_0_0[2:0] ), //o
    .port_state_out_2_0_1  (mixColumns_port_state_out_2_0_1[2:0] ), //o
    .port_state_out_2_0_2  (mixColumns_port_state_out_2_0_2[2:0] ), //o
    .port_state_out_2_0_3  (mixColumns_port_state_out_2_0_3[2:0] ), //o
    .port_state_out_2_0_4  (mixColumns_port_state_out_2_0_4[2:0] ), //o
    .port_state_out_2_0_5  (mixColumns_port_state_out_2_0_5[2:0] ), //o
    .port_state_out_2_0_6  (mixColumns_port_state_out_2_0_6[2:0] ), //o
    .port_state_out_2_0_7  (mixColumns_port_state_out_2_0_7[2:0] ), //o
    .port_state_out_2_1_0  (mixColumns_port_state_out_2_1_0[2:0] ), //o
    .port_state_out_2_1_1  (mixColumns_port_state_out_2_1_1[2:0] ), //o
    .port_state_out_2_1_2  (mixColumns_port_state_out_2_1_2[2:0] ), //o
    .port_state_out_2_1_3  (mixColumns_port_state_out_2_1_3[2:0] ), //o
    .port_state_out_2_1_4  (mixColumns_port_state_out_2_1_4[2:0] ), //o
    .port_state_out_2_1_5  (mixColumns_port_state_out_2_1_5[2:0] ), //o
    .port_state_out_2_1_6  (mixColumns_port_state_out_2_1_6[2:0] ), //o
    .port_state_out_2_1_7  (mixColumns_port_state_out_2_1_7[2:0] ), //o
    .port_state_out_2_2_0  (mixColumns_port_state_out_2_2_0[2:0] ), //o
    .port_state_out_2_2_1  (mixColumns_port_state_out_2_2_1[2:0] ), //o
    .port_state_out_2_2_2  (mixColumns_port_state_out_2_2_2[2:0] ), //o
    .port_state_out_2_2_3  (mixColumns_port_state_out_2_2_3[2:0] ), //o
    .port_state_out_2_2_4  (mixColumns_port_state_out_2_2_4[2:0] ), //o
    .port_state_out_2_2_5  (mixColumns_port_state_out_2_2_5[2:0] ), //o
    .port_state_out_2_2_6  (mixColumns_port_state_out_2_2_6[2:0] ), //o
    .port_state_out_2_2_7  (mixColumns_port_state_out_2_2_7[2:0] ), //o
    .port_state_out_2_3_0  (mixColumns_port_state_out_2_3_0[2:0] ), //o
    .port_state_out_2_3_1  (mixColumns_port_state_out_2_3_1[2:0] ), //o
    .port_state_out_2_3_2  (mixColumns_port_state_out_2_3_2[2:0] ), //o
    .port_state_out_2_3_3  (mixColumns_port_state_out_2_3_3[2:0] ), //o
    .port_state_out_2_3_4  (mixColumns_port_state_out_2_3_4[2:0] ), //o
    .port_state_out_2_3_5  (mixColumns_port_state_out_2_3_5[2:0] ), //o
    .port_state_out_2_3_6  (mixColumns_port_state_out_2_3_6[2:0] ), //o
    .port_state_out_2_3_7  (mixColumns_port_state_out_2_3_7[2:0] ), //o
    .port_state_out_3_0_0  (mixColumns_port_state_out_3_0_0[2:0] ), //o
    .port_state_out_3_0_1  (mixColumns_port_state_out_3_0_1[2:0] ), //o
    .port_state_out_3_0_2  (mixColumns_port_state_out_3_0_2[2:0] ), //o
    .port_state_out_3_0_3  (mixColumns_port_state_out_3_0_3[2:0] ), //o
    .port_state_out_3_0_4  (mixColumns_port_state_out_3_0_4[2:0] ), //o
    .port_state_out_3_0_5  (mixColumns_port_state_out_3_0_5[2:0] ), //o
    .port_state_out_3_0_6  (mixColumns_port_state_out_3_0_6[2:0] ), //o
    .port_state_out_3_0_7  (mixColumns_port_state_out_3_0_7[2:0] ), //o
    .port_state_out_3_1_0  (mixColumns_port_state_out_3_1_0[2:0] ), //o
    .port_state_out_3_1_1  (mixColumns_port_state_out_3_1_1[2:0] ), //o
    .port_state_out_3_1_2  (mixColumns_port_state_out_3_1_2[2:0] ), //o
    .port_state_out_3_1_3  (mixColumns_port_state_out_3_1_3[2:0] ), //o
    .port_state_out_3_1_4  (mixColumns_port_state_out_3_1_4[2:0] ), //o
    .port_state_out_3_1_5  (mixColumns_port_state_out_3_1_5[2:0] ), //o
    .port_state_out_3_1_6  (mixColumns_port_state_out_3_1_6[2:0] ), //o
    .port_state_out_3_1_7  (mixColumns_port_state_out_3_1_7[2:0] ), //o
    .port_state_out_3_2_0  (mixColumns_port_state_out_3_2_0[2:0] ), //o
    .port_state_out_3_2_1  (mixColumns_port_state_out_3_2_1[2:0] ), //o
    .port_state_out_3_2_2  (mixColumns_port_state_out_3_2_2[2:0] ), //o
    .port_state_out_3_2_3  (mixColumns_port_state_out_3_2_3[2:0] ), //o
    .port_state_out_3_2_4  (mixColumns_port_state_out_3_2_4[2:0] ), //o
    .port_state_out_3_2_5  (mixColumns_port_state_out_3_2_5[2:0] ), //o
    .port_state_out_3_2_6  (mixColumns_port_state_out_3_2_6[2:0] ), //o
    .port_state_out_3_2_7  (mixColumns_port_state_out_3_2_7[2:0] ), //o
    .port_state_out_3_3_0  (mixColumns_port_state_out_3_3_0[2:0] ), //o
    .port_state_out_3_3_1  (mixColumns_port_state_out_3_3_1[2:0] ), //o
    .port_state_out_3_3_2  (mixColumns_port_state_out_3_3_2[2:0] ), //o
    .port_state_out_3_3_3  (mixColumns_port_state_out_3_3_3[2:0] ), //o
    .port_state_out_3_3_4  (mixColumns_port_state_out_3_3_4[2:0] ), //o
    .port_state_out_3_3_5  (mixColumns_port_state_out_3_3_5[2:0] ), //o
    .port_state_out_3_3_6  (mixColumns_port_state_out_3_3_6[2:0] ), //o
    .port_state_out_3_3_7  (mixColumns_port_state_out_3_3_7[2:0] ), //o
    .port_state_out_4_0_0  (mixColumns_port_state_out_4_0_0[2:0] ), //o
    .port_state_out_4_0_1  (mixColumns_port_state_out_4_0_1[2:0] ), //o
    .port_state_out_4_0_2  (mixColumns_port_state_out_4_0_2[2:0] ), //o
    .port_state_out_4_0_3  (mixColumns_port_state_out_4_0_3[2:0] ), //o
    .port_state_out_4_0_4  (mixColumns_port_state_out_4_0_4[2:0] ), //o
    .port_state_out_4_0_5  (mixColumns_port_state_out_4_0_5[2:0] ), //o
    .port_state_out_4_0_6  (mixColumns_port_state_out_4_0_6[2:0] ), //o
    .port_state_out_4_0_7  (mixColumns_port_state_out_4_0_7[2:0] ), //o
    .port_state_out_4_1_0  (mixColumns_port_state_out_4_1_0[2:0] ), //o
    .port_state_out_4_1_1  (mixColumns_port_state_out_4_1_1[2:0] ), //o
    .port_state_out_4_1_2  (mixColumns_port_state_out_4_1_2[2:0] ), //o
    .port_state_out_4_1_3  (mixColumns_port_state_out_4_1_3[2:0] ), //o
    .port_state_out_4_1_4  (mixColumns_port_state_out_4_1_4[2:0] ), //o
    .port_state_out_4_1_5  (mixColumns_port_state_out_4_1_5[2:0] ), //o
    .port_state_out_4_1_6  (mixColumns_port_state_out_4_1_6[2:0] ), //o
    .port_state_out_4_1_7  (mixColumns_port_state_out_4_1_7[2:0] ), //o
    .port_state_out_4_2_0  (mixColumns_port_state_out_4_2_0[2:0] ), //o
    .port_state_out_4_2_1  (mixColumns_port_state_out_4_2_1[2:0] ), //o
    .port_state_out_4_2_2  (mixColumns_port_state_out_4_2_2[2:0] ), //o
    .port_state_out_4_2_3  (mixColumns_port_state_out_4_2_3[2:0] ), //o
    .port_state_out_4_2_4  (mixColumns_port_state_out_4_2_4[2:0] ), //o
    .port_state_out_4_2_5  (mixColumns_port_state_out_4_2_5[2:0] ), //o
    .port_state_out_4_2_6  (mixColumns_port_state_out_4_2_6[2:0] ), //o
    .port_state_out_4_2_7  (mixColumns_port_state_out_4_2_7[2:0] ), //o
    .port_state_out_4_3_0  (mixColumns_port_state_out_4_3_0[2:0] ), //o
    .port_state_out_4_3_1  (mixColumns_port_state_out_4_3_1[2:0] ), //o
    .port_state_out_4_3_2  (mixColumns_port_state_out_4_3_2[2:0] ), //o
    .port_state_out_4_3_3  (mixColumns_port_state_out_4_3_3[2:0] ), //o
    .port_state_out_4_3_4  (mixColumns_port_state_out_4_3_4[2:0] ), //o
    .port_state_out_4_3_5  (mixColumns_port_state_out_4_3_5[2:0] ), //o
    .port_state_out_4_3_6  (mixColumns_port_state_out_4_3_6[2:0] ), //o
    .port_state_out_4_3_7  (mixColumns_port_state_out_4_3_7[2:0] ), //o
    .port_state_out_5_0_0  (mixColumns_port_state_out_5_0_0[2:0] ), //o
    .port_state_out_5_0_1  (mixColumns_port_state_out_5_0_1[2:0] ), //o
    .port_state_out_5_0_2  (mixColumns_port_state_out_5_0_2[2:0] ), //o
    .port_state_out_5_0_3  (mixColumns_port_state_out_5_0_3[2:0] ), //o
    .port_state_out_5_0_4  (mixColumns_port_state_out_5_0_4[2:0] ), //o
    .port_state_out_5_0_5  (mixColumns_port_state_out_5_0_5[2:0] ), //o
    .port_state_out_5_0_6  (mixColumns_port_state_out_5_0_6[2:0] ), //o
    .port_state_out_5_0_7  (mixColumns_port_state_out_5_0_7[2:0] ), //o
    .port_state_out_5_1_0  (mixColumns_port_state_out_5_1_0[2:0] ), //o
    .port_state_out_5_1_1  (mixColumns_port_state_out_5_1_1[2:0] ), //o
    .port_state_out_5_1_2  (mixColumns_port_state_out_5_1_2[2:0] ), //o
    .port_state_out_5_1_3  (mixColumns_port_state_out_5_1_3[2:0] ), //o
    .port_state_out_5_1_4  (mixColumns_port_state_out_5_1_4[2:0] ), //o
    .port_state_out_5_1_5  (mixColumns_port_state_out_5_1_5[2:0] ), //o
    .port_state_out_5_1_6  (mixColumns_port_state_out_5_1_6[2:0] ), //o
    .port_state_out_5_1_7  (mixColumns_port_state_out_5_1_7[2:0] ), //o
    .port_state_out_5_2_0  (mixColumns_port_state_out_5_2_0[2:0] ), //o
    .port_state_out_5_2_1  (mixColumns_port_state_out_5_2_1[2:0] ), //o
    .port_state_out_5_2_2  (mixColumns_port_state_out_5_2_2[2:0] ), //o
    .port_state_out_5_2_3  (mixColumns_port_state_out_5_2_3[2:0] ), //o
    .port_state_out_5_2_4  (mixColumns_port_state_out_5_2_4[2:0] ), //o
    .port_state_out_5_2_5  (mixColumns_port_state_out_5_2_5[2:0] ), //o
    .port_state_out_5_2_6  (mixColumns_port_state_out_5_2_6[2:0] ), //o
    .port_state_out_5_2_7  (mixColumns_port_state_out_5_2_7[2:0] ), //o
    .port_state_out_5_3_0  (mixColumns_port_state_out_5_3_0[2:0] ), //o
    .port_state_out_5_3_1  (mixColumns_port_state_out_5_3_1[2:0] ), //o
    .port_state_out_5_3_2  (mixColumns_port_state_out_5_3_2[2:0] ), //o
    .port_state_out_5_3_3  (mixColumns_port_state_out_5_3_3[2:0] ), //o
    .port_state_out_5_3_4  (mixColumns_port_state_out_5_3_4[2:0] ), //o
    .port_state_out_5_3_5  (mixColumns_port_state_out_5_3_5[2:0] ), //o
    .port_state_out_5_3_6  (mixColumns_port_state_out_5_3_6[2:0] ), //o
    .port_state_out_5_3_7  (mixColumns_port_state_out_5_3_7[2:0] ), //o
    .port_state_out_6_0_0  (mixColumns_port_state_out_6_0_0[2:0] ), //o
    .port_state_out_6_0_1  (mixColumns_port_state_out_6_0_1[2:0] ), //o
    .port_state_out_6_0_2  (mixColumns_port_state_out_6_0_2[2:0] ), //o
    .port_state_out_6_0_3  (mixColumns_port_state_out_6_0_3[2:0] ), //o
    .port_state_out_6_0_4  (mixColumns_port_state_out_6_0_4[2:0] ), //o
    .port_state_out_6_0_5  (mixColumns_port_state_out_6_0_5[2:0] ), //o
    .port_state_out_6_0_6  (mixColumns_port_state_out_6_0_6[2:0] ), //o
    .port_state_out_6_0_7  (mixColumns_port_state_out_6_0_7[2:0] ), //o
    .port_state_out_6_1_0  (mixColumns_port_state_out_6_1_0[2:0] ), //o
    .port_state_out_6_1_1  (mixColumns_port_state_out_6_1_1[2:0] ), //o
    .port_state_out_6_1_2  (mixColumns_port_state_out_6_1_2[2:0] ), //o
    .port_state_out_6_1_3  (mixColumns_port_state_out_6_1_3[2:0] ), //o
    .port_state_out_6_1_4  (mixColumns_port_state_out_6_1_4[2:0] ), //o
    .port_state_out_6_1_5  (mixColumns_port_state_out_6_1_5[2:0] ), //o
    .port_state_out_6_1_6  (mixColumns_port_state_out_6_1_6[2:0] ), //o
    .port_state_out_6_1_7  (mixColumns_port_state_out_6_1_7[2:0] ), //o
    .port_state_out_6_2_0  (mixColumns_port_state_out_6_2_0[2:0] ), //o
    .port_state_out_6_2_1  (mixColumns_port_state_out_6_2_1[2:0] ), //o
    .port_state_out_6_2_2  (mixColumns_port_state_out_6_2_2[2:0] ), //o
    .port_state_out_6_2_3  (mixColumns_port_state_out_6_2_3[2:0] ), //o
    .port_state_out_6_2_4  (mixColumns_port_state_out_6_2_4[2:0] ), //o
    .port_state_out_6_2_5  (mixColumns_port_state_out_6_2_5[2:0] ), //o
    .port_state_out_6_2_6  (mixColumns_port_state_out_6_2_6[2:0] ), //o
    .port_state_out_6_2_7  (mixColumns_port_state_out_6_2_7[2:0] ), //o
    .port_state_out_6_3_0  (mixColumns_port_state_out_6_3_0[2:0] ), //o
    .port_state_out_6_3_1  (mixColumns_port_state_out_6_3_1[2:0] ), //o
    .port_state_out_6_3_2  (mixColumns_port_state_out_6_3_2[2:0] ), //o
    .port_state_out_6_3_3  (mixColumns_port_state_out_6_3_3[2:0] ), //o
    .port_state_out_6_3_4  (mixColumns_port_state_out_6_3_4[2:0] ), //o
    .port_state_out_6_3_5  (mixColumns_port_state_out_6_3_5[2:0] ), //o
    .port_state_out_6_3_6  (mixColumns_port_state_out_6_3_6[2:0] ), //o
    .port_state_out_6_3_7  (mixColumns_port_state_out_6_3_7[2:0] ), //o
    .port_state_out_7_0_0  (mixColumns_port_state_out_7_0_0[2:0] ), //o
    .port_state_out_7_0_1  (mixColumns_port_state_out_7_0_1[2:0] ), //o
    .port_state_out_7_0_2  (mixColumns_port_state_out_7_0_2[2:0] ), //o
    .port_state_out_7_0_3  (mixColumns_port_state_out_7_0_3[2:0] ), //o
    .port_state_out_7_0_4  (mixColumns_port_state_out_7_0_4[2:0] ), //o
    .port_state_out_7_0_5  (mixColumns_port_state_out_7_0_5[2:0] ), //o
    .port_state_out_7_0_6  (mixColumns_port_state_out_7_0_6[2:0] ), //o
    .port_state_out_7_0_7  (mixColumns_port_state_out_7_0_7[2:0] ), //o
    .port_state_out_7_1_0  (mixColumns_port_state_out_7_1_0[2:0] ), //o
    .port_state_out_7_1_1  (mixColumns_port_state_out_7_1_1[2:0] ), //o
    .port_state_out_7_1_2  (mixColumns_port_state_out_7_1_2[2:0] ), //o
    .port_state_out_7_1_3  (mixColumns_port_state_out_7_1_3[2:0] ), //o
    .port_state_out_7_1_4  (mixColumns_port_state_out_7_1_4[2:0] ), //o
    .port_state_out_7_1_5  (mixColumns_port_state_out_7_1_5[2:0] ), //o
    .port_state_out_7_1_6  (mixColumns_port_state_out_7_1_6[2:0] ), //o
    .port_state_out_7_1_7  (mixColumns_port_state_out_7_1_7[2:0] ), //o
    .port_state_out_7_2_0  (mixColumns_port_state_out_7_2_0[2:0] ), //o
    .port_state_out_7_2_1  (mixColumns_port_state_out_7_2_1[2:0] ), //o
    .port_state_out_7_2_2  (mixColumns_port_state_out_7_2_2[2:0] ), //o
    .port_state_out_7_2_3  (mixColumns_port_state_out_7_2_3[2:0] ), //o
    .port_state_out_7_2_4  (mixColumns_port_state_out_7_2_4[2:0] ), //o
    .port_state_out_7_2_5  (mixColumns_port_state_out_7_2_5[2:0] ), //o
    .port_state_out_7_2_6  (mixColumns_port_state_out_7_2_6[2:0] ), //o
    .port_state_out_7_2_7  (mixColumns_port_state_out_7_2_7[2:0] ), //o
    .port_state_out_7_3_0  (mixColumns_port_state_out_7_3_0[2:0] ), //o
    .port_state_out_7_3_1  (mixColumns_port_state_out_7_3_1[2:0] ), //o
    .port_state_out_7_3_2  (mixColumns_port_state_out_7_3_2[2:0] ), //o
    .port_state_out_7_3_3  (mixColumns_port_state_out_7_3_3[2:0] ), //o
    .port_state_out_7_3_4  (mixColumns_port_state_out_7_3_4[2:0] ), //o
    .port_state_out_7_3_5  (mixColumns_port_state_out_7_3_5[2:0] ), //o
    .port_state_out_7_3_6  (mixColumns_port_state_out_7_3_6[2:0] ), //o
    .port_state_out_7_3_7  (mixColumns_port_state_out_7_3_7[2:0] ), //o
    .port_state_out_8_0_0  (mixColumns_port_state_out_8_0_0[2:0] ), //o
    .port_state_out_8_0_1  (mixColumns_port_state_out_8_0_1[2:0] ), //o
    .port_state_out_8_0_2  (mixColumns_port_state_out_8_0_2[2:0] ), //o
    .port_state_out_8_0_3  (mixColumns_port_state_out_8_0_3[2:0] ), //o
    .port_state_out_8_0_4  (mixColumns_port_state_out_8_0_4[2:0] ), //o
    .port_state_out_8_0_5  (mixColumns_port_state_out_8_0_5[2:0] ), //o
    .port_state_out_8_0_6  (mixColumns_port_state_out_8_0_6[2:0] ), //o
    .port_state_out_8_0_7  (mixColumns_port_state_out_8_0_7[2:0] ), //o
    .port_state_out_8_1_0  (mixColumns_port_state_out_8_1_0[2:0] ), //o
    .port_state_out_8_1_1  (mixColumns_port_state_out_8_1_1[2:0] ), //o
    .port_state_out_8_1_2  (mixColumns_port_state_out_8_1_2[2:0] ), //o
    .port_state_out_8_1_3  (mixColumns_port_state_out_8_1_3[2:0] ), //o
    .port_state_out_8_1_4  (mixColumns_port_state_out_8_1_4[2:0] ), //o
    .port_state_out_8_1_5  (mixColumns_port_state_out_8_1_5[2:0] ), //o
    .port_state_out_8_1_6  (mixColumns_port_state_out_8_1_6[2:0] ), //o
    .port_state_out_8_1_7  (mixColumns_port_state_out_8_1_7[2:0] ), //o
    .port_state_out_8_2_0  (mixColumns_port_state_out_8_2_0[2:0] ), //o
    .port_state_out_8_2_1  (mixColumns_port_state_out_8_2_1[2:0] ), //o
    .port_state_out_8_2_2  (mixColumns_port_state_out_8_2_2[2:0] ), //o
    .port_state_out_8_2_3  (mixColumns_port_state_out_8_2_3[2:0] ), //o
    .port_state_out_8_2_4  (mixColumns_port_state_out_8_2_4[2:0] ), //o
    .port_state_out_8_2_5  (mixColumns_port_state_out_8_2_5[2:0] ), //o
    .port_state_out_8_2_6  (mixColumns_port_state_out_8_2_6[2:0] ), //o
    .port_state_out_8_2_7  (mixColumns_port_state_out_8_2_7[2:0] ), //o
    .port_state_out_8_3_0  (mixColumns_port_state_out_8_3_0[2:0] ), //o
    .port_state_out_8_3_1  (mixColumns_port_state_out_8_3_1[2:0] ), //o
    .port_state_out_8_3_2  (mixColumns_port_state_out_8_3_2[2:0] ), //o
    .port_state_out_8_3_3  (mixColumns_port_state_out_8_3_3[2:0] ), //o
    .port_state_out_8_3_4  (mixColumns_port_state_out_8_3_4[2:0] ), //o
    .port_state_out_8_3_5  (mixColumns_port_state_out_8_3_5[2:0] ), //o
    .port_state_out_8_3_6  (mixColumns_port_state_out_8_3_6[2:0] ), //o
    .port_state_out_8_3_7  (mixColumns_port_state_out_8_3_7[2:0] ), //o
    .port_state_out_9_0_0  (mixColumns_port_state_out_9_0_0[2:0] ), //o
    .port_state_out_9_0_1  (mixColumns_port_state_out_9_0_1[2:0] ), //o
    .port_state_out_9_0_2  (mixColumns_port_state_out_9_0_2[2:0] ), //o
    .port_state_out_9_0_3  (mixColumns_port_state_out_9_0_3[2:0] ), //o
    .port_state_out_9_0_4  (mixColumns_port_state_out_9_0_4[2:0] ), //o
    .port_state_out_9_0_5  (mixColumns_port_state_out_9_0_5[2:0] ), //o
    .port_state_out_9_0_6  (mixColumns_port_state_out_9_0_6[2:0] ), //o
    .port_state_out_9_0_7  (mixColumns_port_state_out_9_0_7[2:0] ), //o
    .port_state_out_9_1_0  (mixColumns_port_state_out_9_1_0[2:0] ), //o
    .port_state_out_9_1_1  (mixColumns_port_state_out_9_1_1[2:0] ), //o
    .port_state_out_9_1_2  (mixColumns_port_state_out_9_1_2[2:0] ), //o
    .port_state_out_9_1_3  (mixColumns_port_state_out_9_1_3[2:0] ), //o
    .port_state_out_9_1_4  (mixColumns_port_state_out_9_1_4[2:0] ), //o
    .port_state_out_9_1_5  (mixColumns_port_state_out_9_1_5[2:0] ), //o
    .port_state_out_9_1_6  (mixColumns_port_state_out_9_1_6[2:0] ), //o
    .port_state_out_9_1_7  (mixColumns_port_state_out_9_1_7[2:0] ), //o
    .port_state_out_9_2_0  (mixColumns_port_state_out_9_2_0[2:0] ), //o
    .port_state_out_9_2_1  (mixColumns_port_state_out_9_2_1[2:0] ), //o
    .port_state_out_9_2_2  (mixColumns_port_state_out_9_2_2[2:0] ), //o
    .port_state_out_9_2_3  (mixColumns_port_state_out_9_2_3[2:0] ), //o
    .port_state_out_9_2_4  (mixColumns_port_state_out_9_2_4[2:0] ), //o
    .port_state_out_9_2_5  (mixColumns_port_state_out_9_2_5[2:0] ), //o
    .port_state_out_9_2_6  (mixColumns_port_state_out_9_2_6[2:0] ), //o
    .port_state_out_9_2_7  (mixColumns_port_state_out_9_2_7[2:0] ), //o
    .port_state_out_9_3_0  (mixColumns_port_state_out_9_3_0[2:0] ), //o
    .port_state_out_9_3_1  (mixColumns_port_state_out_9_3_1[2:0] ), //o
    .port_state_out_9_3_2  (mixColumns_port_state_out_9_3_2[2:0] ), //o
    .port_state_out_9_3_3  (mixColumns_port_state_out_9_3_3[2:0] ), //o
    .port_state_out_9_3_4  (mixColumns_port_state_out_9_3_4[2:0] ), //o
    .port_state_out_9_3_5  (mixColumns_port_state_out_9_3_5[2:0] ), //o
    .port_state_out_9_3_6  (mixColumns_port_state_out_9_3_6[2:0] ), //o
    .port_state_out_9_3_7  (mixColumns_port_state_out_9_3_7[2:0] ), //o
    .port_state_out_10_0_0 (mixColumns_port_state_out_10_0_0[2:0]), //o
    .port_state_out_10_0_1 (mixColumns_port_state_out_10_0_1[2:0]), //o
    .port_state_out_10_0_2 (mixColumns_port_state_out_10_0_2[2:0]), //o
    .port_state_out_10_0_3 (mixColumns_port_state_out_10_0_3[2:0]), //o
    .port_state_out_10_0_4 (mixColumns_port_state_out_10_0_4[2:0]), //o
    .port_state_out_10_0_5 (mixColumns_port_state_out_10_0_5[2:0]), //o
    .port_state_out_10_0_6 (mixColumns_port_state_out_10_0_6[2:0]), //o
    .port_state_out_10_0_7 (mixColumns_port_state_out_10_0_7[2:0]), //o
    .port_state_out_10_1_0 (mixColumns_port_state_out_10_1_0[2:0]), //o
    .port_state_out_10_1_1 (mixColumns_port_state_out_10_1_1[2:0]), //o
    .port_state_out_10_1_2 (mixColumns_port_state_out_10_1_2[2:0]), //o
    .port_state_out_10_1_3 (mixColumns_port_state_out_10_1_3[2:0]), //o
    .port_state_out_10_1_4 (mixColumns_port_state_out_10_1_4[2:0]), //o
    .port_state_out_10_1_5 (mixColumns_port_state_out_10_1_5[2:0]), //o
    .port_state_out_10_1_6 (mixColumns_port_state_out_10_1_6[2:0]), //o
    .port_state_out_10_1_7 (mixColumns_port_state_out_10_1_7[2:0]), //o
    .port_state_out_10_2_0 (mixColumns_port_state_out_10_2_0[2:0]), //o
    .port_state_out_10_2_1 (mixColumns_port_state_out_10_2_1[2:0]), //o
    .port_state_out_10_2_2 (mixColumns_port_state_out_10_2_2[2:0]), //o
    .port_state_out_10_2_3 (mixColumns_port_state_out_10_2_3[2:0]), //o
    .port_state_out_10_2_4 (mixColumns_port_state_out_10_2_4[2:0]), //o
    .port_state_out_10_2_5 (mixColumns_port_state_out_10_2_5[2:0]), //o
    .port_state_out_10_2_6 (mixColumns_port_state_out_10_2_6[2:0]), //o
    .port_state_out_10_2_7 (mixColumns_port_state_out_10_2_7[2:0]), //o
    .port_state_out_10_3_0 (mixColumns_port_state_out_10_3_0[2:0]), //o
    .port_state_out_10_3_1 (mixColumns_port_state_out_10_3_1[2:0]), //o
    .port_state_out_10_3_2 (mixColumns_port_state_out_10_3_2[2:0]), //o
    .port_state_out_10_3_3 (mixColumns_port_state_out_10_3_3[2:0]), //o
    .port_state_out_10_3_4 (mixColumns_port_state_out_10_3_4[2:0]), //o
    .port_state_out_10_3_5 (mixColumns_port_state_out_10_3_5[2:0]), //o
    .port_state_out_10_3_6 (mixColumns_port_state_out_10_3_6[2:0]), //o
    .port_state_out_10_3_7 (mixColumns_port_state_out_10_3_7[2:0]), //o
    .port_state_out_11_0_0 (mixColumns_port_state_out_11_0_0[2:0]), //o
    .port_state_out_11_0_1 (mixColumns_port_state_out_11_0_1[2:0]), //o
    .port_state_out_11_0_2 (mixColumns_port_state_out_11_0_2[2:0]), //o
    .port_state_out_11_0_3 (mixColumns_port_state_out_11_0_3[2:0]), //o
    .port_state_out_11_0_4 (mixColumns_port_state_out_11_0_4[2:0]), //o
    .port_state_out_11_0_5 (mixColumns_port_state_out_11_0_5[2:0]), //o
    .port_state_out_11_0_6 (mixColumns_port_state_out_11_0_6[2:0]), //o
    .port_state_out_11_0_7 (mixColumns_port_state_out_11_0_7[2:0]), //o
    .port_state_out_11_1_0 (mixColumns_port_state_out_11_1_0[2:0]), //o
    .port_state_out_11_1_1 (mixColumns_port_state_out_11_1_1[2:0]), //o
    .port_state_out_11_1_2 (mixColumns_port_state_out_11_1_2[2:0]), //o
    .port_state_out_11_1_3 (mixColumns_port_state_out_11_1_3[2:0]), //o
    .port_state_out_11_1_4 (mixColumns_port_state_out_11_1_4[2:0]), //o
    .port_state_out_11_1_5 (mixColumns_port_state_out_11_1_5[2:0]), //o
    .port_state_out_11_1_6 (mixColumns_port_state_out_11_1_6[2:0]), //o
    .port_state_out_11_1_7 (mixColumns_port_state_out_11_1_7[2:0]), //o
    .port_state_out_11_2_0 (mixColumns_port_state_out_11_2_0[2:0]), //o
    .port_state_out_11_2_1 (mixColumns_port_state_out_11_2_1[2:0]), //o
    .port_state_out_11_2_2 (mixColumns_port_state_out_11_2_2[2:0]), //o
    .port_state_out_11_2_3 (mixColumns_port_state_out_11_2_3[2:0]), //o
    .port_state_out_11_2_4 (mixColumns_port_state_out_11_2_4[2:0]), //o
    .port_state_out_11_2_5 (mixColumns_port_state_out_11_2_5[2:0]), //o
    .port_state_out_11_2_6 (mixColumns_port_state_out_11_2_6[2:0]), //o
    .port_state_out_11_2_7 (mixColumns_port_state_out_11_2_7[2:0]), //o
    .port_state_out_11_3_0 (mixColumns_port_state_out_11_3_0[2:0]), //o
    .port_state_out_11_3_1 (mixColumns_port_state_out_11_3_1[2:0]), //o
    .port_state_out_11_3_2 (mixColumns_port_state_out_11_3_2[2:0]), //o
    .port_state_out_11_3_3 (mixColumns_port_state_out_11_3_3[2:0]), //o
    .port_state_out_11_3_4 (mixColumns_port_state_out_11_3_4[2:0]), //o
    .port_state_out_11_3_5 (mixColumns_port_state_out_11_3_5[2:0]), //o
    .port_state_out_11_3_6 (mixColumns_port_state_out_11_3_6[2:0]), //o
    .port_state_out_11_3_7 (mixColumns_port_state_out_11_3_7[2:0]), //o
    .port_state_out_12_0_0 (mixColumns_port_state_out_12_0_0[2:0]), //o
    .port_state_out_12_0_1 (mixColumns_port_state_out_12_0_1[2:0]), //o
    .port_state_out_12_0_2 (mixColumns_port_state_out_12_0_2[2:0]), //o
    .port_state_out_12_0_3 (mixColumns_port_state_out_12_0_3[2:0]), //o
    .port_state_out_12_0_4 (mixColumns_port_state_out_12_0_4[2:0]), //o
    .port_state_out_12_0_5 (mixColumns_port_state_out_12_0_5[2:0]), //o
    .port_state_out_12_0_6 (mixColumns_port_state_out_12_0_6[2:0]), //o
    .port_state_out_12_0_7 (mixColumns_port_state_out_12_0_7[2:0]), //o
    .port_state_out_12_1_0 (mixColumns_port_state_out_12_1_0[2:0]), //o
    .port_state_out_12_1_1 (mixColumns_port_state_out_12_1_1[2:0]), //o
    .port_state_out_12_1_2 (mixColumns_port_state_out_12_1_2[2:0]), //o
    .port_state_out_12_1_3 (mixColumns_port_state_out_12_1_3[2:0]), //o
    .port_state_out_12_1_4 (mixColumns_port_state_out_12_1_4[2:0]), //o
    .port_state_out_12_1_5 (mixColumns_port_state_out_12_1_5[2:0]), //o
    .port_state_out_12_1_6 (mixColumns_port_state_out_12_1_6[2:0]), //o
    .port_state_out_12_1_7 (mixColumns_port_state_out_12_1_7[2:0]), //o
    .port_state_out_12_2_0 (mixColumns_port_state_out_12_2_0[2:0]), //o
    .port_state_out_12_2_1 (mixColumns_port_state_out_12_2_1[2:0]), //o
    .port_state_out_12_2_2 (mixColumns_port_state_out_12_2_2[2:0]), //o
    .port_state_out_12_2_3 (mixColumns_port_state_out_12_2_3[2:0]), //o
    .port_state_out_12_2_4 (mixColumns_port_state_out_12_2_4[2:0]), //o
    .port_state_out_12_2_5 (mixColumns_port_state_out_12_2_5[2:0]), //o
    .port_state_out_12_2_6 (mixColumns_port_state_out_12_2_6[2:0]), //o
    .port_state_out_12_2_7 (mixColumns_port_state_out_12_2_7[2:0]), //o
    .port_state_out_12_3_0 (mixColumns_port_state_out_12_3_0[2:0]), //o
    .port_state_out_12_3_1 (mixColumns_port_state_out_12_3_1[2:0]), //o
    .port_state_out_12_3_2 (mixColumns_port_state_out_12_3_2[2:0]), //o
    .port_state_out_12_3_3 (mixColumns_port_state_out_12_3_3[2:0]), //o
    .port_state_out_12_3_4 (mixColumns_port_state_out_12_3_4[2:0]), //o
    .port_state_out_12_3_5 (mixColumns_port_state_out_12_3_5[2:0]), //o
    .port_state_out_12_3_6 (mixColumns_port_state_out_12_3_6[2:0]), //o
    .port_state_out_12_3_7 (mixColumns_port_state_out_12_3_7[2:0]), //o
    .port_state_out_13_0_0 (mixColumns_port_state_out_13_0_0[2:0]), //o
    .port_state_out_13_0_1 (mixColumns_port_state_out_13_0_1[2:0]), //o
    .port_state_out_13_0_2 (mixColumns_port_state_out_13_0_2[2:0]), //o
    .port_state_out_13_0_3 (mixColumns_port_state_out_13_0_3[2:0]), //o
    .port_state_out_13_0_4 (mixColumns_port_state_out_13_0_4[2:0]), //o
    .port_state_out_13_0_5 (mixColumns_port_state_out_13_0_5[2:0]), //o
    .port_state_out_13_0_6 (mixColumns_port_state_out_13_0_6[2:0]), //o
    .port_state_out_13_0_7 (mixColumns_port_state_out_13_0_7[2:0]), //o
    .port_state_out_13_1_0 (mixColumns_port_state_out_13_1_0[2:0]), //o
    .port_state_out_13_1_1 (mixColumns_port_state_out_13_1_1[2:0]), //o
    .port_state_out_13_1_2 (mixColumns_port_state_out_13_1_2[2:0]), //o
    .port_state_out_13_1_3 (mixColumns_port_state_out_13_1_3[2:0]), //o
    .port_state_out_13_1_4 (mixColumns_port_state_out_13_1_4[2:0]), //o
    .port_state_out_13_1_5 (mixColumns_port_state_out_13_1_5[2:0]), //o
    .port_state_out_13_1_6 (mixColumns_port_state_out_13_1_6[2:0]), //o
    .port_state_out_13_1_7 (mixColumns_port_state_out_13_1_7[2:0]), //o
    .port_state_out_13_2_0 (mixColumns_port_state_out_13_2_0[2:0]), //o
    .port_state_out_13_2_1 (mixColumns_port_state_out_13_2_1[2:0]), //o
    .port_state_out_13_2_2 (mixColumns_port_state_out_13_2_2[2:0]), //o
    .port_state_out_13_2_3 (mixColumns_port_state_out_13_2_3[2:0]), //o
    .port_state_out_13_2_4 (mixColumns_port_state_out_13_2_4[2:0]), //o
    .port_state_out_13_2_5 (mixColumns_port_state_out_13_2_5[2:0]), //o
    .port_state_out_13_2_6 (mixColumns_port_state_out_13_2_6[2:0]), //o
    .port_state_out_13_2_7 (mixColumns_port_state_out_13_2_7[2:0]), //o
    .port_state_out_13_3_0 (mixColumns_port_state_out_13_3_0[2:0]), //o
    .port_state_out_13_3_1 (mixColumns_port_state_out_13_3_1[2:0]), //o
    .port_state_out_13_3_2 (mixColumns_port_state_out_13_3_2[2:0]), //o
    .port_state_out_13_3_3 (mixColumns_port_state_out_13_3_3[2:0]), //o
    .port_state_out_13_3_4 (mixColumns_port_state_out_13_3_4[2:0]), //o
    .port_state_out_13_3_5 (mixColumns_port_state_out_13_3_5[2:0]), //o
    .port_state_out_13_3_6 (mixColumns_port_state_out_13_3_6[2:0]), //o
    .port_state_out_13_3_7 (mixColumns_port_state_out_13_3_7[2:0]), //o
    .port_state_out_14_0_0 (mixColumns_port_state_out_14_0_0[2:0]), //o
    .port_state_out_14_0_1 (mixColumns_port_state_out_14_0_1[2:0]), //o
    .port_state_out_14_0_2 (mixColumns_port_state_out_14_0_2[2:0]), //o
    .port_state_out_14_0_3 (mixColumns_port_state_out_14_0_3[2:0]), //o
    .port_state_out_14_0_4 (mixColumns_port_state_out_14_0_4[2:0]), //o
    .port_state_out_14_0_5 (mixColumns_port_state_out_14_0_5[2:0]), //o
    .port_state_out_14_0_6 (mixColumns_port_state_out_14_0_6[2:0]), //o
    .port_state_out_14_0_7 (mixColumns_port_state_out_14_0_7[2:0]), //o
    .port_state_out_14_1_0 (mixColumns_port_state_out_14_1_0[2:0]), //o
    .port_state_out_14_1_1 (mixColumns_port_state_out_14_1_1[2:0]), //o
    .port_state_out_14_1_2 (mixColumns_port_state_out_14_1_2[2:0]), //o
    .port_state_out_14_1_3 (mixColumns_port_state_out_14_1_3[2:0]), //o
    .port_state_out_14_1_4 (mixColumns_port_state_out_14_1_4[2:0]), //o
    .port_state_out_14_1_5 (mixColumns_port_state_out_14_1_5[2:0]), //o
    .port_state_out_14_1_6 (mixColumns_port_state_out_14_1_6[2:0]), //o
    .port_state_out_14_1_7 (mixColumns_port_state_out_14_1_7[2:0]), //o
    .port_state_out_14_2_0 (mixColumns_port_state_out_14_2_0[2:0]), //o
    .port_state_out_14_2_1 (mixColumns_port_state_out_14_2_1[2:0]), //o
    .port_state_out_14_2_2 (mixColumns_port_state_out_14_2_2[2:0]), //o
    .port_state_out_14_2_3 (mixColumns_port_state_out_14_2_3[2:0]), //o
    .port_state_out_14_2_4 (mixColumns_port_state_out_14_2_4[2:0]), //o
    .port_state_out_14_2_5 (mixColumns_port_state_out_14_2_5[2:0]), //o
    .port_state_out_14_2_6 (mixColumns_port_state_out_14_2_6[2:0]), //o
    .port_state_out_14_2_7 (mixColumns_port_state_out_14_2_7[2:0]), //o
    .port_state_out_14_3_0 (mixColumns_port_state_out_14_3_0[2:0]), //o
    .port_state_out_14_3_1 (mixColumns_port_state_out_14_3_1[2:0]), //o
    .port_state_out_14_3_2 (mixColumns_port_state_out_14_3_2[2:0]), //o
    .port_state_out_14_3_3 (mixColumns_port_state_out_14_3_3[2:0]), //o
    .port_state_out_14_3_4 (mixColumns_port_state_out_14_3_4[2:0]), //o
    .port_state_out_14_3_5 (mixColumns_port_state_out_14_3_5[2:0]), //o
    .port_state_out_14_3_6 (mixColumns_port_state_out_14_3_6[2:0]), //o
    .port_state_out_14_3_7 (mixColumns_port_state_out_14_3_7[2:0]), //o
    .port_state_out_15_0_0 (mixColumns_port_state_out_15_0_0[2:0]), //o
    .port_state_out_15_0_1 (mixColumns_port_state_out_15_0_1[2:0]), //o
    .port_state_out_15_0_2 (mixColumns_port_state_out_15_0_2[2:0]), //o
    .port_state_out_15_0_3 (mixColumns_port_state_out_15_0_3[2:0]), //o
    .port_state_out_15_0_4 (mixColumns_port_state_out_15_0_4[2:0]), //o
    .port_state_out_15_0_5 (mixColumns_port_state_out_15_0_5[2:0]), //o
    .port_state_out_15_0_6 (mixColumns_port_state_out_15_0_6[2:0]), //o
    .port_state_out_15_0_7 (mixColumns_port_state_out_15_0_7[2:0]), //o
    .port_state_out_15_1_0 (mixColumns_port_state_out_15_1_0[2:0]), //o
    .port_state_out_15_1_1 (mixColumns_port_state_out_15_1_1[2:0]), //o
    .port_state_out_15_1_2 (mixColumns_port_state_out_15_1_2[2:0]), //o
    .port_state_out_15_1_3 (mixColumns_port_state_out_15_1_3[2:0]), //o
    .port_state_out_15_1_4 (mixColumns_port_state_out_15_1_4[2:0]), //o
    .port_state_out_15_1_5 (mixColumns_port_state_out_15_1_5[2:0]), //o
    .port_state_out_15_1_6 (mixColumns_port_state_out_15_1_6[2:0]), //o
    .port_state_out_15_1_7 (mixColumns_port_state_out_15_1_7[2:0]), //o
    .port_state_out_15_2_0 (mixColumns_port_state_out_15_2_0[2:0]), //o
    .port_state_out_15_2_1 (mixColumns_port_state_out_15_2_1[2:0]), //o
    .port_state_out_15_2_2 (mixColumns_port_state_out_15_2_2[2:0]), //o
    .port_state_out_15_2_3 (mixColumns_port_state_out_15_2_3[2:0]), //o
    .port_state_out_15_2_4 (mixColumns_port_state_out_15_2_4[2:0]), //o
    .port_state_out_15_2_5 (mixColumns_port_state_out_15_2_5[2:0]), //o
    .port_state_out_15_2_6 (mixColumns_port_state_out_15_2_6[2:0]), //o
    .port_state_out_15_2_7 (mixColumns_port_state_out_15_2_7[2:0]), //o
    .port_state_out_15_3_0 (mixColumns_port_state_out_15_3_0[2:0]), //o
    .port_state_out_15_3_1 (mixColumns_port_state_out_15_3_1[2:0]), //o
    .port_state_out_15_3_2 (mixColumns_port_state_out_15_3_2[2:0]), //o
    .port_state_out_15_3_3 (mixColumns_port_state_out_15_3_3[2:0]), //o
    .port_state_out_15_3_4 (mixColumns_port_state_out_15_3_4[2:0]), //o
    .port_state_out_15_3_5 (mixColumns_port_state_out_15_3_5[2:0]), //o
    .port_state_out_15_3_6 (mixColumns_port_state_out_15_3_6[2:0]), //o
    .port_state_out_15_3_7 (mixColumns_port_state_out_15_3_7[2:0])  //o
  );
  Majority majority_4608 (
    .port_i (mixColumns_port_state_out_0_0_0[2:0]), //i
    .port_o (majority_4608_port_o                )  //o
  );
  Majority majority_4609 (
    .port_i (mixColumns_port_state_out_1_0_0[2:0]), //i
    .port_o (majority_4609_port_o                )  //o
  );
  Majority majority_4610 (
    .port_i (mixColumns_port_state_out_2_0_0[2:0]), //i
    .port_o (majority_4610_port_o                )  //o
  );
  Majority majority_4611 (
    .port_i (mixColumns_port_state_out_3_0_0[2:0]), //i
    .port_o (majority_4611_port_o                )  //o
  );
  Majority majority_4612 (
    .port_i (mixColumns_port_state_out_4_0_0[2:0]), //i
    .port_o (majority_4612_port_o                )  //o
  );
  Majority majority_4613 (
    .port_i (mixColumns_port_state_out_5_0_0[2:0]), //i
    .port_o (majority_4613_port_o                )  //o
  );
  Majority majority_4614 (
    .port_i (mixColumns_port_state_out_6_0_0[2:0]), //i
    .port_o (majority_4614_port_o                )  //o
  );
  Majority majority_4615 (
    .port_i (mixColumns_port_state_out_7_0_0[2:0]), //i
    .port_o (majority_4615_port_o                )  //o
  );
  Majority majority_4616 (
    .port_i (mixColumns_port_state_out_8_0_0[2:0]), //i
    .port_o (majority_4616_port_o                )  //o
  );
  Majority majority_4617 (
    .port_i (mixColumns_port_state_out_9_0_0[2:0]), //i
    .port_o (majority_4617_port_o                )  //o
  );
  Majority majority_4618 (
    .port_i (mixColumns_port_state_out_10_0_0[2:0]), //i
    .port_o (majority_4618_port_o                 )  //o
  );
  Majority majority_4619 (
    .port_i (mixColumns_port_state_out_11_0_0[2:0]), //i
    .port_o (majority_4619_port_o                 )  //o
  );
  Majority majority_4620 (
    .port_i (mixColumns_port_state_out_12_0_0[2:0]), //i
    .port_o (majority_4620_port_o                 )  //o
  );
  Majority majority_4621 (
    .port_i (mixColumns_port_state_out_13_0_0[2:0]), //i
    .port_o (majority_4621_port_o                 )  //o
  );
  Majority majority_4622 (
    .port_i (mixColumns_port_state_out_14_0_0[2:0]), //i
    .port_o (majority_4622_port_o                 )  //o
  );
  Majority majority_4623 (
    .port_i (mixColumns_port_state_out_15_0_0[2:0]), //i
    .port_o (majority_4623_port_o                 )  //o
  );
  Majority majority_4624 (
    .port_i (mixColumns_port_state_out_0_1_0[2:0]), //i
    .port_o (majority_4624_port_o                )  //o
  );
  Majority majority_4625 (
    .port_i (mixColumns_port_state_out_1_1_0[2:0]), //i
    .port_o (majority_4625_port_o                )  //o
  );
  Majority majority_4626 (
    .port_i (mixColumns_port_state_out_2_1_0[2:0]), //i
    .port_o (majority_4626_port_o                )  //o
  );
  Majority majority_4627 (
    .port_i (mixColumns_port_state_out_3_1_0[2:0]), //i
    .port_o (majority_4627_port_o                )  //o
  );
  Majority majority_4628 (
    .port_i (mixColumns_port_state_out_4_1_0[2:0]), //i
    .port_o (majority_4628_port_o                )  //o
  );
  Majority majority_4629 (
    .port_i (mixColumns_port_state_out_5_1_0[2:0]), //i
    .port_o (majority_4629_port_o                )  //o
  );
  Majority majority_4630 (
    .port_i (mixColumns_port_state_out_6_1_0[2:0]), //i
    .port_o (majority_4630_port_o                )  //o
  );
  Majority majority_4631 (
    .port_i (mixColumns_port_state_out_7_1_0[2:0]), //i
    .port_o (majority_4631_port_o                )  //o
  );
  Majority majority_4632 (
    .port_i (mixColumns_port_state_out_8_1_0[2:0]), //i
    .port_o (majority_4632_port_o                )  //o
  );
  Majority majority_4633 (
    .port_i (mixColumns_port_state_out_9_1_0[2:0]), //i
    .port_o (majority_4633_port_o                )  //o
  );
  Majority majority_4634 (
    .port_i (mixColumns_port_state_out_10_1_0[2:0]), //i
    .port_o (majority_4634_port_o                 )  //o
  );
  Majority majority_4635 (
    .port_i (mixColumns_port_state_out_11_1_0[2:0]), //i
    .port_o (majority_4635_port_o                 )  //o
  );
  Majority majority_4636 (
    .port_i (mixColumns_port_state_out_12_1_0[2:0]), //i
    .port_o (majority_4636_port_o                 )  //o
  );
  Majority majority_4637 (
    .port_i (mixColumns_port_state_out_13_1_0[2:0]), //i
    .port_o (majority_4637_port_o                 )  //o
  );
  Majority majority_4638 (
    .port_i (mixColumns_port_state_out_14_1_0[2:0]), //i
    .port_o (majority_4638_port_o                 )  //o
  );
  Majority majority_4639 (
    .port_i (mixColumns_port_state_out_15_1_0[2:0]), //i
    .port_o (majority_4639_port_o                 )  //o
  );
  Majority majority_4640 (
    .port_i (mixColumns_port_state_out_0_2_0[2:0]), //i
    .port_o (majority_4640_port_o                )  //o
  );
  Majority majority_4641 (
    .port_i (mixColumns_port_state_out_1_2_0[2:0]), //i
    .port_o (majority_4641_port_o                )  //o
  );
  Majority majority_4642 (
    .port_i (mixColumns_port_state_out_2_2_0[2:0]), //i
    .port_o (majority_4642_port_o                )  //o
  );
  Majority majority_4643 (
    .port_i (mixColumns_port_state_out_3_2_0[2:0]), //i
    .port_o (majority_4643_port_o                )  //o
  );
  Majority majority_4644 (
    .port_i (mixColumns_port_state_out_4_2_0[2:0]), //i
    .port_o (majority_4644_port_o                )  //o
  );
  Majority majority_4645 (
    .port_i (mixColumns_port_state_out_5_2_0[2:0]), //i
    .port_o (majority_4645_port_o                )  //o
  );
  Majority majority_4646 (
    .port_i (mixColumns_port_state_out_6_2_0[2:0]), //i
    .port_o (majority_4646_port_o                )  //o
  );
  Majority majority_4647 (
    .port_i (mixColumns_port_state_out_7_2_0[2:0]), //i
    .port_o (majority_4647_port_o                )  //o
  );
  Majority majority_4648 (
    .port_i (mixColumns_port_state_out_8_2_0[2:0]), //i
    .port_o (majority_4648_port_o                )  //o
  );
  Majority majority_4649 (
    .port_i (mixColumns_port_state_out_9_2_0[2:0]), //i
    .port_o (majority_4649_port_o                )  //o
  );
  Majority majority_4650 (
    .port_i (mixColumns_port_state_out_10_2_0[2:0]), //i
    .port_o (majority_4650_port_o                 )  //o
  );
  Majority majority_4651 (
    .port_i (mixColumns_port_state_out_11_2_0[2:0]), //i
    .port_o (majority_4651_port_o                 )  //o
  );
  Majority majority_4652 (
    .port_i (mixColumns_port_state_out_12_2_0[2:0]), //i
    .port_o (majority_4652_port_o                 )  //o
  );
  Majority majority_4653 (
    .port_i (mixColumns_port_state_out_13_2_0[2:0]), //i
    .port_o (majority_4653_port_o                 )  //o
  );
  Majority majority_4654 (
    .port_i (mixColumns_port_state_out_14_2_0[2:0]), //i
    .port_o (majority_4654_port_o                 )  //o
  );
  Majority majority_4655 (
    .port_i (mixColumns_port_state_out_15_2_0[2:0]), //i
    .port_o (majority_4655_port_o                 )  //o
  );
  Majority majority_4656 (
    .port_i (mixColumns_port_state_out_0_3_0[2:0]), //i
    .port_o (majority_4656_port_o                )  //o
  );
  Majority majority_4657 (
    .port_i (mixColumns_port_state_out_1_3_0[2:0]), //i
    .port_o (majority_4657_port_o                )  //o
  );
  Majority majority_4658 (
    .port_i (mixColumns_port_state_out_2_3_0[2:0]), //i
    .port_o (majority_4658_port_o                )  //o
  );
  Majority majority_4659 (
    .port_i (mixColumns_port_state_out_3_3_0[2:0]), //i
    .port_o (majority_4659_port_o                )  //o
  );
  Majority majority_4660 (
    .port_i (mixColumns_port_state_out_4_3_0[2:0]), //i
    .port_o (majority_4660_port_o                )  //o
  );
  Majority majority_4661 (
    .port_i (mixColumns_port_state_out_5_3_0[2:0]), //i
    .port_o (majority_4661_port_o                )  //o
  );
  Majority majority_4662 (
    .port_i (mixColumns_port_state_out_6_3_0[2:0]), //i
    .port_o (majority_4662_port_o                )  //o
  );
  Majority majority_4663 (
    .port_i (mixColumns_port_state_out_7_3_0[2:0]), //i
    .port_o (majority_4663_port_o                )  //o
  );
  Majority majority_4664 (
    .port_i (mixColumns_port_state_out_8_3_0[2:0]), //i
    .port_o (majority_4664_port_o                )  //o
  );
  Majority majority_4665 (
    .port_i (mixColumns_port_state_out_9_3_0[2:0]), //i
    .port_o (majority_4665_port_o                )  //o
  );
  Majority majority_4666 (
    .port_i (mixColumns_port_state_out_10_3_0[2:0]), //i
    .port_o (majority_4666_port_o                 )  //o
  );
  Majority majority_4667 (
    .port_i (mixColumns_port_state_out_11_3_0[2:0]), //i
    .port_o (majority_4667_port_o                 )  //o
  );
  Majority majority_4668 (
    .port_i (mixColumns_port_state_out_12_3_0[2:0]), //i
    .port_o (majority_4668_port_o                 )  //o
  );
  Majority majority_4669 (
    .port_i (mixColumns_port_state_out_13_3_0[2:0]), //i
    .port_o (majority_4669_port_o                 )  //o
  );
  Majority majority_4670 (
    .port_i (mixColumns_port_state_out_14_3_0[2:0]), //i
    .port_o (majority_4670_port_o                 )  //o
  );
  Majority majority_4671 (
    .port_i (mixColumns_port_state_out_15_3_0[2:0]), //i
    .port_o (majority_4671_port_o                 )  //o
  );
  Majority majority_4672 (
    .port_i (mixColumns_port_state_out_0_0_1[2:0]), //i
    .port_o (majority_4672_port_o                )  //o
  );
  Majority majority_4673 (
    .port_i (mixColumns_port_state_out_1_0_1[2:0]), //i
    .port_o (majority_4673_port_o                )  //o
  );
  Majority majority_4674 (
    .port_i (mixColumns_port_state_out_2_0_1[2:0]), //i
    .port_o (majority_4674_port_o                )  //o
  );
  Majority majority_4675 (
    .port_i (mixColumns_port_state_out_3_0_1[2:0]), //i
    .port_o (majority_4675_port_o                )  //o
  );
  Majority majority_4676 (
    .port_i (mixColumns_port_state_out_4_0_1[2:0]), //i
    .port_o (majority_4676_port_o                )  //o
  );
  Majority majority_4677 (
    .port_i (mixColumns_port_state_out_5_0_1[2:0]), //i
    .port_o (majority_4677_port_o                )  //o
  );
  Majority majority_4678 (
    .port_i (mixColumns_port_state_out_6_0_1[2:0]), //i
    .port_o (majority_4678_port_o                )  //o
  );
  Majority majority_4679 (
    .port_i (mixColumns_port_state_out_7_0_1[2:0]), //i
    .port_o (majority_4679_port_o                )  //o
  );
  Majority majority_4680 (
    .port_i (mixColumns_port_state_out_8_0_1[2:0]), //i
    .port_o (majority_4680_port_o                )  //o
  );
  Majority majority_4681 (
    .port_i (mixColumns_port_state_out_9_0_1[2:0]), //i
    .port_o (majority_4681_port_o                )  //o
  );
  Majority majority_4682 (
    .port_i (mixColumns_port_state_out_10_0_1[2:0]), //i
    .port_o (majority_4682_port_o                 )  //o
  );
  Majority majority_4683 (
    .port_i (mixColumns_port_state_out_11_0_1[2:0]), //i
    .port_o (majority_4683_port_o                 )  //o
  );
  Majority majority_4684 (
    .port_i (mixColumns_port_state_out_12_0_1[2:0]), //i
    .port_o (majority_4684_port_o                 )  //o
  );
  Majority majority_4685 (
    .port_i (mixColumns_port_state_out_13_0_1[2:0]), //i
    .port_o (majority_4685_port_o                 )  //o
  );
  Majority majority_4686 (
    .port_i (mixColumns_port_state_out_14_0_1[2:0]), //i
    .port_o (majority_4686_port_o                 )  //o
  );
  Majority majority_4687 (
    .port_i (mixColumns_port_state_out_15_0_1[2:0]), //i
    .port_o (majority_4687_port_o                 )  //o
  );
  Majority majority_4688 (
    .port_i (mixColumns_port_state_out_0_1_1[2:0]), //i
    .port_o (majority_4688_port_o                )  //o
  );
  Majority majority_4689 (
    .port_i (mixColumns_port_state_out_1_1_1[2:0]), //i
    .port_o (majority_4689_port_o                )  //o
  );
  Majority majority_4690 (
    .port_i (mixColumns_port_state_out_2_1_1[2:0]), //i
    .port_o (majority_4690_port_o                )  //o
  );
  Majority majority_4691 (
    .port_i (mixColumns_port_state_out_3_1_1[2:0]), //i
    .port_o (majority_4691_port_o                )  //o
  );
  Majority majority_4692 (
    .port_i (mixColumns_port_state_out_4_1_1[2:0]), //i
    .port_o (majority_4692_port_o                )  //o
  );
  Majority majority_4693 (
    .port_i (mixColumns_port_state_out_5_1_1[2:0]), //i
    .port_o (majority_4693_port_o                )  //o
  );
  Majority majority_4694 (
    .port_i (mixColumns_port_state_out_6_1_1[2:0]), //i
    .port_o (majority_4694_port_o                )  //o
  );
  Majority majority_4695 (
    .port_i (mixColumns_port_state_out_7_1_1[2:0]), //i
    .port_o (majority_4695_port_o                )  //o
  );
  Majority majority_4696 (
    .port_i (mixColumns_port_state_out_8_1_1[2:0]), //i
    .port_o (majority_4696_port_o                )  //o
  );
  Majority majority_4697 (
    .port_i (mixColumns_port_state_out_9_1_1[2:0]), //i
    .port_o (majority_4697_port_o                )  //o
  );
  Majority majority_4698 (
    .port_i (mixColumns_port_state_out_10_1_1[2:0]), //i
    .port_o (majority_4698_port_o                 )  //o
  );
  Majority majority_4699 (
    .port_i (mixColumns_port_state_out_11_1_1[2:0]), //i
    .port_o (majority_4699_port_o                 )  //o
  );
  Majority majority_4700 (
    .port_i (mixColumns_port_state_out_12_1_1[2:0]), //i
    .port_o (majority_4700_port_o                 )  //o
  );
  Majority majority_4701 (
    .port_i (mixColumns_port_state_out_13_1_1[2:0]), //i
    .port_o (majority_4701_port_o                 )  //o
  );
  Majority majority_4702 (
    .port_i (mixColumns_port_state_out_14_1_1[2:0]), //i
    .port_o (majority_4702_port_o                 )  //o
  );
  Majority majority_4703 (
    .port_i (mixColumns_port_state_out_15_1_1[2:0]), //i
    .port_o (majority_4703_port_o                 )  //o
  );
  Majority majority_4704 (
    .port_i (mixColumns_port_state_out_0_2_1[2:0]), //i
    .port_o (majority_4704_port_o                )  //o
  );
  Majority majority_4705 (
    .port_i (mixColumns_port_state_out_1_2_1[2:0]), //i
    .port_o (majority_4705_port_o                )  //o
  );
  Majority majority_4706 (
    .port_i (mixColumns_port_state_out_2_2_1[2:0]), //i
    .port_o (majority_4706_port_o                )  //o
  );
  Majority majority_4707 (
    .port_i (mixColumns_port_state_out_3_2_1[2:0]), //i
    .port_o (majority_4707_port_o                )  //o
  );
  Majority majority_4708 (
    .port_i (mixColumns_port_state_out_4_2_1[2:0]), //i
    .port_o (majority_4708_port_o                )  //o
  );
  Majority majority_4709 (
    .port_i (mixColumns_port_state_out_5_2_1[2:0]), //i
    .port_o (majority_4709_port_o                )  //o
  );
  Majority majority_4710 (
    .port_i (mixColumns_port_state_out_6_2_1[2:0]), //i
    .port_o (majority_4710_port_o                )  //o
  );
  Majority majority_4711 (
    .port_i (mixColumns_port_state_out_7_2_1[2:0]), //i
    .port_o (majority_4711_port_o                )  //o
  );
  Majority majority_4712 (
    .port_i (mixColumns_port_state_out_8_2_1[2:0]), //i
    .port_o (majority_4712_port_o                )  //o
  );
  Majority majority_4713 (
    .port_i (mixColumns_port_state_out_9_2_1[2:0]), //i
    .port_o (majority_4713_port_o                )  //o
  );
  Majority majority_4714 (
    .port_i (mixColumns_port_state_out_10_2_1[2:0]), //i
    .port_o (majority_4714_port_o                 )  //o
  );
  Majority majority_4715 (
    .port_i (mixColumns_port_state_out_11_2_1[2:0]), //i
    .port_o (majority_4715_port_o                 )  //o
  );
  Majority majority_4716 (
    .port_i (mixColumns_port_state_out_12_2_1[2:0]), //i
    .port_o (majority_4716_port_o                 )  //o
  );
  Majority majority_4717 (
    .port_i (mixColumns_port_state_out_13_2_1[2:0]), //i
    .port_o (majority_4717_port_o                 )  //o
  );
  Majority majority_4718 (
    .port_i (mixColumns_port_state_out_14_2_1[2:0]), //i
    .port_o (majority_4718_port_o                 )  //o
  );
  Majority majority_4719 (
    .port_i (mixColumns_port_state_out_15_2_1[2:0]), //i
    .port_o (majority_4719_port_o                 )  //o
  );
  Majority majority_4720 (
    .port_i (mixColumns_port_state_out_0_3_1[2:0]), //i
    .port_o (majority_4720_port_o                )  //o
  );
  Majority majority_4721 (
    .port_i (mixColumns_port_state_out_1_3_1[2:0]), //i
    .port_o (majority_4721_port_o                )  //o
  );
  Majority majority_4722 (
    .port_i (mixColumns_port_state_out_2_3_1[2:0]), //i
    .port_o (majority_4722_port_o                )  //o
  );
  Majority majority_4723 (
    .port_i (mixColumns_port_state_out_3_3_1[2:0]), //i
    .port_o (majority_4723_port_o                )  //o
  );
  Majority majority_4724 (
    .port_i (mixColumns_port_state_out_4_3_1[2:0]), //i
    .port_o (majority_4724_port_o                )  //o
  );
  Majority majority_4725 (
    .port_i (mixColumns_port_state_out_5_3_1[2:0]), //i
    .port_o (majority_4725_port_o                )  //o
  );
  Majority majority_4726 (
    .port_i (mixColumns_port_state_out_6_3_1[2:0]), //i
    .port_o (majority_4726_port_o                )  //o
  );
  Majority majority_4727 (
    .port_i (mixColumns_port_state_out_7_3_1[2:0]), //i
    .port_o (majority_4727_port_o                )  //o
  );
  Majority majority_4728 (
    .port_i (mixColumns_port_state_out_8_3_1[2:0]), //i
    .port_o (majority_4728_port_o                )  //o
  );
  Majority majority_4729 (
    .port_i (mixColumns_port_state_out_9_3_1[2:0]), //i
    .port_o (majority_4729_port_o                )  //o
  );
  Majority majority_4730 (
    .port_i (mixColumns_port_state_out_10_3_1[2:0]), //i
    .port_o (majority_4730_port_o                 )  //o
  );
  Majority majority_4731 (
    .port_i (mixColumns_port_state_out_11_3_1[2:0]), //i
    .port_o (majority_4731_port_o                 )  //o
  );
  Majority majority_4732 (
    .port_i (mixColumns_port_state_out_12_3_1[2:0]), //i
    .port_o (majority_4732_port_o                 )  //o
  );
  Majority majority_4733 (
    .port_i (mixColumns_port_state_out_13_3_1[2:0]), //i
    .port_o (majority_4733_port_o                 )  //o
  );
  Majority majority_4734 (
    .port_i (mixColumns_port_state_out_14_3_1[2:0]), //i
    .port_o (majority_4734_port_o                 )  //o
  );
  Majority majority_4735 (
    .port_i (mixColumns_port_state_out_15_3_1[2:0]), //i
    .port_o (majority_4735_port_o                 )  //o
  );
  Majority majority_4736 (
    .port_i (mixColumns_port_state_out_0_0_2[2:0]), //i
    .port_o (majority_4736_port_o                )  //o
  );
  Majority majority_4737 (
    .port_i (mixColumns_port_state_out_1_0_2[2:0]), //i
    .port_o (majority_4737_port_o                )  //o
  );
  Majority majority_4738 (
    .port_i (mixColumns_port_state_out_2_0_2[2:0]), //i
    .port_o (majority_4738_port_o                )  //o
  );
  Majority majority_4739 (
    .port_i (mixColumns_port_state_out_3_0_2[2:0]), //i
    .port_o (majority_4739_port_o                )  //o
  );
  Majority majority_4740 (
    .port_i (mixColumns_port_state_out_4_0_2[2:0]), //i
    .port_o (majority_4740_port_o                )  //o
  );
  Majority majority_4741 (
    .port_i (mixColumns_port_state_out_5_0_2[2:0]), //i
    .port_o (majority_4741_port_o                )  //o
  );
  Majority majority_4742 (
    .port_i (mixColumns_port_state_out_6_0_2[2:0]), //i
    .port_o (majority_4742_port_o                )  //o
  );
  Majority majority_4743 (
    .port_i (mixColumns_port_state_out_7_0_2[2:0]), //i
    .port_o (majority_4743_port_o                )  //o
  );
  Majority majority_4744 (
    .port_i (mixColumns_port_state_out_8_0_2[2:0]), //i
    .port_o (majority_4744_port_o                )  //o
  );
  Majority majority_4745 (
    .port_i (mixColumns_port_state_out_9_0_2[2:0]), //i
    .port_o (majority_4745_port_o                )  //o
  );
  Majority majority_4746 (
    .port_i (mixColumns_port_state_out_10_0_2[2:0]), //i
    .port_o (majority_4746_port_o                 )  //o
  );
  Majority majority_4747 (
    .port_i (mixColumns_port_state_out_11_0_2[2:0]), //i
    .port_o (majority_4747_port_o                 )  //o
  );
  Majority majority_4748 (
    .port_i (mixColumns_port_state_out_12_0_2[2:0]), //i
    .port_o (majority_4748_port_o                 )  //o
  );
  Majority majority_4749 (
    .port_i (mixColumns_port_state_out_13_0_2[2:0]), //i
    .port_o (majority_4749_port_o                 )  //o
  );
  Majority majority_4750 (
    .port_i (mixColumns_port_state_out_14_0_2[2:0]), //i
    .port_o (majority_4750_port_o                 )  //o
  );
  Majority majority_4751 (
    .port_i (mixColumns_port_state_out_15_0_2[2:0]), //i
    .port_o (majority_4751_port_o                 )  //o
  );
  Majority majority_4752 (
    .port_i (mixColumns_port_state_out_0_1_2[2:0]), //i
    .port_o (majority_4752_port_o                )  //o
  );
  Majority majority_4753 (
    .port_i (mixColumns_port_state_out_1_1_2[2:0]), //i
    .port_o (majority_4753_port_o                )  //o
  );
  Majority majority_4754 (
    .port_i (mixColumns_port_state_out_2_1_2[2:0]), //i
    .port_o (majority_4754_port_o                )  //o
  );
  Majority majority_4755 (
    .port_i (mixColumns_port_state_out_3_1_2[2:0]), //i
    .port_o (majority_4755_port_o                )  //o
  );
  Majority majority_4756 (
    .port_i (mixColumns_port_state_out_4_1_2[2:0]), //i
    .port_o (majority_4756_port_o                )  //o
  );
  Majority majority_4757 (
    .port_i (mixColumns_port_state_out_5_1_2[2:0]), //i
    .port_o (majority_4757_port_o                )  //o
  );
  Majority majority_4758 (
    .port_i (mixColumns_port_state_out_6_1_2[2:0]), //i
    .port_o (majority_4758_port_o                )  //o
  );
  Majority majority_4759 (
    .port_i (mixColumns_port_state_out_7_1_2[2:0]), //i
    .port_o (majority_4759_port_o                )  //o
  );
  Majority majority_4760 (
    .port_i (mixColumns_port_state_out_8_1_2[2:0]), //i
    .port_o (majority_4760_port_o                )  //o
  );
  Majority majority_4761 (
    .port_i (mixColumns_port_state_out_9_1_2[2:0]), //i
    .port_o (majority_4761_port_o                )  //o
  );
  Majority majority_4762 (
    .port_i (mixColumns_port_state_out_10_1_2[2:0]), //i
    .port_o (majority_4762_port_o                 )  //o
  );
  Majority majority_4763 (
    .port_i (mixColumns_port_state_out_11_1_2[2:0]), //i
    .port_o (majority_4763_port_o                 )  //o
  );
  Majority majority_4764 (
    .port_i (mixColumns_port_state_out_12_1_2[2:0]), //i
    .port_o (majority_4764_port_o                 )  //o
  );
  Majority majority_4765 (
    .port_i (mixColumns_port_state_out_13_1_2[2:0]), //i
    .port_o (majority_4765_port_o                 )  //o
  );
  Majority majority_4766 (
    .port_i (mixColumns_port_state_out_14_1_2[2:0]), //i
    .port_o (majority_4766_port_o                 )  //o
  );
  Majority majority_4767 (
    .port_i (mixColumns_port_state_out_15_1_2[2:0]), //i
    .port_o (majority_4767_port_o                 )  //o
  );
  Majority majority_4768 (
    .port_i (mixColumns_port_state_out_0_2_2[2:0]), //i
    .port_o (majority_4768_port_o                )  //o
  );
  Majority majority_4769 (
    .port_i (mixColumns_port_state_out_1_2_2[2:0]), //i
    .port_o (majority_4769_port_o                )  //o
  );
  Majority majority_4770 (
    .port_i (mixColumns_port_state_out_2_2_2[2:0]), //i
    .port_o (majority_4770_port_o                )  //o
  );
  Majority majority_4771 (
    .port_i (mixColumns_port_state_out_3_2_2[2:0]), //i
    .port_o (majority_4771_port_o                )  //o
  );
  Majority majority_4772 (
    .port_i (mixColumns_port_state_out_4_2_2[2:0]), //i
    .port_o (majority_4772_port_o                )  //o
  );
  Majority majority_4773 (
    .port_i (mixColumns_port_state_out_5_2_2[2:0]), //i
    .port_o (majority_4773_port_o                )  //o
  );
  Majority majority_4774 (
    .port_i (mixColumns_port_state_out_6_2_2[2:0]), //i
    .port_o (majority_4774_port_o                )  //o
  );
  Majority majority_4775 (
    .port_i (mixColumns_port_state_out_7_2_2[2:0]), //i
    .port_o (majority_4775_port_o                )  //o
  );
  Majority majority_4776 (
    .port_i (mixColumns_port_state_out_8_2_2[2:0]), //i
    .port_o (majority_4776_port_o                )  //o
  );
  Majority majority_4777 (
    .port_i (mixColumns_port_state_out_9_2_2[2:0]), //i
    .port_o (majority_4777_port_o                )  //o
  );
  Majority majority_4778 (
    .port_i (mixColumns_port_state_out_10_2_2[2:0]), //i
    .port_o (majority_4778_port_o                 )  //o
  );
  Majority majority_4779 (
    .port_i (mixColumns_port_state_out_11_2_2[2:0]), //i
    .port_o (majority_4779_port_o                 )  //o
  );
  Majority majority_4780 (
    .port_i (mixColumns_port_state_out_12_2_2[2:0]), //i
    .port_o (majority_4780_port_o                 )  //o
  );
  Majority majority_4781 (
    .port_i (mixColumns_port_state_out_13_2_2[2:0]), //i
    .port_o (majority_4781_port_o                 )  //o
  );
  Majority majority_4782 (
    .port_i (mixColumns_port_state_out_14_2_2[2:0]), //i
    .port_o (majority_4782_port_o                 )  //o
  );
  Majority majority_4783 (
    .port_i (mixColumns_port_state_out_15_2_2[2:0]), //i
    .port_o (majority_4783_port_o                 )  //o
  );
  Majority majority_4784 (
    .port_i (mixColumns_port_state_out_0_3_2[2:0]), //i
    .port_o (majority_4784_port_o                )  //o
  );
  Majority majority_4785 (
    .port_i (mixColumns_port_state_out_1_3_2[2:0]), //i
    .port_o (majority_4785_port_o                )  //o
  );
  Majority majority_4786 (
    .port_i (mixColumns_port_state_out_2_3_2[2:0]), //i
    .port_o (majority_4786_port_o                )  //o
  );
  Majority majority_4787 (
    .port_i (mixColumns_port_state_out_3_3_2[2:0]), //i
    .port_o (majority_4787_port_o                )  //o
  );
  Majority majority_4788 (
    .port_i (mixColumns_port_state_out_4_3_2[2:0]), //i
    .port_o (majority_4788_port_o                )  //o
  );
  Majority majority_4789 (
    .port_i (mixColumns_port_state_out_5_3_2[2:0]), //i
    .port_o (majority_4789_port_o                )  //o
  );
  Majority majority_4790 (
    .port_i (mixColumns_port_state_out_6_3_2[2:0]), //i
    .port_o (majority_4790_port_o                )  //o
  );
  Majority majority_4791 (
    .port_i (mixColumns_port_state_out_7_3_2[2:0]), //i
    .port_o (majority_4791_port_o                )  //o
  );
  Majority majority_4792 (
    .port_i (mixColumns_port_state_out_8_3_2[2:0]), //i
    .port_o (majority_4792_port_o                )  //o
  );
  Majority majority_4793 (
    .port_i (mixColumns_port_state_out_9_3_2[2:0]), //i
    .port_o (majority_4793_port_o                )  //o
  );
  Majority majority_4794 (
    .port_i (mixColumns_port_state_out_10_3_2[2:0]), //i
    .port_o (majority_4794_port_o                 )  //o
  );
  Majority majority_4795 (
    .port_i (mixColumns_port_state_out_11_3_2[2:0]), //i
    .port_o (majority_4795_port_o                 )  //o
  );
  Majority majority_4796 (
    .port_i (mixColumns_port_state_out_12_3_2[2:0]), //i
    .port_o (majority_4796_port_o                 )  //o
  );
  Majority majority_4797 (
    .port_i (mixColumns_port_state_out_13_3_2[2:0]), //i
    .port_o (majority_4797_port_o                 )  //o
  );
  Majority majority_4798 (
    .port_i (mixColumns_port_state_out_14_3_2[2:0]), //i
    .port_o (majority_4798_port_o                 )  //o
  );
  Majority majority_4799 (
    .port_i (mixColumns_port_state_out_15_3_2[2:0]), //i
    .port_o (majority_4799_port_o                 )  //o
  );
  Majority majority_4800 (
    .port_i (mixColumns_port_state_out_0_0_3[2:0]), //i
    .port_o (majority_4800_port_o                )  //o
  );
  Majority majority_4801 (
    .port_i (mixColumns_port_state_out_1_0_3[2:0]), //i
    .port_o (majority_4801_port_o                )  //o
  );
  Majority majority_4802 (
    .port_i (mixColumns_port_state_out_2_0_3[2:0]), //i
    .port_o (majority_4802_port_o                )  //o
  );
  Majority majority_4803 (
    .port_i (mixColumns_port_state_out_3_0_3[2:0]), //i
    .port_o (majority_4803_port_o                )  //o
  );
  Majority majority_4804 (
    .port_i (mixColumns_port_state_out_4_0_3[2:0]), //i
    .port_o (majority_4804_port_o                )  //o
  );
  Majority majority_4805 (
    .port_i (mixColumns_port_state_out_5_0_3[2:0]), //i
    .port_o (majority_4805_port_o                )  //o
  );
  Majority majority_4806 (
    .port_i (mixColumns_port_state_out_6_0_3[2:0]), //i
    .port_o (majority_4806_port_o                )  //o
  );
  Majority majority_4807 (
    .port_i (mixColumns_port_state_out_7_0_3[2:0]), //i
    .port_o (majority_4807_port_o                )  //o
  );
  Majority majority_4808 (
    .port_i (mixColumns_port_state_out_8_0_3[2:0]), //i
    .port_o (majority_4808_port_o                )  //o
  );
  Majority majority_4809 (
    .port_i (mixColumns_port_state_out_9_0_3[2:0]), //i
    .port_o (majority_4809_port_o                )  //o
  );
  Majority majority_4810 (
    .port_i (mixColumns_port_state_out_10_0_3[2:0]), //i
    .port_o (majority_4810_port_o                 )  //o
  );
  Majority majority_4811 (
    .port_i (mixColumns_port_state_out_11_0_3[2:0]), //i
    .port_o (majority_4811_port_o                 )  //o
  );
  Majority majority_4812 (
    .port_i (mixColumns_port_state_out_12_0_3[2:0]), //i
    .port_o (majority_4812_port_o                 )  //o
  );
  Majority majority_4813 (
    .port_i (mixColumns_port_state_out_13_0_3[2:0]), //i
    .port_o (majority_4813_port_o                 )  //o
  );
  Majority majority_4814 (
    .port_i (mixColumns_port_state_out_14_0_3[2:0]), //i
    .port_o (majority_4814_port_o                 )  //o
  );
  Majority majority_4815 (
    .port_i (mixColumns_port_state_out_15_0_3[2:0]), //i
    .port_o (majority_4815_port_o                 )  //o
  );
  Majority majority_4816 (
    .port_i (mixColumns_port_state_out_0_1_3[2:0]), //i
    .port_o (majority_4816_port_o                )  //o
  );
  Majority majority_4817 (
    .port_i (mixColumns_port_state_out_1_1_3[2:0]), //i
    .port_o (majority_4817_port_o                )  //o
  );
  Majority majority_4818 (
    .port_i (mixColumns_port_state_out_2_1_3[2:0]), //i
    .port_o (majority_4818_port_o                )  //o
  );
  Majority majority_4819 (
    .port_i (mixColumns_port_state_out_3_1_3[2:0]), //i
    .port_o (majority_4819_port_o                )  //o
  );
  Majority majority_4820 (
    .port_i (mixColumns_port_state_out_4_1_3[2:0]), //i
    .port_o (majority_4820_port_o                )  //o
  );
  Majority majority_4821 (
    .port_i (mixColumns_port_state_out_5_1_3[2:0]), //i
    .port_o (majority_4821_port_o                )  //o
  );
  Majority majority_4822 (
    .port_i (mixColumns_port_state_out_6_1_3[2:0]), //i
    .port_o (majority_4822_port_o                )  //o
  );
  Majority majority_4823 (
    .port_i (mixColumns_port_state_out_7_1_3[2:0]), //i
    .port_o (majority_4823_port_o                )  //o
  );
  Majority majority_4824 (
    .port_i (mixColumns_port_state_out_8_1_3[2:0]), //i
    .port_o (majority_4824_port_o                )  //o
  );
  Majority majority_4825 (
    .port_i (mixColumns_port_state_out_9_1_3[2:0]), //i
    .port_o (majority_4825_port_o                )  //o
  );
  Majority majority_4826 (
    .port_i (mixColumns_port_state_out_10_1_3[2:0]), //i
    .port_o (majority_4826_port_o                 )  //o
  );
  Majority majority_4827 (
    .port_i (mixColumns_port_state_out_11_1_3[2:0]), //i
    .port_o (majority_4827_port_o                 )  //o
  );
  Majority majority_4828 (
    .port_i (mixColumns_port_state_out_12_1_3[2:0]), //i
    .port_o (majority_4828_port_o                 )  //o
  );
  Majority majority_4829 (
    .port_i (mixColumns_port_state_out_13_1_3[2:0]), //i
    .port_o (majority_4829_port_o                 )  //o
  );
  Majority majority_4830 (
    .port_i (mixColumns_port_state_out_14_1_3[2:0]), //i
    .port_o (majority_4830_port_o                 )  //o
  );
  Majority majority_4831 (
    .port_i (mixColumns_port_state_out_15_1_3[2:0]), //i
    .port_o (majority_4831_port_o                 )  //o
  );
  Majority majority_4832 (
    .port_i (mixColumns_port_state_out_0_2_3[2:0]), //i
    .port_o (majority_4832_port_o                )  //o
  );
  Majority majority_4833 (
    .port_i (mixColumns_port_state_out_1_2_3[2:0]), //i
    .port_o (majority_4833_port_o                )  //o
  );
  Majority majority_4834 (
    .port_i (mixColumns_port_state_out_2_2_3[2:0]), //i
    .port_o (majority_4834_port_o                )  //o
  );
  Majority majority_4835 (
    .port_i (mixColumns_port_state_out_3_2_3[2:0]), //i
    .port_o (majority_4835_port_o                )  //o
  );
  Majority majority_4836 (
    .port_i (mixColumns_port_state_out_4_2_3[2:0]), //i
    .port_o (majority_4836_port_o                )  //o
  );
  Majority majority_4837 (
    .port_i (mixColumns_port_state_out_5_2_3[2:0]), //i
    .port_o (majority_4837_port_o                )  //o
  );
  Majority majority_4838 (
    .port_i (mixColumns_port_state_out_6_2_3[2:0]), //i
    .port_o (majority_4838_port_o                )  //o
  );
  Majority majority_4839 (
    .port_i (mixColumns_port_state_out_7_2_3[2:0]), //i
    .port_o (majority_4839_port_o                )  //o
  );
  Majority majority_4840 (
    .port_i (mixColumns_port_state_out_8_2_3[2:0]), //i
    .port_o (majority_4840_port_o                )  //o
  );
  Majority majority_4841 (
    .port_i (mixColumns_port_state_out_9_2_3[2:0]), //i
    .port_o (majority_4841_port_o                )  //o
  );
  Majority majority_4842 (
    .port_i (mixColumns_port_state_out_10_2_3[2:0]), //i
    .port_o (majority_4842_port_o                 )  //o
  );
  Majority majority_4843 (
    .port_i (mixColumns_port_state_out_11_2_3[2:0]), //i
    .port_o (majority_4843_port_o                 )  //o
  );
  Majority majority_4844 (
    .port_i (mixColumns_port_state_out_12_2_3[2:0]), //i
    .port_o (majority_4844_port_o                 )  //o
  );
  Majority majority_4845 (
    .port_i (mixColumns_port_state_out_13_2_3[2:0]), //i
    .port_o (majority_4845_port_o                 )  //o
  );
  Majority majority_4846 (
    .port_i (mixColumns_port_state_out_14_2_3[2:0]), //i
    .port_o (majority_4846_port_o                 )  //o
  );
  Majority majority_4847 (
    .port_i (mixColumns_port_state_out_15_2_3[2:0]), //i
    .port_o (majority_4847_port_o                 )  //o
  );
  Majority majority_4848 (
    .port_i (mixColumns_port_state_out_0_3_3[2:0]), //i
    .port_o (majority_4848_port_o                )  //o
  );
  Majority majority_4849 (
    .port_i (mixColumns_port_state_out_1_3_3[2:0]), //i
    .port_o (majority_4849_port_o                )  //o
  );
  Majority majority_4850 (
    .port_i (mixColumns_port_state_out_2_3_3[2:0]), //i
    .port_o (majority_4850_port_o                )  //o
  );
  Majority majority_4851 (
    .port_i (mixColumns_port_state_out_3_3_3[2:0]), //i
    .port_o (majority_4851_port_o                )  //o
  );
  Majority majority_4852 (
    .port_i (mixColumns_port_state_out_4_3_3[2:0]), //i
    .port_o (majority_4852_port_o                )  //o
  );
  Majority majority_4853 (
    .port_i (mixColumns_port_state_out_5_3_3[2:0]), //i
    .port_o (majority_4853_port_o                )  //o
  );
  Majority majority_4854 (
    .port_i (mixColumns_port_state_out_6_3_3[2:0]), //i
    .port_o (majority_4854_port_o                )  //o
  );
  Majority majority_4855 (
    .port_i (mixColumns_port_state_out_7_3_3[2:0]), //i
    .port_o (majority_4855_port_o                )  //o
  );
  Majority majority_4856 (
    .port_i (mixColumns_port_state_out_8_3_3[2:0]), //i
    .port_o (majority_4856_port_o                )  //o
  );
  Majority majority_4857 (
    .port_i (mixColumns_port_state_out_9_3_3[2:0]), //i
    .port_o (majority_4857_port_o                )  //o
  );
  Majority majority_4858 (
    .port_i (mixColumns_port_state_out_10_3_3[2:0]), //i
    .port_o (majority_4858_port_o                 )  //o
  );
  Majority majority_4859 (
    .port_i (mixColumns_port_state_out_11_3_3[2:0]), //i
    .port_o (majority_4859_port_o                 )  //o
  );
  Majority majority_4860 (
    .port_i (mixColumns_port_state_out_12_3_3[2:0]), //i
    .port_o (majority_4860_port_o                 )  //o
  );
  Majority majority_4861 (
    .port_i (mixColumns_port_state_out_13_3_3[2:0]), //i
    .port_o (majority_4861_port_o                 )  //o
  );
  Majority majority_4862 (
    .port_i (mixColumns_port_state_out_14_3_3[2:0]), //i
    .port_o (majority_4862_port_o                 )  //o
  );
  Majority majority_4863 (
    .port_i (mixColumns_port_state_out_15_3_3[2:0]), //i
    .port_o (majority_4863_port_o                 )  //o
  );
  Majority majority_4864 (
    .port_i (mixColumns_port_state_out_0_0_4[2:0]), //i
    .port_o (majority_4864_port_o                )  //o
  );
  Majority majority_4865 (
    .port_i (mixColumns_port_state_out_1_0_4[2:0]), //i
    .port_o (majority_4865_port_o                )  //o
  );
  Majority majority_4866 (
    .port_i (mixColumns_port_state_out_2_0_4[2:0]), //i
    .port_o (majority_4866_port_o                )  //o
  );
  Majority majority_4867 (
    .port_i (mixColumns_port_state_out_3_0_4[2:0]), //i
    .port_o (majority_4867_port_o                )  //o
  );
  Majority majority_4868 (
    .port_i (mixColumns_port_state_out_4_0_4[2:0]), //i
    .port_o (majority_4868_port_o                )  //o
  );
  Majority majority_4869 (
    .port_i (mixColumns_port_state_out_5_0_4[2:0]), //i
    .port_o (majority_4869_port_o                )  //o
  );
  Majority majority_4870 (
    .port_i (mixColumns_port_state_out_6_0_4[2:0]), //i
    .port_o (majority_4870_port_o                )  //o
  );
  Majority majority_4871 (
    .port_i (mixColumns_port_state_out_7_0_4[2:0]), //i
    .port_o (majority_4871_port_o                )  //o
  );
  Majority majority_4872 (
    .port_i (mixColumns_port_state_out_8_0_4[2:0]), //i
    .port_o (majority_4872_port_o                )  //o
  );
  Majority majority_4873 (
    .port_i (mixColumns_port_state_out_9_0_4[2:0]), //i
    .port_o (majority_4873_port_o                )  //o
  );
  Majority majority_4874 (
    .port_i (mixColumns_port_state_out_10_0_4[2:0]), //i
    .port_o (majority_4874_port_o                 )  //o
  );
  Majority majority_4875 (
    .port_i (mixColumns_port_state_out_11_0_4[2:0]), //i
    .port_o (majority_4875_port_o                 )  //o
  );
  Majority majority_4876 (
    .port_i (mixColumns_port_state_out_12_0_4[2:0]), //i
    .port_o (majority_4876_port_o                 )  //o
  );
  Majority majority_4877 (
    .port_i (mixColumns_port_state_out_13_0_4[2:0]), //i
    .port_o (majority_4877_port_o                 )  //o
  );
  Majority majority_4878 (
    .port_i (mixColumns_port_state_out_14_0_4[2:0]), //i
    .port_o (majority_4878_port_o                 )  //o
  );
  Majority majority_4879 (
    .port_i (mixColumns_port_state_out_15_0_4[2:0]), //i
    .port_o (majority_4879_port_o                 )  //o
  );
  Majority majority_4880 (
    .port_i (mixColumns_port_state_out_0_1_4[2:0]), //i
    .port_o (majority_4880_port_o                )  //o
  );
  Majority majority_4881 (
    .port_i (mixColumns_port_state_out_1_1_4[2:0]), //i
    .port_o (majority_4881_port_o                )  //o
  );
  Majority majority_4882 (
    .port_i (mixColumns_port_state_out_2_1_4[2:0]), //i
    .port_o (majority_4882_port_o                )  //o
  );
  Majority majority_4883 (
    .port_i (mixColumns_port_state_out_3_1_4[2:0]), //i
    .port_o (majority_4883_port_o                )  //o
  );
  Majority majority_4884 (
    .port_i (mixColumns_port_state_out_4_1_4[2:0]), //i
    .port_o (majority_4884_port_o                )  //o
  );
  Majority majority_4885 (
    .port_i (mixColumns_port_state_out_5_1_4[2:0]), //i
    .port_o (majority_4885_port_o                )  //o
  );
  Majority majority_4886 (
    .port_i (mixColumns_port_state_out_6_1_4[2:0]), //i
    .port_o (majority_4886_port_o                )  //o
  );
  Majority majority_4887 (
    .port_i (mixColumns_port_state_out_7_1_4[2:0]), //i
    .port_o (majority_4887_port_o                )  //o
  );
  Majority majority_4888 (
    .port_i (mixColumns_port_state_out_8_1_4[2:0]), //i
    .port_o (majority_4888_port_o                )  //o
  );
  Majority majority_4889 (
    .port_i (mixColumns_port_state_out_9_1_4[2:0]), //i
    .port_o (majority_4889_port_o                )  //o
  );
  Majority majority_4890 (
    .port_i (mixColumns_port_state_out_10_1_4[2:0]), //i
    .port_o (majority_4890_port_o                 )  //o
  );
  Majority majority_4891 (
    .port_i (mixColumns_port_state_out_11_1_4[2:0]), //i
    .port_o (majority_4891_port_o                 )  //o
  );
  Majority majority_4892 (
    .port_i (mixColumns_port_state_out_12_1_4[2:0]), //i
    .port_o (majority_4892_port_o                 )  //o
  );
  Majority majority_4893 (
    .port_i (mixColumns_port_state_out_13_1_4[2:0]), //i
    .port_o (majority_4893_port_o                 )  //o
  );
  Majority majority_4894 (
    .port_i (mixColumns_port_state_out_14_1_4[2:0]), //i
    .port_o (majority_4894_port_o                 )  //o
  );
  Majority majority_4895 (
    .port_i (mixColumns_port_state_out_15_1_4[2:0]), //i
    .port_o (majority_4895_port_o                 )  //o
  );
  Majority majority_4896 (
    .port_i (mixColumns_port_state_out_0_2_4[2:0]), //i
    .port_o (majority_4896_port_o                )  //o
  );
  Majority majority_4897 (
    .port_i (mixColumns_port_state_out_1_2_4[2:0]), //i
    .port_o (majority_4897_port_o                )  //o
  );
  Majority majority_4898 (
    .port_i (mixColumns_port_state_out_2_2_4[2:0]), //i
    .port_o (majority_4898_port_o                )  //o
  );
  Majority majority_4899 (
    .port_i (mixColumns_port_state_out_3_2_4[2:0]), //i
    .port_o (majority_4899_port_o                )  //o
  );
  Majority majority_4900 (
    .port_i (mixColumns_port_state_out_4_2_4[2:0]), //i
    .port_o (majority_4900_port_o                )  //o
  );
  Majority majority_4901 (
    .port_i (mixColumns_port_state_out_5_2_4[2:0]), //i
    .port_o (majority_4901_port_o                )  //o
  );
  Majority majority_4902 (
    .port_i (mixColumns_port_state_out_6_2_4[2:0]), //i
    .port_o (majority_4902_port_o                )  //o
  );
  Majority majority_4903 (
    .port_i (mixColumns_port_state_out_7_2_4[2:0]), //i
    .port_o (majority_4903_port_o                )  //o
  );
  Majority majority_4904 (
    .port_i (mixColumns_port_state_out_8_2_4[2:0]), //i
    .port_o (majority_4904_port_o                )  //o
  );
  Majority majority_4905 (
    .port_i (mixColumns_port_state_out_9_2_4[2:0]), //i
    .port_o (majority_4905_port_o                )  //o
  );
  Majority majority_4906 (
    .port_i (mixColumns_port_state_out_10_2_4[2:0]), //i
    .port_o (majority_4906_port_o                 )  //o
  );
  Majority majority_4907 (
    .port_i (mixColumns_port_state_out_11_2_4[2:0]), //i
    .port_o (majority_4907_port_o                 )  //o
  );
  Majority majority_4908 (
    .port_i (mixColumns_port_state_out_12_2_4[2:0]), //i
    .port_o (majority_4908_port_o                 )  //o
  );
  Majority majority_4909 (
    .port_i (mixColumns_port_state_out_13_2_4[2:0]), //i
    .port_o (majority_4909_port_o                 )  //o
  );
  Majority majority_4910 (
    .port_i (mixColumns_port_state_out_14_2_4[2:0]), //i
    .port_o (majority_4910_port_o                 )  //o
  );
  Majority majority_4911 (
    .port_i (mixColumns_port_state_out_15_2_4[2:0]), //i
    .port_o (majority_4911_port_o                 )  //o
  );
  Majority majority_4912 (
    .port_i (mixColumns_port_state_out_0_3_4[2:0]), //i
    .port_o (majority_4912_port_o                )  //o
  );
  Majority majority_4913 (
    .port_i (mixColumns_port_state_out_1_3_4[2:0]), //i
    .port_o (majority_4913_port_o                )  //o
  );
  Majority majority_4914 (
    .port_i (mixColumns_port_state_out_2_3_4[2:0]), //i
    .port_o (majority_4914_port_o                )  //o
  );
  Majority majority_4915 (
    .port_i (mixColumns_port_state_out_3_3_4[2:0]), //i
    .port_o (majority_4915_port_o                )  //o
  );
  Majority majority_4916 (
    .port_i (mixColumns_port_state_out_4_3_4[2:0]), //i
    .port_o (majority_4916_port_o                )  //o
  );
  Majority majority_4917 (
    .port_i (mixColumns_port_state_out_5_3_4[2:0]), //i
    .port_o (majority_4917_port_o                )  //o
  );
  Majority majority_4918 (
    .port_i (mixColumns_port_state_out_6_3_4[2:0]), //i
    .port_o (majority_4918_port_o                )  //o
  );
  Majority majority_4919 (
    .port_i (mixColumns_port_state_out_7_3_4[2:0]), //i
    .port_o (majority_4919_port_o                )  //o
  );
  Majority majority_4920 (
    .port_i (mixColumns_port_state_out_8_3_4[2:0]), //i
    .port_o (majority_4920_port_o                )  //o
  );
  Majority majority_4921 (
    .port_i (mixColumns_port_state_out_9_3_4[2:0]), //i
    .port_o (majority_4921_port_o                )  //o
  );
  Majority majority_4922 (
    .port_i (mixColumns_port_state_out_10_3_4[2:0]), //i
    .port_o (majority_4922_port_o                 )  //o
  );
  Majority majority_4923 (
    .port_i (mixColumns_port_state_out_11_3_4[2:0]), //i
    .port_o (majority_4923_port_o                 )  //o
  );
  Majority majority_4924 (
    .port_i (mixColumns_port_state_out_12_3_4[2:0]), //i
    .port_o (majority_4924_port_o                 )  //o
  );
  Majority majority_4925 (
    .port_i (mixColumns_port_state_out_13_3_4[2:0]), //i
    .port_o (majority_4925_port_o                 )  //o
  );
  Majority majority_4926 (
    .port_i (mixColumns_port_state_out_14_3_4[2:0]), //i
    .port_o (majority_4926_port_o                 )  //o
  );
  Majority majority_4927 (
    .port_i (mixColumns_port_state_out_15_3_4[2:0]), //i
    .port_o (majority_4927_port_o                 )  //o
  );
  Majority majority_4928 (
    .port_i (mixColumns_port_state_out_0_0_5[2:0]), //i
    .port_o (majority_4928_port_o                )  //o
  );
  Majority majority_4929 (
    .port_i (mixColumns_port_state_out_1_0_5[2:0]), //i
    .port_o (majority_4929_port_o                )  //o
  );
  Majority majority_4930 (
    .port_i (mixColumns_port_state_out_2_0_5[2:0]), //i
    .port_o (majority_4930_port_o                )  //o
  );
  Majority majority_4931 (
    .port_i (mixColumns_port_state_out_3_0_5[2:0]), //i
    .port_o (majority_4931_port_o                )  //o
  );
  Majority majority_4932 (
    .port_i (mixColumns_port_state_out_4_0_5[2:0]), //i
    .port_o (majority_4932_port_o                )  //o
  );
  Majority majority_4933 (
    .port_i (mixColumns_port_state_out_5_0_5[2:0]), //i
    .port_o (majority_4933_port_o                )  //o
  );
  Majority majority_4934 (
    .port_i (mixColumns_port_state_out_6_0_5[2:0]), //i
    .port_o (majority_4934_port_o                )  //o
  );
  Majority majority_4935 (
    .port_i (mixColumns_port_state_out_7_0_5[2:0]), //i
    .port_o (majority_4935_port_o                )  //o
  );
  Majority majority_4936 (
    .port_i (mixColumns_port_state_out_8_0_5[2:0]), //i
    .port_o (majority_4936_port_o                )  //o
  );
  Majority majority_4937 (
    .port_i (mixColumns_port_state_out_9_0_5[2:0]), //i
    .port_o (majority_4937_port_o                )  //o
  );
  Majority majority_4938 (
    .port_i (mixColumns_port_state_out_10_0_5[2:0]), //i
    .port_o (majority_4938_port_o                 )  //o
  );
  Majority majority_4939 (
    .port_i (mixColumns_port_state_out_11_0_5[2:0]), //i
    .port_o (majority_4939_port_o                 )  //o
  );
  Majority majority_4940 (
    .port_i (mixColumns_port_state_out_12_0_5[2:0]), //i
    .port_o (majority_4940_port_o                 )  //o
  );
  Majority majority_4941 (
    .port_i (mixColumns_port_state_out_13_0_5[2:0]), //i
    .port_o (majority_4941_port_o                 )  //o
  );
  Majority majority_4942 (
    .port_i (mixColumns_port_state_out_14_0_5[2:0]), //i
    .port_o (majority_4942_port_o                 )  //o
  );
  Majority majority_4943 (
    .port_i (mixColumns_port_state_out_15_0_5[2:0]), //i
    .port_o (majority_4943_port_o                 )  //o
  );
  Majority majority_4944 (
    .port_i (mixColumns_port_state_out_0_1_5[2:0]), //i
    .port_o (majority_4944_port_o                )  //o
  );
  Majority majority_4945 (
    .port_i (mixColumns_port_state_out_1_1_5[2:0]), //i
    .port_o (majority_4945_port_o                )  //o
  );
  Majority majority_4946 (
    .port_i (mixColumns_port_state_out_2_1_5[2:0]), //i
    .port_o (majority_4946_port_o                )  //o
  );
  Majority majority_4947 (
    .port_i (mixColumns_port_state_out_3_1_5[2:0]), //i
    .port_o (majority_4947_port_o                )  //o
  );
  Majority majority_4948 (
    .port_i (mixColumns_port_state_out_4_1_5[2:0]), //i
    .port_o (majority_4948_port_o                )  //o
  );
  Majority majority_4949 (
    .port_i (mixColumns_port_state_out_5_1_5[2:0]), //i
    .port_o (majority_4949_port_o                )  //o
  );
  Majority majority_4950 (
    .port_i (mixColumns_port_state_out_6_1_5[2:0]), //i
    .port_o (majority_4950_port_o                )  //o
  );
  Majority majority_4951 (
    .port_i (mixColumns_port_state_out_7_1_5[2:0]), //i
    .port_o (majority_4951_port_o                )  //o
  );
  Majority majority_4952 (
    .port_i (mixColumns_port_state_out_8_1_5[2:0]), //i
    .port_o (majority_4952_port_o                )  //o
  );
  Majority majority_4953 (
    .port_i (mixColumns_port_state_out_9_1_5[2:0]), //i
    .port_o (majority_4953_port_o                )  //o
  );
  Majority majority_4954 (
    .port_i (mixColumns_port_state_out_10_1_5[2:0]), //i
    .port_o (majority_4954_port_o                 )  //o
  );
  Majority majority_4955 (
    .port_i (mixColumns_port_state_out_11_1_5[2:0]), //i
    .port_o (majority_4955_port_o                 )  //o
  );
  Majority majority_4956 (
    .port_i (mixColumns_port_state_out_12_1_5[2:0]), //i
    .port_o (majority_4956_port_o                 )  //o
  );
  Majority majority_4957 (
    .port_i (mixColumns_port_state_out_13_1_5[2:0]), //i
    .port_o (majority_4957_port_o                 )  //o
  );
  Majority majority_4958 (
    .port_i (mixColumns_port_state_out_14_1_5[2:0]), //i
    .port_o (majority_4958_port_o                 )  //o
  );
  Majority majority_4959 (
    .port_i (mixColumns_port_state_out_15_1_5[2:0]), //i
    .port_o (majority_4959_port_o                 )  //o
  );
  Majority majority_4960 (
    .port_i (mixColumns_port_state_out_0_2_5[2:0]), //i
    .port_o (majority_4960_port_o                )  //o
  );
  Majority majority_4961 (
    .port_i (mixColumns_port_state_out_1_2_5[2:0]), //i
    .port_o (majority_4961_port_o                )  //o
  );
  Majority majority_4962 (
    .port_i (mixColumns_port_state_out_2_2_5[2:0]), //i
    .port_o (majority_4962_port_o                )  //o
  );
  Majority majority_4963 (
    .port_i (mixColumns_port_state_out_3_2_5[2:0]), //i
    .port_o (majority_4963_port_o                )  //o
  );
  Majority majority_4964 (
    .port_i (mixColumns_port_state_out_4_2_5[2:0]), //i
    .port_o (majority_4964_port_o                )  //o
  );
  Majority majority_4965 (
    .port_i (mixColumns_port_state_out_5_2_5[2:0]), //i
    .port_o (majority_4965_port_o                )  //o
  );
  Majority majority_4966 (
    .port_i (mixColumns_port_state_out_6_2_5[2:0]), //i
    .port_o (majority_4966_port_o                )  //o
  );
  Majority majority_4967 (
    .port_i (mixColumns_port_state_out_7_2_5[2:0]), //i
    .port_o (majority_4967_port_o                )  //o
  );
  Majority majority_4968 (
    .port_i (mixColumns_port_state_out_8_2_5[2:0]), //i
    .port_o (majority_4968_port_o                )  //o
  );
  Majority majority_4969 (
    .port_i (mixColumns_port_state_out_9_2_5[2:0]), //i
    .port_o (majority_4969_port_o                )  //o
  );
  Majority majority_4970 (
    .port_i (mixColumns_port_state_out_10_2_5[2:0]), //i
    .port_o (majority_4970_port_o                 )  //o
  );
  Majority majority_4971 (
    .port_i (mixColumns_port_state_out_11_2_5[2:0]), //i
    .port_o (majority_4971_port_o                 )  //o
  );
  Majority majority_4972 (
    .port_i (mixColumns_port_state_out_12_2_5[2:0]), //i
    .port_o (majority_4972_port_o                 )  //o
  );
  Majority majority_4973 (
    .port_i (mixColumns_port_state_out_13_2_5[2:0]), //i
    .port_o (majority_4973_port_o                 )  //o
  );
  Majority majority_4974 (
    .port_i (mixColumns_port_state_out_14_2_5[2:0]), //i
    .port_o (majority_4974_port_o                 )  //o
  );
  Majority majority_4975 (
    .port_i (mixColumns_port_state_out_15_2_5[2:0]), //i
    .port_o (majority_4975_port_o                 )  //o
  );
  Majority majority_4976 (
    .port_i (mixColumns_port_state_out_0_3_5[2:0]), //i
    .port_o (majority_4976_port_o                )  //o
  );
  Majority majority_4977 (
    .port_i (mixColumns_port_state_out_1_3_5[2:0]), //i
    .port_o (majority_4977_port_o                )  //o
  );
  Majority majority_4978 (
    .port_i (mixColumns_port_state_out_2_3_5[2:0]), //i
    .port_o (majority_4978_port_o                )  //o
  );
  Majority majority_4979 (
    .port_i (mixColumns_port_state_out_3_3_5[2:0]), //i
    .port_o (majority_4979_port_o                )  //o
  );
  Majority majority_4980 (
    .port_i (mixColumns_port_state_out_4_3_5[2:0]), //i
    .port_o (majority_4980_port_o                )  //o
  );
  Majority majority_4981 (
    .port_i (mixColumns_port_state_out_5_3_5[2:0]), //i
    .port_o (majority_4981_port_o                )  //o
  );
  Majority majority_4982 (
    .port_i (mixColumns_port_state_out_6_3_5[2:0]), //i
    .port_o (majority_4982_port_o                )  //o
  );
  Majority majority_4983 (
    .port_i (mixColumns_port_state_out_7_3_5[2:0]), //i
    .port_o (majority_4983_port_o                )  //o
  );
  Majority majority_4984 (
    .port_i (mixColumns_port_state_out_8_3_5[2:0]), //i
    .port_o (majority_4984_port_o                )  //o
  );
  Majority majority_4985 (
    .port_i (mixColumns_port_state_out_9_3_5[2:0]), //i
    .port_o (majority_4985_port_o                )  //o
  );
  Majority majority_4986 (
    .port_i (mixColumns_port_state_out_10_3_5[2:0]), //i
    .port_o (majority_4986_port_o                 )  //o
  );
  Majority majority_4987 (
    .port_i (mixColumns_port_state_out_11_3_5[2:0]), //i
    .port_o (majority_4987_port_o                 )  //o
  );
  Majority majority_4988 (
    .port_i (mixColumns_port_state_out_12_3_5[2:0]), //i
    .port_o (majority_4988_port_o                 )  //o
  );
  Majority majority_4989 (
    .port_i (mixColumns_port_state_out_13_3_5[2:0]), //i
    .port_o (majority_4989_port_o                 )  //o
  );
  Majority majority_4990 (
    .port_i (mixColumns_port_state_out_14_3_5[2:0]), //i
    .port_o (majority_4990_port_o                 )  //o
  );
  Majority majority_4991 (
    .port_i (mixColumns_port_state_out_15_3_5[2:0]), //i
    .port_o (majority_4991_port_o                 )  //o
  );
  Majority majority_4992 (
    .port_i (mixColumns_port_state_out_0_0_6[2:0]), //i
    .port_o (majority_4992_port_o                )  //o
  );
  Majority majority_4993 (
    .port_i (mixColumns_port_state_out_1_0_6[2:0]), //i
    .port_o (majority_4993_port_o                )  //o
  );
  Majority majority_4994 (
    .port_i (mixColumns_port_state_out_2_0_6[2:0]), //i
    .port_o (majority_4994_port_o                )  //o
  );
  Majority majority_4995 (
    .port_i (mixColumns_port_state_out_3_0_6[2:0]), //i
    .port_o (majority_4995_port_o                )  //o
  );
  Majority majority_4996 (
    .port_i (mixColumns_port_state_out_4_0_6[2:0]), //i
    .port_o (majority_4996_port_o                )  //o
  );
  Majority majority_4997 (
    .port_i (mixColumns_port_state_out_5_0_6[2:0]), //i
    .port_o (majority_4997_port_o                )  //o
  );
  Majority majority_4998 (
    .port_i (mixColumns_port_state_out_6_0_6[2:0]), //i
    .port_o (majority_4998_port_o                )  //o
  );
  Majority majority_4999 (
    .port_i (mixColumns_port_state_out_7_0_6[2:0]), //i
    .port_o (majority_4999_port_o                )  //o
  );
  Majority majority_5000 (
    .port_i (mixColumns_port_state_out_8_0_6[2:0]), //i
    .port_o (majority_5000_port_o                )  //o
  );
  Majority majority_5001 (
    .port_i (mixColumns_port_state_out_9_0_6[2:0]), //i
    .port_o (majority_5001_port_o                )  //o
  );
  Majority majority_5002 (
    .port_i (mixColumns_port_state_out_10_0_6[2:0]), //i
    .port_o (majority_5002_port_o                 )  //o
  );
  Majority majority_5003 (
    .port_i (mixColumns_port_state_out_11_0_6[2:0]), //i
    .port_o (majority_5003_port_o                 )  //o
  );
  Majority majority_5004 (
    .port_i (mixColumns_port_state_out_12_0_6[2:0]), //i
    .port_o (majority_5004_port_o                 )  //o
  );
  Majority majority_5005 (
    .port_i (mixColumns_port_state_out_13_0_6[2:0]), //i
    .port_o (majority_5005_port_o                 )  //o
  );
  Majority majority_5006 (
    .port_i (mixColumns_port_state_out_14_0_6[2:0]), //i
    .port_o (majority_5006_port_o                 )  //o
  );
  Majority majority_5007 (
    .port_i (mixColumns_port_state_out_15_0_6[2:0]), //i
    .port_o (majority_5007_port_o                 )  //o
  );
  Majority majority_5008 (
    .port_i (mixColumns_port_state_out_0_1_6[2:0]), //i
    .port_o (majority_5008_port_o                )  //o
  );
  Majority majority_5009 (
    .port_i (mixColumns_port_state_out_1_1_6[2:0]), //i
    .port_o (majority_5009_port_o                )  //o
  );
  Majority majority_5010 (
    .port_i (mixColumns_port_state_out_2_1_6[2:0]), //i
    .port_o (majority_5010_port_o                )  //o
  );
  Majority majority_5011 (
    .port_i (mixColumns_port_state_out_3_1_6[2:0]), //i
    .port_o (majority_5011_port_o                )  //o
  );
  Majority majority_5012 (
    .port_i (mixColumns_port_state_out_4_1_6[2:0]), //i
    .port_o (majority_5012_port_o                )  //o
  );
  Majority majority_5013 (
    .port_i (mixColumns_port_state_out_5_1_6[2:0]), //i
    .port_o (majority_5013_port_o                )  //o
  );
  Majority majority_5014 (
    .port_i (mixColumns_port_state_out_6_1_6[2:0]), //i
    .port_o (majority_5014_port_o                )  //o
  );
  Majority majority_5015 (
    .port_i (mixColumns_port_state_out_7_1_6[2:0]), //i
    .port_o (majority_5015_port_o                )  //o
  );
  Majority majority_5016 (
    .port_i (mixColumns_port_state_out_8_1_6[2:0]), //i
    .port_o (majority_5016_port_o                )  //o
  );
  Majority majority_5017 (
    .port_i (mixColumns_port_state_out_9_1_6[2:0]), //i
    .port_o (majority_5017_port_o                )  //o
  );
  Majority majority_5018 (
    .port_i (mixColumns_port_state_out_10_1_6[2:0]), //i
    .port_o (majority_5018_port_o                 )  //o
  );
  Majority majority_5019 (
    .port_i (mixColumns_port_state_out_11_1_6[2:0]), //i
    .port_o (majority_5019_port_o                 )  //o
  );
  Majority majority_5020 (
    .port_i (mixColumns_port_state_out_12_1_6[2:0]), //i
    .port_o (majority_5020_port_o                 )  //o
  );
  Majority majority_5021 (
    .port_i (mixColumns_port_state_out_13_1_6[2:0]), //i
    .port_o (majority_5021_port_o                 )  //o
  );
  Majority majority_5022 (
    .port_i (mixColumns_port_state_out_14_1_6[2:0]), //i
    .port_o (majority_5022_port_o                 )  //o
  );
  Majority majority_5023 (
    .port_i (mixColumns_port_state_out_15_1_6[2:0]), //i
    .port_o (majority_5023_port_o                 )  //o
  );
  Majority majority_5024 (
    .port_i (mixColumns_port_state_out_0_2_6[2:0]), //i
    .port_o (majority_5024_port_o                )  //o
  );
  Majority majority_5025 (
    .port_i (mixColumns_port_state_out_1_2_6[2:0]), //i
    .port_o (majority_5025_port_o                )  //o
  );
  Majority majority_5026 (
    .port_i (mixColumns_port_state_out_2_2_6[2:0]), //i
    .port_o (majority_5026_port_o                )  //o
  );
  Majority majority_5027 (
    .port_i (mixColumns_port_state_out_3_2_6[2:0]), //i
    .port_o (majority_5027_port_o                )  //o
  );
  Majority majority_5028 (
    .port_i (mixColumns_port_state_out_4_2_6[2:0]), //i
    .port_o (majority_5028_port_o                )  //o
  );
  Majority majority_5029 (
    .port_i (mixColumns_port_state_out_5_2_6[2:0]), //i
    .port_o (majority_5029_port_o                )  //o
  );
  Majority majority_5030 (
    .port_i (mixColumns_port_state_out_6_2_6[2:0]), //i
    .port_o (majority_5030_port_o                )  //o
  );
  Majority majority_5031 (
    .port_i (mixColumns_port_state_out_7_2_6[2:0]), //i
    .port_o (majority_5031_port_o                )  //o
  );
  Majority majority_5032 (
    .port_i (mixColumns_port_state_out_8_2_6[2:0]), //i
    .port_o (majority_5032_port_o                )  //o
  );
  Majority majority_5033 (
    .port_i (mixColumns_port_state_out_9_2_6[2:0]), //i
    .port_o (majority_5033_port_o                )  //o
  );
  Majority majority_5034 (
    .port_i (mixColumns_port_state_out_10_2_6[2:0]), //i
    .port_o (majority_5034_port_o                 )  //o
  );
  Majority majority_5035 (
    .port_i (mixColumns_port_state_out_11_2_6[2:0]), //i
    .port_o (majority_5035_port_o                 )  //o
  );
  Majority majority_5036 (
    .port_i (mixColumns_port_state_out_12_2_6[2:0]), //i
    .port_o (majority_5036_port_o                 )  //o
  );
  Majority majority_5037 (
    .port_i (mixColumns_port_state_out_13_2_6[2:0]), //i
    .port_o (majority_5037_port_o                 )  //o
  );
  Majority majority_5038 (
    .port_i (mixColumns_port_state_out_14_2_6[2:0]), //i
    .port_o (majority_5038_port_o                 )  //o
  );
  Majority majority_5039 (
    .port_i (mixColumns_port_state_out_15_2_6[2:0]), //i
    .port_o (majority_5039_port_o                 )  //o
  );
  Majority majority_5040 (
    .port_i (mixColumns_port_state_out_0_3_6[2:0]), //i
    .port_o (majority_5040_port_o                )  //o
  );
  Majority majority_5041 (
    .port_i (mixColumns_port_state_out_1_3_6[2:0]), //i
    .port_o (majority_5041_port_o                )  //o
  );
  Majority majority_5042 (
    .port_i (mixColumns_port_state_out_2_3_6[2:0]), //i
    .port_o (majority_5042_port_o                )  //o
  );
  Majority majority_5043 (
    .port_i (mixColumns_port_state_out_3_3_6[2:0]), //i
    .port_o (majority_5043_port_o                )  //o
  );
  Majority majority_5044 (
    .port_i (mixColumns_port_state_out_4_3_6[2:0]), //i
    .port_o (majority_5044_port_o                )  //o
  );
  Majority majority_5045 (
    .port_i (mixColumns_port_state_out_5_3_6[2:0]), //i
    .port_o (majority_5045_port_o                )  //o
  );
  Majority majority_5046 (
    .port_i (mixColumns_port_state_out_6_3_6[2:0]), //i
    .port_o (majority_5046_port_o                )  //o
  );
  Majority majority_5047 (
    .port_i (mixColumns_port_state_out_7_3_6[2:0]), //i
    .port_o (majority_5047_port_o                )  //o
  );
  Majority majority_5048 (
    .port_i (mixColumns_port_state_out_8_3_6[2:0]), //i
    .port_o (majority_5048_port_o                )  //o
  );
  Majority majority_5049 (
    .port_i (mixColumns_port_state_out_9_3_6[2:0]), //i
    .port_o (majority_5049_port_o                )  //o
  );
  Majority majority_5050 (
    .port_i (mixColumns_port_state_out_10_3_6[2:0]), //i
    .port_o (majority_5050_port_o                 )  //o
  );
  Majority majority_5051 (
    .port_i (mixColumns_port_state_out_11_3_6[2:0]), //i
    .port_o (majority_5051_port_o                 )  //o
  );
  Majority majority_5052 (
    .port_i (mixColumns_port_state_out_12_3_6[2:0]), //i
    .port_o (majority_5052_port_o                 )  //o
  );
  Majority majority_5053 (
    .port_i (mixColumns_port_state_out_13_3_6[2:0]), //i
    .port_o (majority_5053_port_o                 )  //o
  );
  Majority majority_5054 (
    .port_i (mixColumns_port_state_out_14_3_6[2:0]), //i
    .port_o (majority_5054_port_o                 )  //o
  );
  Majority majority_5055 (
    .port_i (mixColumns_port_state_out_15_3_6[2:0]), //i
    .port_o (majority_5055_port_o                 )  //o
  );
  Majority majority_5056 (
    .port_i (mixColumns_port_state_out_0_0_7[2:0]), //i
    .port_o (majority_5056_port_o                )  //o
  );
  Majority majority_5057 (
    .port_i (mixColumns_port_state_out_1_0_7[2:0]), //i
    .port_o (majority_5057_port_o                )  //o
  );
  Majority majority_5058 (
    .port_i (mixColumns_port_state_out_2_0_7[2:0]), //i
    .port_o (majority_5058_port_o                )  //o
  );
  Majority majority_5059 (
    .port_i (mixColumns_port_state_out_3_0_7[2:0]), //i
    .port_o (majority_5059_port_o                )  //o
  );
  Majority majority_5060 (
    .port_i (mixColumns_port_state_out_4_0_7[2:0]), //i
    .port_o (majority_5060_port_o                )  //o
  );
  Majority majority_5061 (
    .port_i (mixColumns_port_state_out_5_0_7[2:0]), //i
    .port_o (majority_5061_port_o                )  //o
  );
  Majority majority_5062 (
    .port_i (mixColumns_port_state_out_6_0_7[2:0]), //i
    .port_o (majority_5062_port_o                )  //o
  );
  Majority majority_5063 (
    .port_i (mixColumns_port_state_out_7_0_7[2:0]), //i
    .port_o (majority_5063_port_o                )  //o
  );
  Majority majority_5064 (
    .port_i (mixColumns_port_state_out_8_0_7[2:0]), //i
    .port_o (majority_5064_port_o                )  //o
  );
  Majority majority_5065 (
    .port_i (mixColumns_port_state_out_9_0_7[2:0]), //i
    .port_o (majority_5065_port_o                )  //o
  );
  Majority majority_5066 (
    .port_i (mixColumns_port_state_out_10_0_7[2:0]), //i
    .port_o (majority_5066_port_o                 )  //o
  );
  Majority majority_5067 (
    .port_i (mixColumns_port_state_out_11_0_7[2:0]), //i
    .port_o (majority_5067_port_o                 )  //o
  );
  Majority majority_5068 (
    .port_i (mixColumns_port_state_out_12_0_7[2:0]), //i
    .port_o (majority_5068_port_o                 )  //o
  );
  Majority majority_5069 (
    .port_i (mixColumns_port_state_out_13_0_7[2:0]), //i
    .port_o (majority_5069_port_o                 )  //o
  );
  Majority majority_5070 (
    .port_i (mixColumns_port_state_out_14_0_7[2:0]), //i
    .port_o (majority_5070_port_o                 )  //o
  );
  Majority majority_5071 (
    .port_i (mixColumns_port_state_out_15_0_7[2:0]), //i
    .port_o (majority_5071_port_o                 )  //o
  );
  Majority majority_5072 (
    .port_i (mixColumns_port_state_out_0_1_7[2:0]), //i
    .port_o (majority_5072_port_o                )  //o
  );
  Majority majority_5073 (
    .port_i (mixColumns_port_state_out_1_1_7[2:0]), //i
    .port_o (majority_5073_port_o                )  //o
  );
  Majority majority_5074 (
    .port_i (mixColumns_port_state_out_2_1_7[2:0]), //i
    .port_o (majority_5074_port_o                )  //o
  );
  Majority majority_5075 (
    .port_i (mixColumns_port_state_out_3_1_7[2:0]), //i
    .port_o (majority_5075_port_o                )  //o
  );
  Majority majority_5076 (
    .port_i (mixColumns_port_state_out_4_1_7[2:0]), //i
    .port_o (majority_5076_port_o                )  //o
  );
  Majority majority_5077 (
    .port_i (mixColumns_port_state_out_5_1_7[2:0]), //i
    .port_o (majority_5077_port_o                )  //o
  );
  Majority majority_5078 (
    .port_i (mixColumns_port_state_out_6_1_7[2:0]), //i
    .port_o (majority_5078_port_o                )  //o
  );
  Majority majority_5079 (
    .port_i (mixColumns_port_state_out_7_1_7[2:0]), //i
    .port_o (majority_5079_port_o                )  //o
  );
  Majority majority_5080 (
    .port_i (mixColumns_port_state_out_8_1_7[2:0]), //i
    .port_o (majority_5080_port_o                )  //o
  );
  Majority majority_5081 (
    .port_i (mixColumns_port_state_out_9_1_7[2:0]), //i
    .port_o (majority_5081_port_o                )  //o
  );
  Majority majority_5082 (
    .port_i (mixColumns_port_state_out_10_1_7[2:0]), //i
    .port_o (majority_5082_port_o                 )  //o
  );
  Majority majority_5083 (
    .port_i (mixColumns_port_state_out_11_1_7[2:0]), //i
    .port_o (majority_5083_port_o                 )  //o
  );
  Majority majority_5084 (
    .port_i (mixColumns_port_state_out_12_1_7[2:0]), //i
    .port_o (majority_5084_port_o                 )  //o
  );
  Majority majority_5085 (
    .port_i (mixColumns_port_state_out_13_1_7[2:0]), //i
    .port_o (majority_5085_port_o                 )  //o
  );
  Majority majority_5086 (
    .port_i (mixColumns_port_state_out_14_1_7[2:0]), //i
    .port_o (majority_5086_port_o                 )  //o
  );
  Majority majority_5087 (
    .port_i (mixColumns_port_state_out_15_1_7[2:0]), //i
    .port_o (majority_5087_port_o                 )  //o
  );
  Majority majority_5088 (
    .port_i (mixColumns_port_state_out_0_2_7[2:0]), //i
    .port_o (majority_5088_port_o                )  //o
  );
  Majority majority_5089 (
    .port_i (mixColumns_port_state_out_1_2_7[2:0]), //i
    .port_o (majority_5089_port_o                )  //o
  );
  Majority majority_5090 (
    .port_i (mixColumns_port_state_out_2_2_7[2:0]), //i
    .port_o (majority_5090_port_o                )  //o
  );
  Majority majority_5091 (
    .port_i (mixColumns_port_state_out_3_2_7[2:0]), //i
    .port_o (majority_5091_port_o                )  //o
  );
  Majority majority_5092 (
    .port_i (mixColumns_port_state_out_4_2_7[2:0]), //i
    .port_o (majority_5092_port_o                )  //o
  );
  Majority majority_5093 (
    .port_i (mixColumns_port_state_out_5_2_7[2:0]), //i
    .port_o (majority_5093_port_o                )  //o
  );
  Majority majority_5094 (
    .port_i (mixColumns_port_state_out_6_2_7[2:0]), //i
    .port_o (majority_5094_port_o                )  //o
  );
  Majority majority_5095 (
    .port_i (mixColumns_port_state_out_7_2_7[2:0]), //i
    .port_o (majority_5095_port_o                )  //o
  );
  Majority majority_5096 (
    .port_i (mixColumns_port_state_out_8_2_7[2:0]), //i
    .port_o (majority_5096_port_o                )  //o
  );
  Majority majority_5097 (
    .port_i (mixColumns_port_state_out_9_2_7[2:0]), //i
    .port_o (majority_5097_port_o                )  //o
  );
  Majority majority_5098 (
    .port_i (mixColumns_port_state_out_10_2_7[2:0]), //i
    .port_o (majority_5098_port_o                 )  //o
  );
  Majority majority_5099 (
    .port_i (mixColumns_port_state_out_11_2_7[2:0]), //i
    .port_o (majority_5099_port_o                 )  //o
  );
  Majority majority_5100 (
    .port_i (mixColumns_port_state_out_12_2_7[2:0]), //i
    .port_o (majority_5100_port_o                 )  //o
  );
  Majority majority_5101 (
    .port_i (mixColumns_port_state_out_13_2_7[2:0]), //i
    .port_o (majority_5101_port_o                 )  //o
  );
  Majority majority_5102 (
    .port_i (mixColumns_port_state_out_14_2_7[2:0]), //i
    .port_o (majority_5102_port_o                 )  //o
  );
  Majority majority_5103 (
    .port_i (mixColumns_port_state_out_15_2_7[2:0]), //i
    .port_o (majority_5103_port_o                 )  //o
  );
  Majority majority_5104 (
    .port_i (mixColumns_port_state_out_0_3_7[2:0]), //i
    .port_o (majority_5104_port_o                )  //o
  );
  Majority majority_5105 (
    .port_i (mixColumns_port_state_out_1_3_7[2:0]), //i
    .port_o (majority_5105_port_o                )  //o
  );
  Majority majority_5106 (
    .port_i (mixColumns_port_state_out_2_3_7[2:0]), //i
    .port_o (majority_5106_port_o                )  //o
  );
  Majority majority_5107 (
    .port_i (mixColumns_port_state_out_3_3_7[2:0]), //i
    .port_o (majority_5107_port_o                )  //o
  );
  Majority majority_5108 (
    .port_i (mixColumns_port_state_out_4_3_7[2:0]), //i
    .port_o (majority_5108_port_o                )  //o
  );
  Majority majority_5109 (
    .port_i (mixColumns_port_state_out_5_3_7[2:0]), //i
    .port_o (majority_5109_port_o                )  //o
  );
  Majority majority_5110 (
    .port_i (mixColumns_port_state_out_6_3_7[2:0]), //i
    .port_o (majority_5110_port_o                )  //o
  );
  Majority majority_5111 (
    .port_i (mixColumns_port_state_out_7_3_7[2:0]), //i
    .port_o (majority_5111_port_o                )  //o
  );
  Majority majority_5112 (
    .port_i (mixColumns_port_state_out_8_3_7[2:0]), //i
    .port_o (majority_5112_port_o                )  //o
  );
  Majority majority_5113 (
    .port_i (mixColumns_port_state_out_9_3_7[2:0]), //i
    .port_o (majority_5113_port_o                )  //o
  );
  Majority majority_5114 (
    .port_i (mixColumns_port_state_out_10_3_7[2:0]), //i
    .port_o (majority_5114_port_o                 )  //o
  );
  Majority majority_5115 (
    .port_i (mixColumns_port_state_out_11_3_7[2:0]), //i
    .port_o (majority_5115_port_o                 )  //o
  );
  Majority majority_5116 (
    .port_i (mixColumns_port_state_out_12_3_7[2:0]), //i
    .port_o (majority_5116_port_o                 )  //o
  );
  Majority majority_5117 (
    .port_i (mixColumns_port_state_out_13_3_7[2:0]), //i
    .port_o (majority_5117_port_o                 )  //o
  );
  Majority majority_5118 (
    .port_i (mixColumns_port_state_out_14_3_7[2:0]), //i
    .port_o (majority_5118_port_o                 )  //o
  );
  Majority majority_5119 (
    .port_i (mixColumns_port_state_out_15_3_7[2:0]), //i
    .port_o (majority_5119_port_o                 )  //o
  );
  Majority majority_5120 (
    .port_i (mixColumns_port_state_out_0_0_0[2:0]), //i
    .port_o (majority_5120_port_o                )  //o
  );
  Majority majority_5121 (
    .port_i (mixColumns_port_state_out_1_0_0[2:0]), //i
    .port_o (majority_5121_port_o                )  //o
  );
  Majority majority_5122 (
    .port_i (mixColumns_port_state_out_2_0_0[2:0]), //i
    .port_o (majority_5122_port_o                )  //o
  );
  Majority majority_5123 (
    .port_i (mixColumns_port_state_out_3_0_0[2:0]), //i
    .port_o (majority_5123_port_o                )  //o
  );
  Majority majority_5124 (
    .port_i (mixColumns_port_state_out_4_0_0[2:0]), //i
    .port_o (majority_5124_port_o                )  //o
  );
  Majority majority_5125 (
    .port_i (mixColumns_port_state_out_5_0_0[2:0]), //i
    .port_o (majority_5125_port_o                )  //o
  );
  Majority majority_5126 (
    .port_i (mixColumns_port_state_out_6_0_0[2:0]), //i
    .port_o (majority_5126_port_o                )  //o
  );
  Majority majority_5127 (
    .port_i (mixColumns_port_state_out_7_0_0[2:0]), //i
    .port_o (majority_5127_port_o                )  //o
  );
  Majority majority_5128 (
    .port_i (mixColumns_port_state_out_8_0_0[2:0]), //i
    .port_o (majority_5128_port_o                )  //o
  );
  Majority majority_5129 (
    .port_i (mixColumns_port_state_out_9_0_0[2:0]), //i
    .port_o (majority_5129_port_o                )  //o
  );
  Majority majority_5130 (
    .port_i (mixColumns_port_state_out_10_0_0[2:0]), //i
    .port_o (majority_5130_port_o                 )  //o
  );
  Majority majority_5131 (
    .port_i (mixColumns_port_state_out_11_0_0[2:0]), //i
    .port_o (majority_5131_port_o                 )  //o
  );
  Majority majority_5132 (
    .port_i (mixColumns_port_state_out_12_0_0[2:0]), //i
    .port_o (majority_5132_port_o                 )  //o
  );
  Majority majority_5133 (
    .port_i (mixColumns_port_state_out_13_0_0[2:0]), //i
    .port_o (majority_5133_port_o                 )  //o
  );
  Majority majority_5134 (
    .port_i (mixColumns_port_state_out_14_0_0[2:0]), //i
    .port_o (majority_5134_port_o                 )  //o
  );
  Majority majority_5135 (
    .port_i (mixColumns_port_state_out_15_0_0[2:0]), //i
    .port_o (majority_5135_port_o                 )  //o
  );
  Majority majority_5136 (
    .port_i (mixColumns_port_state_out_0_1_0[2:0]), //i
    .port_o (majority_5136_port_o                )  //o
  );
  Majority majority_5137 (
    .port_i (mixColumns_port_state_out_1_1_0[2:0]), //i
    .port_o (majority_5137_port_o                )  //o
  );
  Majority majority_5138 (
    .port_i (mixColumns_port_state_out_2_1_0[2:0]), //i
    .port_o (majority_5138_port_o                )  //o
  );
  Majority majority_5139 (
    .port_i (mixColumns_port_state_out_3_1_0[2:0]), //i
    .port_o (majority_5139_port_o                )  //o
  );
  Majority majority_5140 (
    .port_i (mixColumns_port_state_out_4_1_0[2:0]), //i
    .port_o (majority_5140_port_o                )  //o
  );
  Majority majority_5141 (
    .port_i (mixColumns_port_state_out_5_1_0[2:0]), //i
    .port_o (majority_5141_port_o                )  //o
  );
  Majority majority_5142 (
    .port_i (mixColumns_port_state_out_6_1_0[2:0]), //i
    .port_o (majority_5142_port_o                )  //o
  );
  Majority majority_5143 (
    .port_i (mixColumns_port_state_out_7_1_0[2:0]), //i
    .port_o (majority_5143_port_o                )  //o
  );
  Majority majority_5144 (
    .port_i (mixColumns_port_state_out_8_1_0[2:0]), //i
    .port_o (majority_5144_port_o                )  //o
  );
  Majority majority_5145 (
    .port_i (mixColumns_port_state_out_9_1_0[2:0]), //i
    .port_o (majority_5145_port_o                )  //o
  );
  Majority majority_5146 (
    .port_i (mixColumns_port_state_out_10_1_0[2:0]), //i
    .port_o (majority_5146_port_o                 )  //o
  );
  Majority majority_5147 (
    .port_i (mixColumns_port_state_out_11_1_0[2:0]), //i
    .port_o (majority_5147_port_o                 )  //o
  );
  Majority majority_5148 (
    .port_i (mixColumns_port_state_out_12_1_0[2:0]), //i
    .port_o (majority_5148_port_o                 )  //o
  );
  Majority majority_5149 (
    .port_i (mixColumns_port_state_out_13_1_0[2:0]), //i
    .port_o (majority_5149_port_o                 )  //o
  );
  Majority majority_5150 (
    .port_i (mixColumns_port_state_out_14_1_0[2:0]), //i
    .port_o (majority_5150_port_o                 )  //o
  );
  Majority majority_5151 (
    .port_i (mixColumns_port_state_out_15_1_0[2:0]), //i
    .port_o (majority_5151_port_o                 )  //o
  );
  Majority majority_5152 (
    .port_i (mixColumns_port_state_out_0_2_0[2:0]), //i
    .port_o (majority_5152_port_o                )  //o
  );
  Majority majority_5153 (
    .port_i (mixColumns_port_state_out_1_2_0[2:0]), //i
    .port_o (majority_5153_port_o                )  //o
  );
  Majority majority_5154 (
    .port_i (mixColumns_port_state_out_2_2_0[2:0]), //i
    .port_o (majority_5154_port_o                )  //o
  );
  Majority majority_5155 (
    .port_i (mixColumns_port_state_out_3_2_0[2:0]), //i
    .port_o (majority_5155_port_o                )  //o
  );
  Majority majority_5156 (
    .port_i (mixColumns_port_state_out_4_2_0[2:0]), //i
    .port_o (majority_5156_port_o                )  //o
  );
  Majority majority_5157 (
    .port_i (mixColumns_port_state_out_5_2_0[2:0]), //i
    .port_o (majority_5157_port_o                )  //o
  );
  Majority majority_5158 (
    .port_i (mixColumns_port_state_out_6_2_0[2:0]), //i
    .port_o (majority_5158_port_o                )  //o
  );
  Majority majority_5159 (
    .port_i (mixColumns_port_state_out_7_2_0[2:0]), //i
    .port_o (majority_5159_port_o                )  //o
  );
  Majority majority_5160 (
    .port_i (mixColumns_port_state_out_8_2_0[2:0]), //i
    .port_o (majority_5160_port_o                )  //o
  );
  Majority majority_5161 (
    .port_i (mixColumns_port_state_out_9_2_0[2:0]), //i
    .port_o (majority_5161_port_o                )  //o
  );
  Majority majority_5162 (
    .port_i (mixColumns_port_state_out_10_2_0[2:0]), //i
    .port_o (majority_5162_port_o                 )  //o
  );
  Majority majority_5163 (
    .port_i (mixColumns_port_state_out_11_2_0[2:0]), //i
    .port_o (majority_5163_port_o                 )  //o
  );
  Majority majority_5164 (
    .port_i (mixColumns_port_state_out_12_2_0[2:0]), //i
    .port_o (majority_5164_port_o                 )  //o
  );
  Majority majority_5165 (
    .port_i (mixColumns_port_state_out_13_2_0[2:0]), //i
    .port_o (majority_5165_port_o                 )  //o
  );
  Majority majority_5166 (
    .port_i (mixColumns_port_state_out_14_2_0[2:0]), //i
    .port_o (majority_5166_port_o                 )  //o
  );
  Majority majority_5167 (
    .port_i (mixColumns_port_state_out_15_2_0[2:0]), //i
    .port_o (majority_5167_port_o                 )  //o
  );
  Majority majority_5168 (
    .port_i (mixColumns_port_state_out_0_3_0[2:0]), //i
    .port_o (majority_5168_port_o                )  //o
  );
  Majority majority_5169 (
    .port_i (mixColumns_port_state_out_1_3_0[2:0]), //i
    .port_o (majority_5169_port_o                )  //o
  );
  Majority majority_5170 (
    .port_i (mixColumns_port_state_out_2_3_0[2:0]), //i
    .port_o (majority_5170_port_o                )  //o
  );
  Majority majority_5171 (
    .port_i (mixColumns_port_state_out_3_3_0[2:0]), //i
    .port_o (majority_5171_port_o                )  //o
  );
  Majority majority_5172 (
    .port_i (mixColumns_port_state_out_4_3_0[2:0]), //i
    .port_o (majority_5172_port_o                )  //o
  );
  Majority majority_5173 (
    .port_i (mixColumns_port_state_out_5_3_0[2:0]), //i
    .port_o (majority_5173_port_o                )  //o
  );
  Majority majority_5174 (
    .port_i (mixColumns_port_state_out_6_3_0[2:0]), //i
    .port_o (majority_5174_port_o                )  //o
  );
  Majority majority_5175 (
    .port_i (mixColumns_port_state_out_7_3_0[2:0]), //i
    .port_o (majority_5175_port_o                )  //o
  );
  Majority majority_5176 (
    .port_i (mixColumns_port_state_out_8_3_0[2:0]), //i
    .port_o (majority_5176_port_o                )  //o
  );
  Majority majority_5177 (
    .port_i (mixColumns_port_state_out_9_3_0[2:0]), //i
    .port_o (majority_5177_port_o                )  //o
  );
  Majority majority_5178 (
    .port_i (mixColumns_port_state_out_10_3_0[2:0]), //i
    .port_o (majority_5178_port_o                 )  //o
  );
  Majority majority_5179 (
    .port_i (mixColumns_port_state_out_11_3_0[2:0]), //i
    .port_o (majority_5179_port_o                 )  //o
  );
  Majority majority_5180 (
    .port_i (mixColumns_port_state_out_12_3_0[2:0]), //i
    .port_o (majority_5180_port_o                 )  //o
  );
  Majority majority_5181 (
    .port_i (mixColumns_port_state_out_13_3_0[2:0]), //i
    .port_o (majority_5181_port_o                 )  //o
  );
  Majority majority_5182 (
    .port_i (mixColumns_port_state_out_14_3_0[2:0]), //i
    .port_o (majority_5182_port_o                 )  //o
  );
  Majority majority_5183 (
    .port_i (mixColumns_port_state_out_15_3_0[2:0]), //i
    .port_o (majority_5183_port_o                 )  //o
  );
  Majority majority_5184 (
    .port_i (mixColumns_port_state_out_0_0_1[2:0]), //i
    .port_o (majority_5184_port_o                )  //o
  );
  Majority majority_5185 (
    .port_i (mixColumns_port_state_out_1_0_1[2:0]), //i
    .port_o (majority_5185_port_o                )  //o
  );
  Majority majority_5186 (
    .port_i (mixColumns_port_state_out_2_0_1[2:0]), //i
    .port_o (majority_5186_port_o                )  //o
  );
  Majority majority_5187 (
    .port_i (mixColumns_port_state_out_3_0_1[2:0]), //i
    .port_o (majority_5187_port_o                )  //o
  );
  Majority majority_5188 (
    .port_i (mixColumns_port_state_out_4_0_1[2:0]), //i
    .port_o (majority_5188_port_o                )  //o
  );
  Majority majority_5189 (
    .port_i (mixColumns_port_state_out_5_0_1[2:0]), //i
    .port_o (majority_5189_port_o                )  //o
  );
  Majority majority_5190 (
    .port_i (mixColumns_port_state_out_6_0_1[2:0]), //i
    .port_o (majority_5190_port_o                )  //o
  );
  Majority majority_5191 (
    .port_i (mixColumns_port_state_out_7_0_1[2:0]), //i
    .port_o (majority_5191_port_o                )  //o
  );
  Majority majority_5192 (
    .port_i (mixColumns_port_state_out_8_0_1[2:0]), //i
    .port_o (majority_5192_port_o                )  //o
  );
  Majority majority_5193 (
    .port_i (mixColumns_port_state_out_9_0_1[2:0]), //i
    .port_o (majority_5193_port_o                )  //o
  );
  Majority majority_5194 (
    .port_i (mixColumns_port_state_out_10_0_1[2:0]), //i
    .port_o (majority_5194_port_o                 )  //o
  );
  Majority majority_5195 (
    .port_i (mixColumns_port_state_out_11_0_1[2:0]), //i
    .port_o (majority_5195_port_o                 )  //o
  );
  Majority majority_5196 (
    .port_i (mixColumns_port_state_out_12_0_1[2:0]), //i
    .port_o (majority_5196_port_o                 )  //o
  );
  Majority majority_5197 (
    .port_i (mixColumns_port_state_out_13_0_1[2:0]), //i
    .port_o (majority_5197_port_o                 )  //o
  );
  Majority majority_5198 (
    .port_i (mixColumns_port_state_out_14_0_1[2:0]), //i
    .port_o (majority_5198_port_o                 )  //o
  );
  Majority majority_5199 (
    .port_i (mixColumns_port_state_out_15_0_1[2:0]), //i
    .port_o (majority_5199_port_o                 )  //o
  );
  Majority majority_5200 (
    .port_i (mixColumns_port_state_out_0_1_1[2:0]), //i
    .port_o (majority_5200_port_o                )  //o
  );
  Majority majority_5201 (
    .port_i (mixColumns_port_state_out_1_1_1[2:0]), //i
    .port_o (majority_5201_port_o                )  //o
  );
  Majority majority_5202 (
    .port_i (mixColumns_port_state_out_2_1_1[2:0]), //i
    .port_o (majority_5202_port_o                )  //o
  );
  Majority majority_5203 (
    .port_i (mixColumns_port_state_out_3_1_1[2:0]), //i
    .port_o (majority_5203_port_o                )  //o
  );
  Majority majority_5204 (
    .port_i (mixColumns_port_state_out_4_1_1[2:0]), //i
    .port_o (majority_5204_port_o                )  //o
  );
  Majority majority_5205 (
    .port_i (mixColumns_port_state_out_5_1_1[2:0]), //i
    .port_o (majority_5205_port_o                )  //o
  );
  Majority majority_5206 (
    .port_i (mixColumns_port_state_out_6_1_1[2:0]), //i
    .port_o (majority_5206_port_o                )  //o
  );
  Majority majority_5207 (
    .port_i (mixColumns_port_state_out_7_1_1[2:0]), //i
    .port_o (majority_5207_port_o                )  //o
  );
  Majority majority_5208 (
    .port_i (mixColumns_port_state_out_8_1_1[2:0]), //i
    .port_o (majority_5208_port_o                )  //o
  );
  Majority majority_5209 (
    .port_i (mixColumns_port_state_out_9_1_1[2:0]), //i
    .port_o (majority_5209_port_o                )  //o
  );
  Majority majority_5210 (
    .port_i (mixColumns_port_state_out_10_1_1[2:0]), //i
    .port_o (majority_5210_port_o                 )  //o
  );
  Majority majority_5211 (
    .port_i (mixColumns_port_state_out_11_1_1[2:0]), //i
    .port_o (majority_5211_port_o                 )  //o
  );
  Majority majority_5212 (
    .port_i (mixColumns_port_state_out_12_1_1[2:0]), //i
    .port_o (majority_5212_port_o                 )  //o
  );
  Majority majority_5213 (
    .port_i (mixColumns_port_state_out_13_1_1[2:0]), //i
    .port_o (majority_5213_port_o                 )  //o
  );
  Majority majority_5214 (
    .port_i (mixColumns_port_state_out_14_1_1[2:0]), //i
    .port_o (majority_5214_port_o                 )  //o
  );
  Majority majority_5215 (
    .port_i (mixColumns_port_state_out_15_1_1[2:0]), //i
    .port_o (majority_5215_port_o                 )  //o
  );
  Majority majority_5216 (
    .port_i (mixColumns_port_state_out_0_2_1[2:0]), //i
    .port_o (majority_5216_port_o                )  //o
  );
  Majority majority_5217 (
    .port_i (mixColumns_port_state_out_1_2_1[2:0]), //i
    .port_o (majority_5217_port_o                )  //o
  );
  Majority majority_5218 (
    .port_i (mixColumns_port_state_out_2_2_1[2:0]), //i
    .port_o (majority_5218_port_o                )  //o
  );
  Majority majority_5219 (
    .port_i (mixColumns_port_state_out_3_2_1[2:0]), //i
    .port_o (majority_5219_port_o                )  //o
  );
  Majority majority_5220 (
    .port_i (mixColumns_port_state_out_4_2_1[2:0]), //i
    .port_o (majority_5220_port_o                )  //o
  );
  Majority majority_5221 (
    .port_i (mixColumns_port_state_out_5_2_1[2:0]), //i
    .port_o (majority_5221_port_o                )  //o
  );
  Majority majority_5222 (
    .port_i (mixColumns_port_state_out_6_2_1[2:0]), //i
    .port_o (majority_5222_port_o                )  //o
  );
  Majority majority_5223 (
    .port_i (mixColumns_port_state_out_7_2_1[2:0]), //i
    .port_o (majority_5223_port_o                )  //o
  );
  Majority majority_5224 (
    .port_i (mixColumns_port_state_out_8_2_1[2:0]), //i
    .port_o (majority_5224_port_o                )  //o
  );
  Majority majority_5225 (
    .port_i (mixColumns_port_state_out_9_2_1[2:0]), //i
    .port_o (majority_5225_port_o                )  //o
  );
  Majority majority_5226 (
    .port_i (mixColumns_port_state_out_10_2_1[2:0]), //i
    .port_o (majority_5226_port_o                 )  //o
  );
  Majority majority_5227 (
    .port_i (mixColumns_port_state_out_11_2_1[2:0]), //i
    .port_o (majority_5227_port_o                 )  //o
  );
  Majority majority_5228 (
    .port_i (mixColumns_port_state_out_12_2_1[2:0]), //i
    .port_o (majority_5228_port_o                 )  //o
  );
  Majority majority_5229 (
    .port_i (mixColumns_port_state_out_13_2_1[2:0]), //i
    .port_o (majority_5229_port_o                 )  //o
  );
  Majority majority_5230 (
    .port_i (mixColumns_port_state_out_14_2_1[2:0]), //i
    .port_o (majority_5230_port_o                 )  //o
  );
  Majority majority_5231 (
    .port_i (mixColumns_port_state_out_15_2_1[2:0]), //i
    .port_o (majority_5231_port_o                 )  //o
  );
  Majority majority_5232 (
    .port_i (mixColumns_port_state_out_0_3_1[2:0]), //i
    .port_o (majority_5232_port_o                )  //o
  );
  Majority majority_5233 (
    .port_i (mixColumns_port_state_out_1_3_1[2:0]), //i
    .port_o (majority_5233_port_o                )  //o
  );
  Majority majority_5234 (
    .port_i (mixColumns_port_state_out_2_3_1[2:0]), //i
    .port_o (majority_5234_port_o                )  //o
  );
  Majority majority_5235 (
    .port_i (mixColumns_port_state_out_3_3_1[2:0]), //i
    .port_o (majority_5235_port_o                )  //o
  );
  Majority majority_5236 (
    .port_i (mixColumns_port_state_out_4_3_1[2:0]), //i
    .port_o (majority_5236_port_o                )  //o
  );
  Majority majority_5237 (
    .port_i (mixColumns_port_state_out_5_3_1[2:0]), //i
    .port_o (majority_5237_port_o                )  //o
  );
  Majority majority_5238 (
    .port_i (mixColumns_port_state_out_6_3_1[2:0]), //i
    .port_o (majority_5238_port_o                )  //o
  );
  Majority majority_5239 (
    .port_i (mixColumns_port_state_out_7_3_1[2:0]), //i
    .port_o (majority_5239_port_o                )  //o
  );
  Majority majority_5240 (
    .port_i (mixColumns_port_state_out_8_3_1[2:0]), //i
    .port_o (majority_5240_port_o                )  //o
  );
  Majority majority_5241 (
    .port_i (mixColumns_port_state_out_9_3_1[2:0]), //i
    .port_o (majority_5241_port_o                )  //o
  );
  Majority majority_5242 (
    .port_i (mixColumns_port_state_out_10_3_1[2:0]), //i
    .port_o (majority_5242_port_o                 )  //o
  );
  Majority majority_5243 (
    .port_i (mixColumns_port_state_out_11_3_1[2:0]), //i
    .port_o (majority_5243_port_o                 )  //o
  );
  Majority majority_5244 (
    .port_i (mixColumns_port_state_out_12_3_1[2:0]), //i
    .port_o (majority_5244_port_o                 )  //o
  );
  Majority majority_5245 (
    .port_i (mixColumns_port_state_out_13_3_1[2:0]), //i
    .port_o (majority_5245_port_o                 )  //o
  );
  Majority majority_5246 (
    .port_i (mixColumns_port_state_out_14_3_1[2:0]), //i
    .port_o (majority_5246_port_o                 )  //o
  );
  Majority majority_5247 (
    .port_i (mixColumns_port_state_out_15_3_1[2:0]), //i
    .port_o (majority_5247_port_o                 )  //o
  );
  Majority majority_5248 (
    .port_i (mixColumns_port_state_out_0_0_2[2:0]), //i
    .port_o (majority_5248_port_o                )  //o
  );
  Majority majority_5249 (
    .port_i (mixColumns_port_state_out_1_0_2[2:0]), //i
    .port_o (majority_5249_port_o                )  //o
  );
  Majority majority_5250 (
    .port_i (mixColumns_port_state_out_2_0_2[2:0]), //i
    .port_o (majority_5250_port_o                )  //o
  );
  Majority majority_5251 (
    .port_i (mixColumns_port_state_out_3_0_2[2:0]), //i
    .port_o (majority_5251_port_o                )  //o
  );
  Majority majority_5252 (
    .port_i (mixColumns_port_state_out_4_0_2[2:0]), //i
    .port_o (majority_5252_port_o                )  //o
  );
  Majority majority_5253 (
    .port_i (mixColumns_port_state_out_5_0_2[2:0]), //i
    .port_o (majority_5253_port_o                )  //o
  );
  Majority majority_5254 (
    .port_i (mixColumns_port_state_out_6_0_2[2:0]), //i
    .port_o (majority_5254_port_o                )  //o
  );
  Majority majority_5255 (
    .port_i (mixColumns_port_state_out_7_0_2[2:0]), //i
    .port_o (majority_5255_port_o                )  //o
  );
  Majority majority_5256 (
    .port_i (mixColumns_port_state_out_8_0_2[2:0]), //i
    .port_o (majority_5256_port_o                )  //o
  );
  Majority majority_5257 (
    .port_i (mixColumns_port_state_out_9_0_2[2:0]), //i
    .port_o (majority_5257_port_o                )  //o
  );
  Majority majority_5258 (
    .port_i (mixColumns_port_state_out_10_0_2[2:0]), //i
    .port_o (majority_5258_port_o                 )  //o
  );
  Majority majority_5259 (
    .port_i (mixColumns_port_state_out_11_0_2[2:0]), //i
    .port_o (majority_5259_port_o                 )  //o
  );
  Majority majority_5260 (
    .port_i (mixColumns_port_state_out_12_0_2[2:0]), //i
    .port_o (majority_5260_port_o                 )  //o
  );
  Majority majority_5261 (
    .port_i (mixColumns_port_state_out_13_0_2[2:0]), //i
    .port_o (majority_5261_port_o                 )  //o
  );
  Majority majority_5262 (
    .port_i (mixColumns_port_state_out_14_0_2[2:0]), //i
    .port_o (majority_5262_port_o                 )  //o
  );
  Majority majority_5263 (
    .port_i (mixColumns_port_state_out_15_0_2[2:0]), //i
    .port_o (majority_5263_port_o                 )  //o
  );
  Majority majority_5264 (
    .port_i (mixColumns_port_state_out_0_1_2[2:0]), //i
    .port_o (majority_5264_port_o                )  //o
  );
  Majority majority_5265 (
    .port_i (mixColumns_port_state_out_1_1_2[2:0]), //i
    .port_o (majority_5265_port_o                )  //o
  );
  Majority majority_5266 (
    .port_i (mixColumns_port_state_out_2_1_2[2:0]), //i
    .port_o (majority_5266_port_o                )  //o
  );
  Majority majority_5267 (
    .port_i (mixColumns_port_state_out_3_1_2[2:0]), //i
    .port_o (majority_5267_port_o                )  //o
  );
  Majority majority_5268 (
    .port_i (mixColumns_port_state_out_4_1_2[2:0]), //i
    .port_o (majority_5268_port_o                )  //o
  );
  Majority majority_5269 (
    .port_i (mixColumns_port_state_out_5_1_2[2:0]), //i
    .port_o (majority_5269_port_o                )  //o
  );
  Majority majority_5270 (
    .port_i (mixColumns_port_state_out_6_1_2[2:0]), //i
    .port_o (majority_5270_port_o                )  //o
  );
  Majority majority_5271 (
    .port_i (mixColumns_port_state_out_7_1_2[2:0]), //i
    .port_o (majority_5271_port_o                )  //o
  );
  Majority majority_5272 (
    .port_i (mixColumns_port_state_out_8_1_2[2:0]), //i
    .port_o (majority_5272_port_o                )  //o
  );
  Majority majority_5273 (
    .port_i (mixColumns_port_state_out_9_1_2[2:0]), //i
    .port_o (majority_5273_port_o                )  //o
  );
  Majority majority_5274 (
    .port_i (mixColumns_port_state_out_10_1_2[2:0]), //i
    .port_o (majority_5274_port_o                 )  //o
  );
  Majority majority_5275 (
    .port_i (mixColumns_port_state_out_11_1_2[2:0]), //i
    .port_o (majority_5275_port_o                 )  //o
  );
  Majority majority_5276 (
    .port_i (mixColumns_port_state_out_12_1_2[2:0]), //i
    .port_o (majority_5276_port_o                 )  //o
  );
  Majority majority_5277 (
    .port_i (mixColumns_port_state_out_13_1_2[2:0]), //i
    .port_o (majority_5277_port_o                 )  //o
  );
  Majority majority_5278 (
    .port_i (mixColumns_port_state_out_14_1_2[2:0]), //i
    .port_o (majority_5278_port_o                 )  //o
  );
  Majority majority_5279 (
    .port_i (mixColumns_port_state_out_15_1_2[2:0]), //i
    .port_o (majority_5279_port_o                 )  //o
  );
  Majority majority_5280 (
    .port_i (mixColumns_port_state_out_0_2_2[2:0]), //i
    .port_o (majority_5280_port_o                )  //o
  );
  Majority majority_5281 (
    .port_i (mixColumns_port_state_out_1_2_2[2:0]), //i
    .port_o (majority_5281_port_o                )  //o
  );
  Majority majority_5282 (
    .port_i (mixColumns_port_state_out_2_2_2[2:0]), //i
    .port_o (majority_5282_port_o                )  //o
  );
  Majority majority_5283 (
    .port_i (mixColumns_port_state_out_3_2_2[2:0]), //i
    .port_o (majority_5283_port_o                )  //o
  );
  Majority majority_5284 (
    .port_i (mixColumns_port_state_out_4_2_2[2:0]), //i
    .port_o (majority_5284_port_o                )  //o
  );
  Majority majority_5285 (
    .port_i (mixColumns_port_state_out_5_2_2[2:0]), //i
    .port_o (majority_5285_port_o                )  //o
  );
  Majority majority_5286 (
    .port_i (mixColumns_port_state_out_6_2_2[2:0]), //i
    .port_o (majority_5286_port_o                )  //o
  );
  Majority majority_5287 (
    .port_i (mixColumns_port_state_out_7_2_2[2:0]), //i
    .port_o (majority_5287_port_o                )  //o
  );
  Majority majority_5288 (
    .port_i (mixColumns_port_state_out_8_2_2[2:0]), //i
    .port_o (majority_5288_port_o                )  //o
  );
  Majority majority_5289 (
    .port_i (mixColumns_port_state_out_9_2_2[2:0]), //i
    .port_o (majority_5289_port_o                )  //o
  );
  Majority majority_5290 (
    .port_i (mixColumns_port_state_out_10_2_2[2:0]), //i
    .port_o (majority_5290_port_o                 )  //o
  );
  Majority majority_5291 (
    .port_i (mixColumns_port_state_out_11_2_2[2:0]), //i
    .port_o (majority_5291_port_o                 )  //o
  );
  Majority majority_5292 (
    .port_i (mixColumns_port_state_out_12_2_2[2:0]), //i
    .port_o (majority_5292_port_o                 )  //o
  );
  Majority majority_5293 (
    .port_i (mixColumns_port_state_out_13_2_2[2:0]), //i
    .port_o (majority_5293_port_o                 )  //o
  );
  Majority majority_5294 (
    .port_i (mixColumns_port_state_out_14_2_2[2:0]), //i
    .port_o (majority_5294_port_o                 )  //o
  );
  Majority majority_5295 (
    .port_i (mixColumns_port_state_out_15_2_2[2:0]), //i
    .port_o (majority_5295_port_o                 )  //o
  );
  Majority majority_5296 (
    .port_i (mixColumns_port_state_out_0_3_2[2:0]), //i
    .port_o (majority_5296_port_o                )  //o
  );
  Majority majority_5297 (
    .port_i (mixColumns_port_state_out_1_3_2[2:0]), //i
    .port_o (majority_5297_port_o                )  //o
  );
  Majority majority_5298 (
    .port_i (mixColumns_port_state_out_2_3_2[2:0]), //i
    .port_o (majority_5298_port_o                )  //o
  );
  Majority majority_5299 (
    .port_i (mixColumns_port_state_out_3_3_2[2:0]), //i
    .port_o (majority_5299_port_o                )  //o
  );
  Majority majority_5300 (
    .port_i (mixColumns_port_state_out_4_3_2[2:0]), //i
    .port_o (majority_5300_port_o                )  //o
  );
  Majority majority_5301 (
    .port_i (mixColumns_port_state_out_5_3_2[2:0]), //i
    .port_o (majority_5301_port_o                )  //o
  );
  Majority majority_5302 (
    .port_i (mixColumns_port_state_out_6_3_2[2:0]), //i
    .port_o (majority_5302_port_o                )  //o
  );
  Majority majority_5303 (
    .port_i (mixColumns_port_state_out_7_3_2[2:0]), //i
    .port_o (majority_5303_port_o                )  //o
  );
  Majority majority_5304 (
    .port_i (mixColumns_port_state_out_8_3_2[2:0]), //i
    .port_o (majority_5304_port_o                )  //o
  );
  Majority majority_5305 (
    .port_i (mixColumns_port_state_out_9_3_2[2:0]), //i
    .port_o (majority_5305_port_o                )  //o
  );
  Majority majority_5306 (
    .port_i (mixColumns_port_state_out_10_3_2[2:0]), //i
    .port_o (majority_5306_port_o                 )  //o
  );
  Majority majority_5307 (
    .port_i (mixColumns_port_state_out_11_3_2[2:0]), //i
    .port_o (majority_5307_port_o                 )  //o
  );
  Majority majority_5308 (
    .port_i (mixColumns_port_state_out_12_3_2[2:0]), //i
    .port_o (majority_5308_port_o                 )  //o
  );
  Majority majority_5309 (
    .port_i (mixColumns_port_state_out_13_3_2[2:0]), //i
    .port_o (majority_5309_port_o                 )  //o
  );
  Majority majority_5310 (
    .port_i (mixColumns_port_state_out_14_3_2[2:0]), //i
    .port_o (majority_5310_port_o                 )  //o
  );
  Majority majority_5311 (
    .port_i (mixColumns_port_state_out_15_3_2[2:0]), //i
    .port_o (majority_5311_port_o                 )  //o
  );
  Majority majority_5312 (
    .port_i (mixColumns_port_state_out_0_0_3[2:0]), //i
    .port_o (majority_5312_port_o                )  //o
  );
  Majority majority_5313 (
    .port_i (mixColumns_port_state_out_1_0_3[2:0]), //i
    .port_o (majority_5313_port_o                )  //o
  );
  Majority majority_5314 (
    .port_i (mixColumns_port_state_out_2_0_3[2:0]), //i
    .port_o (majority_5314_port_o                )  //o
  );
  Majority majority_5315 (
    .port_i (mixColumns_port_state_out_3_0_3[2:0]), //i
    .port_o (majority_5315_port_o                )  //o
  );
  Majority majority_5316 (
    .port_i (mixColumns_port_state_out_4_0_3[2:0]), //i
    .port_o (majority_5316_port_o                )  //o
  );
  Majority majority_5317 (
    .port_i (mixColumns_port_state_out_5_0_3[2:0]), //i
    .port_o (majority_5317_port_o                )  //o
  );
  Majority majority_5318 (
    .port_i (mixColumns_port_state_out_6_0_3[2:0]), //i
    .port_o (majority_5318_port_o                )  //o
  );
  Majority majority_5319 (
    .port_i (mixColumns_port_state_out_7_0_3[2:0]), //i
    .port_o (majority_5319_port_o                )  //o
  );
  Majority majority_5320 (
    .port_i (mixColumns_port_state_out_8_0_3[2:0]), //i
    .port_o (majority_5320_port_o                )  //o
  );
  Majority majority_5321 (
    .port_i (mixColumns_port_state_out_9_0_3[2:0]), //i
    .port_o (majority_5321_port_o                )  //o
  );
  Majority majority_5322 (
    .port_i (mixColumns_port_state_out_10_0_3[2:0]), //i
    .port_o (majority_5322_port_o                 )  //o
  );
  Majority majority_5323 (
    .port_i (mixColumns_port_state_out_11_0_3[2:0]), //i
    .port_o (majority_5323_port_o                 )  //o
  );
  Majority majority_5324 (
    .port_i (mixColumns_port_state_out_12_0_3[2:0]), //i
    .port_o (majority_5324_port_o                 )  //o
  );
  Majority majority_5325 (
    .port_i (mixColumns_port_state_out_13_0_3[2:0]), //i
    .port_o (majority_5325_port_o                 )  //o
  );
  Majority majority_5326 (
    .port_i (mixColumns_port_state_out_14_0_3[2:0]), //i
    .port_o (majority_5326_port_o                 )  //o
  );
  Majority majority_5327 (
    .port_i (mixColumns_port_state_out_15_0_3[2:0]), //i
    .port_o (majority_5327_port_o                 )  //o
  );
  Majority majority_5328 (
    .port_i (mixColumns_port_state_out_0_1_3[2:0]), //i
    .port_o (majority_5328_port_o                )  //o
  );
  Majority majority_5329 (
    .port_i (mixColumns_port_state_out_1_1_3[2:0]), //i
    .port_o (majority_5329_port_o                )  //o
  );
  Majority majority_5330 (
    .port_i (mixColumns_port_state_out_2_1_3[2:0]), //i
    .port_o (majority_5330_port_o                )  //o
  );
  Majority majority_5331 (
    .port_i (mixColumns_port_state_out_3_1_3[2:0]), //i
    .port_o (majority_5331_port_o                )  //o
  );
  Majority majority_5332 (
    .port_i (mixColumns_port_state_out_4_1_3[2:0]), //i
    .port_o (majority_5332_port_o                )  //o
  );
  Majority majority_5333 (
    .port_i (mixColumns_port_state_out_5_1_3[2:0]), //i
    .port_o (majority_5333_port_o                )  //o
  );
  Majority majority_5334 (
    .port_i (mixColumns_port_state_out_6_1_3[2:0]), //i
    .port_o (majority_5334_port_o                )  //o
  );
  Majority majority_5335 (
    .port_i (mixColumns_port_state_out_7_1_3[2:0]), //i
    .port_o (majority_5335_port_o                )  //o
  );
  Majority majority_5336 (
    .port_i (mixColumns_port_state_out_8_1_3[2:0]), //i
    .port_o (majority_5336_port_o                )  //o
  );
  Majority majority_5337 (
    .port_i (mixColumns_port_state_out_9_1_3[2:0]), //i
    .port_o (majority_5337_port_o                )  //o
  );
  Majority majority_5338 (
    .port_i (mixColumns_port_state_out_10_1_3[2:0]), //i
    .port_o (majority_5338_port_o                 )  //o
  );
  Majority majority_5339 (
    .port_i (mixColumns_port_state_out_11_1_3[2:0]), //i
    .port_o (majority_5339_port_o                 )  //o
  );
  Majority majority_5340 (
    .port_i (mixColumns_port_state_out_12_1_3[2:0]), //i
    .port_o (majority_5340_port_o                 )  //o
  );
  Majority majority_5341 (
    .port_i (mixColumns_port_state_out_13_1_3[2:0]), //i
    .port_o (majority_5341_port_o                 )  //o
  );
  Majority majority_5342 (
    .port_i (mixColumns_port_state_out_14_1_3[2:0]), //i
    .port_o (majority_5342_port_o                 )  //o
  );
  Majority majority_5343 (
    .port_i (mixColumns_port_state_out_15_1_3[2:0]), //i
    .port_o (majority_5343_port_o                 )  //o
  );
  Majority majority_5344 (
    .port_i (mixColumns_port_state_out_0_2_3[2:0]), //i
    .port_o (majority_5344_port_o                )  //o
  );
  Majority majority_5345 (
    .port_i (mixColumns_port_state_out_1_2_3[2:0]), //i
    .port_o (majority_5345_port_o                )  //o
  );
  Majority majority_5346 (
    .port_i (mixColumns_port_state_out_2_2_3[2:0]), //i
    .port_o (majority_5346_port_o                )  //o
  );
  Majority majority_5347 (
    .port_i (mixColumns_port_state_out_3_2_3[2:0]), //i
    .port_o (majority_5347_port_o                )  //o
  );
  Majority majority_5348 (
    .port_i (mixColumns_port_state_out_4_2_3[2:0]), //i
    .port_o (majority_5348_port_o                )  //o
  );
  Majority majority_5349 (
    .port_i (mixColumns_port_state_out_5_2_3[2:0]), //i
    .port_o (majority_5349_port_o                )  //o
  );
  Majority majority_5350 (
    .port_i (mixColumns_port_state_out_6_2_3[2:0]), //i
    .port_o (majority_5350_port_o                )  //o
  );
  Majority majority_5351 (
    .port_i (mixColumns_port_state_out_7_2_3[2:0]), //i
    .port_o (majority_5351_port_o                )  //o
  );
  Majority majority_5352 (
    .port_i (mixColumns_port_state_out_8_2_3[2:0]), //i
    .port_o (majority_5352_port_o                )  //o
  );
  Majority majority_5353 (
    .port_i (mixColumns_port_state_out_9_2_3[2:0]), //i
    .port_o (majority_5353_port_o                )  //o
  );
  Majority majority_5354 (
    .port_i (mixColumns_port_state_out_10_2_3[2:0]), //i
    .port_o (majority_5354_port_o                 )  //o
  );
  Majority majority_5355 (
    .port_i (mixColumns_port_state_out_11_2_3[2:0]), //i
    .port_o (majority_5355_port_o                 )  //o
  );
  Majority majority_5356 (
    .port_i (mixColumns_port_state_out_12_2_3[2:0]), //i
    .port_o (majority_5356_port_o                 )  //o
  );
  Majority majority_5357 (
    .port_i (mixColumns_port_state_out_13_2_3[2:0]), //i
    .port_o (majority_5357_port_o                 )  //o
  );
  Majority majority_5358 (
    .port_i (mixColumns_port_state_out_14_2_3[2:0]), //i
    .port_o (majority_5358_port_o                 )  //o
  );
  Majority majority_5359 (
    .port_i (mixColumns_port_state_out_15_2_3[2:0]), //i
    .port_o (majority_5359_port_o                 )  //o
  );
  Majority majority_5360 (
    .port_i (mixColumns_port_state_out_0_3_3[2:0]), //i
    .port_o (majority_5360_port_o                )  //o
  );
  Majority majority_5361 (
    .port_i (mixColumns_port_state_out_1_3_3[2:0]), //i
    .port_o (majority_5361_port_o                )  //o
  );
  Majority majority_5362 (
    .port_i (mixColumns_port_state_out_2_3_3[2:0]), //i
    .port_o (majority_5362_port_o                )  //o
  );
  Majority majority_5363 (
    .port_i (mixColumns_port_state_out_3_3_3[2:0]), //i
    .port_o (majority_5363_port_o                )  //o
  );
  Majority majority_5364 (
    .port_i (mixColumns_port_state_out_4_3_3[2:0]), //i
    .port_o (majority_5364_port_o                )  //o
  );
  Majority majority_5365 (
    .port_i (mixColumns_port_state_out_5_3_3[2:0]), //i
    .port_o (majority_5365_port_o                )  //o
  );
  Majority majority_5366 (
    .port_i (mixColumns_port_state_out_6_3_3[2:0]), //i
    .port_o (majority_5366_port_o                )  //o
  );
  Majority majority_5367 (
    .port_i (mixColumns_port_state_out_7_3_3[2:0]), //i
    .port_o (majority_5367_port_o                )  //o
  );
  Majority majority_5368 (
    .port_i (mixColumns_port_state_out_8_3_3[2:0]), //i
    .port_o (majority_5368_port_o                )  //o
  );
  Majority majority_5369 (
    .port_i (mixColumns_port_state_out_9_3_3[2:0]), //i
    .port_o (majority_5369_port_o                )  //o
  );
  Majority majority_5370 (
    .port_i (mixColumns_port_state_out_10_3_3[2:0]), //i
    .port_o (majority_5370_port_o                 )  //o
  );
  Majority majority_5371 (
    .port_i (mixColumns_port_state_out_11_3_3[2:0]), //i
    .port_o (majority_5371_port_o                 )  //o
  );
  Majority majority_5372 (
    .port_i (mixColumns_port_state_out_12_3_3[2:0]), //i
    .port_o (majority_5372_port_o                 )  //o
  );
  Majority majority_5373 (
    .port_i (mixColumns_port_state_out_13_3_3[2:0]), //i
    .port_o (majority_5373_port_o                 )  //o
  );
  Majority majority_5374 (
    .port_i (mixColumns_port_state_out_14_3_3[2:0]), //i
    .port_o (majority_5374_port_o                 )  //o
  );
  Majority majority_5375 (
    .port_i (mixColumns_port_state_out_15_3_3[2:0]), //i
    .port_o (majority_5375_port_o                 )  //o
  );
  Majority majority_5376 (
    .port_i (mixColumns_port_state_out_0_0_4[2:0]), //i
    .port_o (majority_5376_port_o                )  //o
  );
  Majority majority_5377 (
    .port_i (mixColumns_port_state_out_1_0_4[2:0]), //i
    .port_o (majority_5377_port_o                )  //o
  );
  Majority majority_5378 (
    .port_i (mixColumns_port_state_out_2_0_4[2:0]), //i
    .port_o (majority_5378_port_o                )  //o
  );
  Majority majority_5379 (
    .port_i (mixColumns_port_state_out_3_0_4[2:0]), //i
    .port_o (majority_5379_port_o                )  //o
  );
  Majority majority_5380 (
    .port_i (mixColumns_port_state_out_4_0_4[2:0]), //i
    .port_o (majority_5380_port_o                )  //o
  );
  Majority majority_5381 (
    .port_i (mixColumns_port_state_out_5_0_4[2:0]), //i
    .port_o (majority_5381_port_o                )  //o
  );
  Majority majority_5382 (
    .port_i (mixColumns_port_state_out_6_0_4[2:0]), //i
    .port_o (majority_5382_port_o                )  //o
  );
  Majority majority_5383 (
    .port_i (mixColumns_port_state_out_7_0_4[2:0]), //i
    .port_o (majority_5383_port_o                )  //o
  );
  Majority majority_5384 (
    .port_i (mixColumns_port_state_out_8_0_4[2:0]), //i
    .port_o (majority_5384_port_o                )  //o
  );
  Majority majority_5385 (
    .port_i (mixColumns_port_state_out_9_0_4[2:0]), //i
    .port_o (majority_5385_port_o                )  //o
  );
  Majority majority_5386 (
    .port_i (mixColumns_port_state_out_10_0_4[2:0]), //i
    .port_o (majority_5386_port_o                 )  //o
  );
  Majority majority_5387 (
    .port_i (mixColumns_port_state_out_11_0_4[2:0]), //i
    .port_o (majority_5387_port_o                 )  //o
  );
  Majority majority_5388 (
    .port_i (mixColumns_port_state_out_12_0_4[2:0]), //i
    .port_o (majority_5388_port_o                 )  //o
  );
  Majority majority_5389 (
    .port_i (mixColumns_port_state_out_13_0_4[2:0]), //i
    .port_o (majority_5389_port_o                 )  //o
  );
  Majority majority_5390 (
    .port_i (mixColumns_port_state_out_14_0_4[2:0]), //i
    .port_o (majority_5390_port_o                 )  //o
  );
  Majority majority_5391 (
    .port_i (mixColumns_port_state_out_15_0_4[2:0]), //i
    .port_o (majority_5391_port_o                 )  //o
  );
  Majority majority_5392 (
    .port_i (mixColumns_port_state_out_0_1_4[2:0]), //i
    .port_o (majority_5392_port_o                )  //o
  );
  Majority majority_5393 (
    .port_i (mixColumns_port_state_out_1_1_4[2:0]), //i
    .port_o (majority_5393_port_o                )  //o
  );
  Majority majority_5394 (
    .port_i (mixColumns_port_state_out_2_1_4[2:0]), //i
    .port_o (majority_5394_port_o                )  //o
  );
  Majority majority_5395 (
    .port_i (mixColumns_port_state_out_3_1_4[2:0]), //i
    .port_o (majority_5395_port_o                )  //o
  );
  Majority majority_5396 (
    .port_i (mixColumns_port_state_out_4_1_4[2:0]), //i
    .port_o (majority_5396_port_o                )  //o
  );
  Majority majority_5397 (
    .port_i (mixColumns_port_state_out_5_1_4[2:0]), //i
    .port_o (majority_5397_port_o                )  //o
  );
  Majority majority_5398 (
    .port_i (mixColumns_port_state_out_6_1_4[2:0]), //i
    .port_o (majority_5398_port_o                )  //o
  );
  Majority majority_5399 (
    .port_i (mixColumns_port_state_out_7_1_4[2:0]), //i
    .port_o (majority_5399_port_o                )  //o
  );
  Majority majority_5400 (
    .port_i (mixColumns_port_state_out_8_1_4[2:0]), //i
    .port_o (majority_5400_port_o                )  //o
  );
  Majority majority_5401 (
    .port_i (mixColumns_port_state_out_9_1_4[2:0]), //i
    .port_o (majority_5401_port_o                )  //o
  );
  Majority majority_5402 (
    .port_i (mixColumns_port_state_out_10_1_4[2:0]), //i
    .port_o (majority_5402_port_o                 )  //o
  );
  Majority majority_5403 (
    .port_i (mixColumns_port_state_out_11_1_4[2:0]), //i
    .port_o (majority_5403_port_o                 )  //o
  );
  Majority majority_5404 (
    .port_i (mixColumns_port_state_out_12_1_4[2:0]), //i
    .port_o (majority_5404_port_o                 )  //o
  );
  Majority majority_5405 (
    .port_i (mixColumns_port_state_out_13_1_4[2:0]), //i
    .port_o (majority_5405_port_o                 )  //o
  );
  Majority majority_5406 (
    .port_i (mixColumns_port_state_out_14_1_4[2:0]), //i
    .port_o (majority_5406_port_o                 )  //o
  );
  Majority majority_5407 (
    .port_i (mixColumns_port_state_out_15_1_4[2:0]), //i
    .port_o (majority_5407_port_o                 )  //o
  );
  Majority majority_5408 (
    .port_i (mixColumns_port_state_out_0_2_4[2:0]), //i
    .port_o (majority_5408_port_o                )  //o
  );
  Majority majority_5409 (
    .port_i (mixColumns_port_state_out_1_2_4[2:0]), //i
    .port_o (majority_5409_port_o                )  //o
  );
  Majority majority_5410 (
    .port_i (mixColumns_port_state_out_2_2_4[2:0]), //i
    .port_o (majority_5410_port_o                )  //o
  );
  Majority majority_5411 (
    .port_i (mixColumns_port_state_out_3_2_4[2:0]), //i
    .port_o (majority_5411_port_o                )  //o
  );
  Majority majority_5412 (
    .port_i (mixColumns_port_state_out_4_2_4[2:0]), //i
    .port_o (majority_5412_port_o                )  //o
  );
  Majority majority_5413 (
    .port_i (mixColumns_port_state_out_5_2_4[2:0]), //i
    .port_o (majority_5413_port_o                )  //o
  );
  Majority majority_5414 (
    .port_i (mixColumns_port_state_out_6_2_4[2:0]), //i
    .port_o (majority_5414_port_o                )  //o
  );
  Majority majority_5415 (
    .port_i (mixColumns_port_state_out_7_2_4[2:0]), //i
    .port_o (majority_5415_port_o                )  //o
  );
  Majority majority_5416 (
    .port_i (mixColumns_port_state_out_8_2_4[2:0]), //i
    .port_o (majority_5416_port_o                )  //o
  );
  Majority majority_5417 (
    .port_i (mixColumns_port_state_out_9_2_4[2:0]), //i
    .port_o (majority_5417_port_o                )  //o
  );
  Majority majority_5418 (
    .port_i (mixColumns_port_state_out_10_2_4[2:0]), //i
    .port_o (majority_5418_port_o                 )  //o
  );
  Majority majority_5419 (
    .port_i (mixColumns_port_state_out_11_2_4[2:0]), //i
    .port_o (majority_5419_port_o                 )  //o
  );
  Majority majority_5420 (
    .port_i (mixColumns_port_state_out_12_2_4[2:0]), //i
    .port_o (majority_5420_port_o                 )  //o
  );
  Majority majority_5421 (
    .port_i (mixColumns_port_state_out_13_2_4[2:0]), //i
    .port_o (majority_5421_port_o                 )  //o
  );
  Majority majority_5422 (
    .port_i (mixColumns_port_state_out_14_2_4[2:0]), //i
    .port_o (majority_5422_port_o                 )  //o
  );
  Majority majority_5423 (
    .port_i (mixColumns_port_state_out_15_2_4[2:0]), //i
    .port_o (majority_5423_port_o                 )  //o
  );
  Majority majority_5424 (
    .port_i (mixColumns_port_state_out_0_3_4[2:0]), //i
    .port_o (majority_5424_port_o                )  //o
  );
  Majority majority_5425 (
    .port_i (mixColumns_port_state_out_1_3_4[2:0]), //i
    .port_o (majority_5425_port_o                )  //o
  );
  Majority majority_5426 (
    .port_i (mixColumns_port_state_out_2_3_4[2:0]), //i
    .port_o (majority_5426_port_o                )  //o
  );
  Majority majority_5427 (
    .port_i (mixColumns_port_state_out_3_3_4[2:0]), //i
    .port_o (majority_5427_port_o                )  //o
  );
  Majority majority_5428 (
    .port_i (mixColumns_port_state_out_4_3_4[2:0]), //i
    .port_o (majority_5428_port_o                )  //o
  );
  Majority majority_5429 (
    .port_i (mixColumns_port_state_out_5_3_4[2:0]), //i
    .port_o (majority_5429_port_o                )  //o
  );
  Majority majority_5430 (
    .port_i (mixColumns_port_state_out_6_3_4[2:0]), //i
    .port_o (majority_5430_port_o                )  //o
  );
  Majority majority_5431 (
    .port_i (mixColumns_port_state_out_7_3_4[2:0]), //i
    .port_o (majority_5431_port_o                )  //o
  );
  Majority majority_5432 (
    .port_i (mixColumns_port_state_out_8_3_4[2:0]), //i
    .port_o (majority_5432_port_o                )  //o
  );
  Majority majority_5433 (
    .port_i (mixColumns_port_state_out_9_3_4[2:0]), //i
    .port_o (majority_5433_port_o                )  //o
  );
  Majority majority_5434 (
    .port_i (mixColumns_port_state_out_10_3_4[2:0]), //i
    .port_o (majority_5434_port_o                 )  //o
  );
  Majority majority_5435 (
    .port_i (mixColumns_port_state_out_11_3_4[2:0]), //i
    .port_o (majority_5435_port_o                 )  //o
  );
  Majority majority_5436 (
    .port_i (mixColumns_port_state_out_12_3_4[2:0]), //i
    .port_o (majority_5436_port_o                 )  //o
  );
  Majority majority_5437 (
    .port_i (mixColumns_port_state_out_13_3_4[2:0]), //i
    .port_o (majority_5437_port_o                 )  //o
  );
  Majority majority_5438 (
    .port_i (mixColumns_port_state_out_14_3_4[2:0]), //i
    .port_o (majority_5438_port_o                 )  //o
  );
  Majority majority_5439 (
    .port_i (mixColumns_port_state_out_15_3_4[2:0]), //i
    .port_o (majority_5439_port_o                 )  //o
  );
  Majority majority_5440 (
    .port_i (mixColumns_port_state_out_0_0_5[2:0]), //i
    .port_o (majority_5440_port_o                )  //o
  );
  Majority majority_5441 (
    .port_i (mixColumns_port_state_out_1_0_5[2:0]), //i
    .port_o (majority_5441_port_o                )  //o
  );
  Majority majority_5442 (
    .port_i (mixColumns_port_state_out_2_0_5[2:0]), //i
    .port_o (majority_5442_port_o                )  //o
  );
  Majority majority_5443 (
    .port_i (mixColumns_port_state_out_3_0_5[2:0]), //i
    .port_o (majority_5443_port_o                )  //o
  );
  Majority majority_5444 (
    .port_i (mixColumns_port_state_out_4_0_5[2:0]), //i
    .port_o (majority_5444_port_o                )  //o
  );
  Majority majority_5445 (
    .port_i (mixColumns_port_state_out_5_0_5[2:0]), //i
    .port_o (majority_5445_port_o                )  //o
  );
  Majority majority_5446 (
    .port_i (mixColumns_port_state_out_6_0_5[2:0]), //i
    .port_o (majority_5446_port_o                )  //o
  );
  Majority majority_5447 (
    .port_i (mixColumns_port_state_out_7_0_5[2:0]), //i
    .port_o (majority_5447_port_o                )  //o
  );
  Majority majority_5448 (
    .port_i (mixColumns_port_state_out_8_0_5[2:0]), //i
    .port_o (majority_5448_port_o                )  //o
  );
  Majority majority_5449 (
    .port_i (mixColumns_port_state_out_9_0_5[2:0]), //i
    .port_o (majority_5449_port_o                )  //o
  );
  Majority majority_5450 (
    .port_i (mixColumns_port_state_out_10_0_5[2:0]), //i
    .port_o (majority_5450_port_o                 )  //o
  );
  Majority majority_5451 (
    .port_i (mixColumns_port_state_out_11_0_5[2:0]), //i
    .port_o (majority_5451_port_o                 )  //o
  );
  Majority majority_5452 (
    .port_i (mixColumns_port_state_out_12_0_5[2:0]), //i
    .port_o (majority_5452_port_o                 )  //o
  );
  Majority majority_5453 (
    .port_i (mixColumns_port_state_out_13_0_5[2:0]), //i
    .port_o (majority_5453_port_o                 )  //o
  );
  Majority majority_5454 (
    .port_i (mixColumns_port_state_out_14_0_5[2:0]), //i
    .port_o (majority_5454_port_o                 )  //o
  );
  Majority majority_5455 (
    .port_i (mixColumns_port_state_out_15_0_5[2:0]), //i
    .port_o (majority_5455_port_o                 )  //o
  );
  Majority majority_5456 (
    .port_i (mixColumns_port_state_out_0_1_5[2:0]), //i
    .port_o (majority_5456_port_o                )  //o
  );
  Majority majority_5457 (
    .port_i (mixColumns_port_state_out_1_1_5[2:0]), //i
    .port_o (majority_5457_port_o                )  //o
  );
  Majority majority_5458 (
    .port_i (mixColumns_port_state_out_2_1_5[2:0]), //i
    .port_o (majority_5458_port_o                )  //o
  );
  Majority majority_5459 (
    .port_i (mixColumns_port_state_out_3_1_5[2:0]), //i
    .port_o (majority_5459_port_o                )  //o
  );
  Majority majority_5460 (
    .port_i (mixColumns_port_state_out_4_1_5[2:0]), //i
    .port_o (majority_5460_port_o                )  //o
  );
  Majority majority_5461 (
    .port_i (mixColumns_port_state_out_5_1_5[2:0]), //i
    .port_o (majority_5461_port_o                )  //o
  );
  Majority majority_5462 (
    .port_i (mixColumns_port_state_out_6_1_5[2:0]), //i
    .port_o (majority_5462_port_o                )  //o
  );
  Majority majority_5463 (
    .port_i (mixColumns_port_state_out_7_1_5[2:0]), //i
    .port_o (majority_5463_port_o                )  //o
  );
  Majority majority_5464 (
    .port_i (mixColumns_port_state_out_8_1_5[2:0]), //i
    .port_o (majority_5464_port_o                )  //o
  );
  Majority majority_5465 (
    .port_i (mixColumns_port_state_out_9_1_5[2:0]), //i
    .port_o (majority_5465_port_o                )  //o
  );
  Majority majority_5466 (
    .port_i (mixColumns_port_state_out_10_1_5[2:0]), //i
    .port_o (majority_5466_port_o                 )  //o
  );
  Majority majority_5467 (
    .port_i (mixColumns_port_state_out_11_1_5[2:0]), //i
    .port_o (majority_5467_port_o                 )  //o
  );
  Majority majority_5468 (
    .port_i (mixColumns_port_state_out_12_1_5[2:0]), //i
    .port_o (majority_5468_port_o                 )  //o
  );
  Majority majority_5469 (
    .port_i (mixColumns_port_state_out_13_1_5[2:0]), //i
    .port_o (majority_5469_port_o                 )  //o
  );
  Majority majority_5470 (
    .port_i (mixColumns_port_state_out_14_1_5[2:0]), //i
    .port_o (majority_5470_port_o                 )  //o
  );
  Majority majority_5471 (
    .port_i (mixColumns_port_state_out_15_1_5[2:0]), //i
    .port_o (majority_5471_port_o                 )  //o
  );
  Majority majority_5472 (
    .port_i (mixColumns_port_state_out_0_2_5[2:0]), //i
    .port_o (majority_5472_port_o                )  //o
  );
  Majority majority_5473 (
    .port_i (mixColumns_port_state_out_1_2_5[2:0]), //i
    .port_o (majority_5473_port_o                )  //o
  );
  Majority majority_5474 (
    .port_i (mixColumns_port_state_out_2_2_5[2:0]), //i
    .port_o (majority_5474_port_o                )  //o
  );
  Majority majority_5475 (
    .port_i (mixColumns_port_state_out_3_2_5[2:0]), //i
    .port_o (majority_5475_port_o                )  //o
  );
  Majority majority_5476 (
    .port_i (mixColumns_port_state_out_4_2_5[2:0]), //i
    .port_o (majority_5476_port_o                )  //o
  );
  Majority majority_5477 (
    .port_i (mixColumns_port_state_out_5_2_5[2:0]), //i
    .port_o (majority_5477_port_o                )  //o
  );
  Majority majority_5478 (
    .port_i (mixColumns_port_state_out_6_2_5[2:0]), //i
    .port_o (majority_5478_port_o                )  //o
  );
  Majority majority_5479 (
    .port_i (mixColumns_port_state_out_7_2_5[2:0]), //i
    .port_o (majority_5479_port_o                )  //o
  );
  Majority majority_5480 (
    .port_i (mixColumns_port_state_out_8_2_5[2:0]), //i
    .port_o (majority_5480_port_o                )  //o
  );
  Majority majority_5481 (
    .port_i (mixColumns_port_state_out_9_2_5[2:0]), //i
    .port_o (majority_5481_port_o                )  //o
  );
  Majority majority_5482 (
    .port_i (mixColumns_port_state_out_10_2_5[2:0]), //i
    .port_o (majority_5482_port_o                 )  //o
  );
  Majority majority_5483 (
    .port_i (mixColumns_port_state_out_11_2_5[2:0]), //i
    .port_o (majority_5483_port_o                 )  //o
  );
  Majority majority_5484 (
    .port_i (mixColumns_port_state_out_12_2_5[2:0]), //i
    .port_o (majority_5484_port_o                 )  //o
  );
  Majority majority_5485 (
    .port_i (mixColumns_port_state_out_13_2_5[2:0]), //i
    .port_o (majority_5485_port_o                 )  //o
  );
  Majority majority_5486 (
    .port_i (mixColumns_port_state_out_14_2_5[2:0]), //i
    .port_o (majority_5486_port_o                 )  //o
  );
  Majority majority_5487 (
    .port_i (mixColumns_port_state_out_15_2_5[2:0]), //i
    .port_o (majority_5487_port_o                 )  //o
  );
  Majority majority_5488 (
    .port_i (mixColumns_port_state_out_0_3_5[2:0]), //i
    .port_o (majority_5488_port_o                )  //o
  );
  Majority majority_5489 (
    .port_i (mixColumns_port_state_out_1_3_5[2:0]), //i
    .port_o (majority_5489_port_o                )  //o
  );
  Majority majority_5490 (
    .port_i (mixColumns_port_state_out_2_3_5[2:0]), //i
    .port_o (majority_5490_port_o                )  //o
  );
  Majority majority_5491 (
    .port_i (mixColumns_port_state_out_3_3_5[2:0]), //i
    .port_o (majority_5491_port_o                )  //o
  );
  Majority majority_5492 (
    .port_i (mixColumns_port_state_out_4_3_5[2:0]), //i
    .port_o (majority_5492_port_o                )  //o
  );
  Majority majority_5493 (
    .port_i (mixColumns_port_state_out_5_3_5[2:0]), //i
    .port_o (majority_5493_port_o                )  //o
  );
  Majority majority_5494 (
    .port_i (mixColumns_port_state_out_6_3_5[2:0]), //i
    .port_o (majority_5494_port_o                )  //o
  );
  Majority majority_5495 (
    .port_i (mixColumns_port_state_out_7_3_5[2:0]), //i
    .port_o (majority_5495_port_o                )  //o
  );
  Majority majority_5496 (
    .port_i (mixColumns_port_state_out_8_3_5[2:0]), //i
    .port_o (majority_5496_port_o                )  //o
  );
  Majority majority_5497 (
    .port_i (mixColumns_port_state_out_9_3_5[2:0]), //i
    .port_o (majority_5497_port_o                )  //o
  );
  Majority majority_5498 (
    .port_i (mixColumns_port_state_out_10_3_5[2:0]), //i
    .port_o (majority_5498_port_o                 )  //o
  );
  Majority majority_5499 (
    .port_i (mixColumns_port_state_out_11_3_5[2:0]), //i
    .port_o (majority_5499_port_o                 )  //o
  );
  Majority majority_5500 (
    .port_i (mixColumns_port_state_out_12_3_5[2:0]), //i
    .port_o (majority_5500_port_o                 )  //o
  );
  Majority majority_5501 (
    .port_i (mixColumns_port_state_out_13_3_5[2:0]), //i
    .port_o (majority_5501_port_o                 )  //o
  );
  Majority majority_5502 (
    .port_i (mixColumns_port_state_out_14_3_5[2:0]), //i
    .port_o (majority_5502_port_o                 )  //o
  );
  Majority majority_5503 (
    .port_i (mixColumns_port_state_out_15_3_5[2:0]), //i
    .port_o (majority_5503_port_o                 )  //o
  );
  Majority majority_5504 (
    .port_i (mixColumns_port_state_out_0_0_6[2:0]), //i
    .port_o (majority_5504_port_o                )  //o
  );
  Majority majority_5505 (
    .port_i (mixColumns_port_state_out_1_0_6[2:0]), //i
    .port_o (majority_5505_port_o                )  //o
  );
  Majority majority_5506 (
    .port_i (mixColumns_port_state_out_2_0_6[2:0]), //i
    .port_o (majority_5506_port_o                )  //o
  );
  Majority majority_5507 (
    .port_i (mixColumns_port_state_out_3_0_6[2:0]), //i
    .port_o (majority_5507_port_o                )  //o
  );
  Majority majority_5508 (
    .port_i (mixColumns_port_state_out_4_0_6[2:0]), //i
    .port_o (majority_5508_port_o                )  //o
  );
  Majority majority_5509 (
    .port_i (mixColumns_port_state_out_5_0_6[2:0]), //i
    .port_o (majority_5509_port_o                )  //o
  );
  Majority majority_5510 (
    .port_i (mixColumns_port_state_out_6_0_6[2:0]), //i
    .port_o (majority_5510_port_o                )  //o
  );
  Majority majority_5511 (
    .port_i (mixColumns_port_state_out_7_0_6[2:0]), //i
    .port_o (majority_5511_port_o                )  //o
  );
  Majority majority_5512 (
    .port_i (mixColumns_port_state_out_8_0_6[2:0]), //i
    .port_o (majority_5512_port_o                )  //o
  );
  Majority majority_5513 (
    .port_i (mixColumns_port_state_out_9_0_6[2:0]), //i
    .port_o (majority_5513_port_o                )  //o
  );
  Majority majority_5514 (
    .port_i (mixColumns_port_state_out_10_0_6[2:0]), //i
    .port_o (majority_5514_port_o                 )  //o
  );
  Majority majority_5515 (
    .port_i (mixColumns_port_state_out_11_0_6[2:0]), //i
    .port_o (majority_5515_port_o                 )  //o
  );
  Majority majority_5516 (
    .port_i (mixColumns_port_state_out_12_0_6[2:0]), //i
    .port_o (majority_5516_port_o                 )  //o
  );
  Majority majority_5517 (
    .port_i (mixColumns_port_state_out_13_0_6[2:0]), //i
    .port_o (majority_5517_port_o                 )  //o
  );
  Majority majority_5518 (
    .port_i (mixColumns_port_state_out_14_0_6[2:0]), //i
    .port_o (majority_5518_port_o                 )  //o
  );
  Majority majority_5519 (
    .port_i (mixColumns_port_state_out_15_0_6[2:0]), //i
    .port_o (majority_5519_port_o                 )  //o
  );
  Majority majority_5520 (
    .port_i (mixColumns_port_state_out_0_1_6[2:0]), //i
    .port_o (majority_5520_port_o                )  //o
  );
  Majority majority_5521 (
    .port_i (mixColumns_port_state_out_1_1_6[2:0]), //i
    .port_o (majority_5521_port_o                )  //o
  );
  Majority majority_5522 (
    .port_i (mixColumns_port_state_out_2_1_6[2:0]), //i
    .port_o (majority_5522_port_o                )  //o
  );
  Majority majority_5523 (
    .port_i (mixColumns_port_state_out_3_1_6[2:0]), //i
    .port_o (majority_5523_port_o                )  //o
  );
  Majority majority_5524 (
    .port_i (mixColumns_port_state_out_4_1_6[2:0]), //i
    .port_o (majority_5524_port_o                )  //o
  );
  Majority majority_5525 (
    .port_i (mixColumns_port_state_out_5_1_6[2:0]), //i
    .port_o (majority_5525_port_o                )  //o
  );
  Majority majority_5526 (
    .port_i (mixColumns_port_state_out_6_1_6[2:0]), //i
    .port_o (majority_5526_port_o                )  //o
  );
  Majority majority_5527 (
    .port_i (mixColumns_port_state_out_7_1_6[2:0]), //i
    .port_o (majority_5527_port_o                )  //o
  );
  Majority majority_5528 (
    .port_i (mixColumns_port_state_out_8_1_6[2:0]), //i
    .port_o (majority_5528_port_o                )  //o
  );
  Majority majority_5529 (
    .port_i (mixColumns_port_state_out_9_1_6[2:0]), //i
    .port_o (majority_5529_port_o                )  //o
  );
  Majority majority_5530 (
    .port_i (mixColumns_port_state_out_10_1_6[2:0]), //i
    .port_o (majority_5530_port_o                 )  //o
  );
  Majority majority_5531 (
    .port_i (mixColumns_port_state_out_11_1_6[2:0]), //i
    .port_o (majority_5531_port_o                 )  //o
  );
  Majority majority_5532 (
    .port_i (mixColumns_port_state_out_12_1_6[2:0]), //i
    .port_o (majority_5532_port_o                 )  //o
  );
  Majority majority_5533 (
    .port_i (mixColumns_port_state_out_13_1_6[2:0]), //i
    .port_o (majority_5533_port_o                 )  //o
  );
  Majority majority_5534 (
    .port_i (mixColumns_port_state_out_14_1_6[2:0]), //i
    .port_o (majority_5534_port_o                 )  //o
  );
  Majority majority_5535 (
    .port_i (mixColumns_port_state_out_15_1_6[2:0]), //i
    .port_o (majority_5535_port_o                 )  //o
  );
  Majority majority_5536 (
    .port_i (mixColumns_port_state_out_0_2_6[2:0]), //i
    .port_o (majority_5536_port_o                )  //o
  );
  Majority majority_5537 (
    .port_i (mixColumns_port_state_out_1_2_6[2:0]), //i
    .port_o (majority_5537_port_o                )  //o
  );
  Majority majority_5538 (
    .port_i (mixColumns_port_state_out_2_2_6[2:0]), //i
    .port_o (majority_5538_port_o                )  //o
  );
  Majority majority_5539 (
    .port_i (mixColumns_port_state_out_3_2_6[2:0]), //i
    .port_o (majority_5539_port_o                )  //o
  );
  Majority majority_5540 (
    .port_i (mixColumns_port_state_out_4_2_6[2:0]), //i
    .port_o (majority_5540_port_o                )  //o
  );
  Majority majority_5541 (
    .port_i (mixColumns_port_state_out_5_2_6[2:0]), //i
    .port_o (majority_5541_port_o                )  //o
  );
  Majority majority_5542 (
    .port_i (mixColumns_port_state_out_6_2_6[2:0]), //i
    .port_o (majority_5542_port_o                )  //o
  );
  Majority majority_5543 (
    .port_i (mixColumns_port_state_out_7_2_6[2:0]), //i
    .port_o (majority_5543_port_o                )  //o
  );
  Majority majority_5544 (
    .port_i (mixColumns_port_state_out_8_2_6[2:0]), //i
    .port_o (majority_5544_port_o                )  //o
  );
  Majority majority_5545 (
    .port_i (mixColumns_port_state_out_9_2_6[2:0]), //i
    .port_o (majority_5545_port_o                )  //o
  );
  Majority majority_5546 (
    .port_i (mixColumns_port_state_out_10_2_6[2:0]), //i
    .port_o (majority_5546_port_o                 )  //o
  );
  Majority majority_5547 (
    .port_i (mixColumns_port_state_out_11_2_6[2:0]), //i
    .port_o (majority_5547_port_o                 )  //o
  );
  Majority majority_5548 (
    .port_i (mixColumns_port_state_out_12_2_6[2:0]), //i
    .port_o (majority_5548_port_o                 )  //o
  );
  Majority majority_5549 (
    .port_i (mixColumns_port_state_out_13_2_6[2:0]), //i
    .port_o (majority_5549_port_o                 )  //o
  );
  Majority majority_5550 (
    .port_i (mixColumns_port_state_out_14_2_6[2:0]), //i
    .port_o (majority_5550_port_o                 )  //o
  );
  Majority majority_5551 (
    .port_i (mixColumns_port_state_out_15_2_6[2:0]), //i
    .port_o (majority_5551_port_o                 )  //o
  );
  Majority majority_5552 (
    .port_i (mixColumns_port_state_out_0_3_6[2:0]), //i
    .port_o (majority_5552_port_o                )  //o
  );
  Majority majority_5553 (
    .port_i (mixColumns_port_state_out_1_3_6[2:0]), //i
    .port_o (majority_5553_port_o                )  //o
  );
  Majority majority_5554 (
    .port_i (mixColumns_port_state_out_2_3_6[2:0]), //i
    .port_o (majority_5554_port_o                )  //o
  );
  Majority majority_5555 (
    .port_i (mixColumns_port_state_out_3_3_6[2:0]), //i
    .port_o (majority_5555_port_o                )  //o
  );
  Majority majority_5556 (
    .port_i (mixColumns_port_state_out_4_3_6[2:0]), //i
    .port_o (majority_5556_port_o                )  //o
  );
  Majority majority_5557 (
    .port_i (mixColumns_port_state_out_5_3_6[2:0]), //i
    .port_o (majority_5557_port_o                )  //o
  );
  Majority majority_5558 (
    .port_i (mixColumns_port_state_out_6_3_6[2:0]), //i
    .port_o (majority_5558_port_o                )  //o
  );
  Majority majority_5559 (
    .port_i (mixColumns_port_state_out_7_3_6[2:0]), //i
    .port_o (majority_5559_port_o                )  //o
  );
  Majority majority_5560 (
    .port_i (mixColumns_port_state_out_8_3_6[2:0]), //i
    .port_o (majority_5560_port_o                )  //o
  );
  Majority majority_5561 (
    .port_i (mixColumns_port_state_out_9_3_6[2:0]), //i
    .port_o (majority_5561_port_o                )  //o
  );
  Majority majority_5562 (
    .port_i (mixColumns_port_state_out_10_3_6[2:0]), //i
    .port_o (majority_5562_port_o                 )  //o
  );
  Majority majority_5563 (
    .port_i (mixColumns_port_state_out_11_3_6[2:0]), //i
    .port_o (majority_5563_port_o                 )  //o
  );
  Majority majority_5564 (
    .port_i (mixColumns_port_state_out_12_3_6[2:0]), //i
    .port_o (majority_5564_port_o                 )  //o
  );
  Majority majority_5565 (
    .port_i (mixColumns_port_state_out_13_3_6[2:0]), //i
    .port_o (majority_5565_port_o                 )  //o
  );
  Majority majority_5566 (
    .port_i (mixColumns_port_state_out_14_3_6[2:0]), //i
    .port_o (majority_5566_port_o                 )  //o
  );
  Majority majority_5567 (
    .port_i (mixColumns_port_state_out_15_3_6[2:0]), //i
    .port_o (majority_5567_port_o                 )  //o
  );
  Majority majority_5568 (
    .port_i (mixColumns_port_state_out_0_0_7[2:0]), //i
    .port_o (majority_5568_port_o                )  //o
  );
  Majority majority_5569 (
    .port_i (mixColumns_port_state_out_1_0_7[2:0]), //i
    .port_o (majority_5569_port_o                )  //o
  );
  Majority majority_5570 (
    .port_i (mixColumns_port_state_out_2_0_7[2:0]), //i
    .port_o (majority_5570_port_o                )  //o
  );
  Majority majority_5571 (
    .port_i (mixColumns_port_state_out_3_0_7[2:0]), //i
    .port_o (majority_5571_port_o                )  //o
  );
  Majority majority_5572 (
    .port_i (mixColumns_port_state_out_4_0_7[2:0]), //i
    .port_o (majority_5572_port_o                )  //o
  );
  Majority majority_5573 (
    .port_i (mixColumns_port_state_out_5_0_7[2:0]), //i
    .port_o (majority_5573_port_o                )  //o
  );
  Majority majority_5574 (
    .port_i (mixColumns_port_state_out_6_0_7[2:0]), //i
    .port_o (majority_5574_port_o                )  //o
  );
  Majority majority_5575 (
    .port_i (mixColumns_port_state_out_7_0_7[2:0]), //i
    .port_o (majority_5575_port_o                )  //o
  );
  Majority majority_5576 (
    .port_i (mixColumns_port_state_out_8_0_7[2:0]), //i
    .port_o (majority_5576_port_o                )  //o
  );
  Majority majority_5577 (
    .port_i (mixColumns_port_state_out_9_0_7[2:0]), //i
    .port_o (majority_5577_port_o                )  //o
  );
  Majority majority_5578 (
    .port_i (mixColumns_port_state_out_10_0_7[2:0]), //i
    .port_o (majority_5578_port_o                 )  //o
  );
  Majority majority_5579 (
    .port_i (mixColumns_port_state_out_11_0_7[2:0]), //i
    .port_o (majority_5579_port_o                 )  //o
  );
  Majority majority_5580 (
    .port_i (mixColumns_port_state_out_12_0_7[2:0]), //i
    .port_o (majority_5580_port_o                 )  //o
  );
  Majority majority_5581 (
    .port_i (mixColumns_port_state_out_13_0_7[2:0]), //i
    .port_o (majority_5581_port_o                 )  //o
  );
  Majority majority_5582 (
    .port_i (mixColumns_port_state_out_14_0_7[2:0]), //i
    .port_o (majority_5582_port_o                 )  //o
  );
  Majority majority_5583 (
    .port_i (mixColumns_port_state_out_15_0_7[2:0]), //i
    .port_o (majority_5583_port_o                 )  //o
  );
  Majority majority_5584 (
    .port_i (mixColumns_port_state_out_0_1_7[2:0]), //i
    .port_o (majority_5584_port_o                )  //o
  );
  Majority majority_5585 (
    .port_i (mixColumns_port_state_out_1_1_7[2:0]), //i
    .port_o (majority_5585_port_o                )  //o
  );
  Majority majority_5586 (
    .port_i (mixColumns_port_state_out_2_1_7[2:0]), //i
    .port_o (majority_5586_port_o                )  //o
  );
  Majority majority_5587 (
    .port_i (mixColumns_port_state_out_3_1_7[2:0]), //i
    .port_o (majority_5587_port_o                )  //o
  );
  Majority majority_5588 (
    .port_i (mixColumns_port_state_out_4_1_7[2:0]), //i
    .port_o (majority_5588_port_o                )  //o
  );
  Majority majority_5589 (
    .port_i (mixColumns_port_state_out_5_1_7[2:0]), //i
    .port_o (majority_5589_port_o                )  //o
  );
  Majority majority_5590 (
    .port_i (mixColumns_port_state_out_6_1_7[2:0]), //i
    .port_o (majority_5590_port_o                )  //o
  );
  Majority majority_5591 (
    .port_i (mixColumns_port_state_out_7_1_7[2:0]), //i
    .port_o (majority_5591_port_o                )  //o
  );
  Majority majority_5592 (
    .port_i (mixColumns_port_state_out_8_1_7[2:0]), //i
    .port_o (majority_5592_port_o                )  //o
  );
  Majority majority_5593 (
    .port_i (mixColumns_port_state_out_9_1_7[2:0]), //i
    .port_o (majority_5593_port_o                )  //o
  );
  Majority majority_5594 (
    .port_i (mixColumns_port_state_out_10_1_7[2:0]), //i
    .port_o (majority_5594_port_o                 )  //o
  );
  Majority majority_5595 (
    .port_i (mixColumns_port_state_out_11_1_7[2:0]), //i
    .port_o (majority_5595_port_o                 )  //o
  );
  Majority majority_5596 (
    .port_i (mixColumns_port_state_out_12_1_7[2:0]), //i
    .port_o (majority_5596_port_o                 )  //o
  );
  Majority majority_5597 (
    .port_i (mixColumns_port_state_out_13_1_7[2:0]), //i
    .port_o (majority_5597_port_o                 )  //o
  );
  Majority majority_5598 (
    .port_i (mixColumns_port_state_out_14_1_7[2:0]), //i
    .port_o (majority_5598_port_o                 )  //o
  );
  Majority majority_5599 (
    .port_i (mixColumns_port_state_out_15_1_7[2:0]), //i
    .port_o (majority_5599_port_o                 )  //o
  );
  Majority majority_5600 (
    .port_i (mixColumns_port_state_out_0_2_7[2:0]), //i
    .port_o (majority_5600_port_o                )  //o
  );
  Majority majority_5601 (
    .port_i (mixColumns_port_state_out_1_2_7[2:0]), //i
    .port_o (majority_5601_port_o                )  //o
  );
  Majority majority_5602 (
    .port_i (mixColumns_port_state_out_2_2_7[2:0]), //i
    .port_o (majority_5602_port_o                )  //o
  );
  Majority majority_5603 (
    .port_i (mixColumns_port_state_out_3_2_7[2:0]), //i
    .port_o (majority_5603_port_o                )  //o
  );
  Majority majority_5604 (
    .port_i (mixColumns_port_state_out_4_2_7[2:0]), //i
    .port_o (majority_5604_port_o                )  //o
  );
  Majority majority_5605 (
    .port_i (mixColumns_port_state_out_5_2_7[2:0]), //i
    .port_o (majority_5605_port_o                )  //o
  );
  Majority majority_5606 (
    .port_i (mixColumns_port_state_out_6_2_7[2:0]), //i
    .port_o (majority_5606_port_o                )  //o
  );
  Majority majority_5607 (
    .port_i (mixColumns_port_state_out_7_2_7[2:0]), //i
    .port_o (majority_5607_port_o                )  //o
  );
  Majority majority_5608 (
    .port_i (mixColumns_port_state_out_8_2_7[2:0]), //i
    .port_o (majority_5608_port_o                )  //o
  );
  Majority majority_5609 (
    .port_i (mixColumns_port_state_out_9_2_7[2:0]), //i
    .port_o (majority_5609_port_o                )  //o
  );
  Majority majority_5610 (
    .port_i (mixColumns_port_state_out_10_2_7[2:0]), //i
    .port_o (majority_5610_port_o                 )  //o
  );
  Majority majority_5611 (
    .port_i (mixColumns_port_state_out_11_2_7[2:0]), //i
    .port_o (majority_5611_port_o                 )  //o
  );
  Majority majority_5612 (
    .port_i (mixColumns_port_state_out_12_2_7[2:0]), //i
    .port_o (majority_5612_port_o                 )  //o
  );
  Majority majority_5613 (
    .port_i (mixColumns_port_state_out_13_2_7[2:0]), //i
    .port_o (majority_5613_port_o                 )  //o
  );
  Majority majority_5614 (
    .port_i (mixColumns_port_state_out_14_2_7[2:0]), //i
    .port_o (majority_5614_port_o                 )  //o
  );
  Majority majority_5615 (
    .port_i (mixColumns_port_state_out_15_2_7[2:0]), //i
    .port_o (majority_5615_port_o                 )  //o
  );
  Majority majority_5616 (
    .port_i (mixColumns_port_state_out_0_3_7[2:0]), //i
    .port_o (majority_5616_port_o                )  //o
  );
  Majority majority_5617 (
    .port_i (mixColumns_port_state_out_1_3_7[2:0]), //i
    .port_o (majority_5617_port_o                )  //o
  );
  Majority majority_5618 (
    .port_i (mixColumns_port_state_out_2_3_7[2:0]), //i
    .port_o (majority_5618_port_o                )  //o
  );
  Majority majority_5619 (
    .port_i (mixColumns_port_state_out_3_3_7[2:0]), //i
    .port_o (majority_5619_port_o                )  //o
  );
  Majority majority_5620 (
    .port_i (mixColumns_port_state_out_4_3_7[2:0]), //i
    .port_o (majority_5620_port_o                )  //o
  );
  Majority majority_5621 (
    .port_i (mixColumns_port_state_out_5_3_7[2:0]), //i
    .port_o (majority_5621_port_o                )  //o
  );
  Majority majority_5622 (
    .port_i (mixColumns_port_state_out_6_3_7[2:0]), //i
    .port_o (majority_5622_port_o                )  //o
  );
  Majority majority_5623 (
    .port_i (mixColumns_port_state_out_7_3_7[2:0]), //i
    .port_o (majority_5623_port_o                )  //o
  );
  Majority majority_5624 (
    .port_i (mixColumns_port_state_out_8_3_7[2:0]), //i
    .port_o (majority_5624_port_o                )  //o
  );
  Majority majority_5625 (
    .port_i (mixColumns_port_state_out_9_3_7[2:0]), //i
    .port_o (majority_5625_port_o                )  //o
  );
  Majority majority_5626 (
    .port_i (mixColumns_port_state_out_10_3_7[2:0]), //i
    .port_o (majority_5626_port_o                 )  //o
  );
  Majority majority_5627 (
    .port_i (mixColumns_port_state_out_11_3_7[2:0]), //i
    .port_o (majority_5627_port_o                 )  //o
  );
  Majority majority_5628 (
    .port_i (mixColumns_port_state_out_12_3_7[2:0]), //i
    .port_o (majority_5628_port_o                 )  //o
  );
  Majority majority_5629 (
    .port_i (mixColumns_port_state_out_13_3_7[2:0]), //i
    .port_o (majority_5629_port_o                 )  //o
  );
  Majority majority_5630 (
    .port_i (mixColumns_port_state_out_14_3_7[2:0]), //i
    .port_o (majority_5630_port_o                 )  //o
  );
  Majority majority_5631 (
    .port_i (mixColumns_port_state_out_15_3_7[2:0]), //i
    .port_o (majority_5631_port_o                 )  //o
  );
  Majority majority_5632 (
    .port_i (mixColumns_port_state_out_0_0_0[2:0]), //i
    .port_o (majority_5632_port_o                )  //o
  );
  Majority majority_5633 (
    .port_i (mixColumns_port_state_out_1_0_0[2:0]), //i
    .port_o (majority_5633_port_o                )  //o
  );
  Majority majority_5634 (
    .port_i (mixColumns_port_state_out_2_0_0[2:0]), //i
    .port_o (majority_5634_port_o                )  //o
  );
  Majority majority_5635 (
    .port_i (mixColumns_port_state_out_3_0_0[2:0]), //i
    .port_o (majority_5635_port_o                )  //o
  );
  Majority majority_5636 (
    .port_i (mixColumns_port_state_out_4_0_0[2:0]), //i
    .port_o (majority_5636_port_o                )  //o
  );
  Majority majority_5637 (
    .port_i (mixColumns_port_state_out_5_0_0[2:0]), //i
    .port_o (majority_5637_port_o                )  //o
  );
  Majority majority_5638 (
    .port_i (mixColumns_port_state_out_6_0_0[2:0]), //i
    .port_o (majority_5638_port_o                )  //o
  );
  Majority majority_5639 (
    .port_i (mixColumns_port_state_out_7_0_0[2:0]), //i
    .port_o (majority_5639_port_o                )  //o
  );
  Majority majority_5640 (
    .port_i (mixColumns_port_state_out_8_0_0[2:0]), //i
    .port_o (majority_5640_port_o                )  //o
  );
  Majority majority_5641 (
    .port_i (mixColumns_port_state_out_9_0_0[2:0]), //i
    .port_o (majority_5641_port_o                )  //o
  );
  Majority majority_5642 (
    .port_i (mixColumns_port_state_out_10_0_0[2:0]), //i
    .port_o (majority_5642_port_o                 )  //o
  );
  Majority majority_5643 (
    .port_i (mixColumns_port_state_out_11_0_0[2:0]), //i
    .port_o (majority_5643_port_o                 )  //o
  );
  Majority majority_5644 (
    .port_i (mixColumns_port_state_out_12_0_0[2:0]), //i
    .port_o (majority_5644_port_o                 )  //o
  );
  Majority majority_5645 (
    .port_i (mixColumns_port_state_out_13_0_0[2:0]), //i
    .port_o (majority_5645_port_o                 )  //o
  );
  Majority majority_5646 (
    .port_i (mixColumns_port_state_out_14_0_0[2:0]), //i
    .port_o (majority_5646_port_o                 )  //o
  );
  Majority majority_5647 (
    .port_i (mixColumns_port_state_out_15_0_0[2:0]), //i
    .port_o (majority_5647_port_o                 )  //o
  );
  Majority majority_5648 (
    .port_i (mixColumns_port_state_out_0_1_0[2:0]), //i
    .port_o (majority_5648_port_o                )  //o
  );
  Majority majority_5649 (
    .port_i (mixColumns_port_state_out_1_1_0[2:0]), //i
    .port_o (majority_5649_port_o                )  //o
  );
  Majority majority_5650 (
    .port_i (mixColumns_port_state_out_2_1_0[2:0]), //i
    .port_o (majority_5650_port_o                )  //o
  );
  Majority majority_5651 (
    .port_i (mixColumns_port_state_out_3_1_0[2:0]), //i
    .port_o (majority_5651_port_o                )  //o
  );
  Majority majority_5652 (
    .port_i (mixColumns_port_state_out_4_1_0[2:0]), //i
    .port_o (majority_5652_port_o                )  //o
  );
  Majority majority_5653 (
    .port_i (mixColumns_port_state_out_5_1_0[2:0]), //i
    .port_o (majority_5653_port_o                )  //o
  );
  Majority majority_5654 (
    .port_i (mixColumns_port_state_out_6_1_0[2:0]), //i
    .port_o (majority_5654_port_o                )  //o
  );
  Majority majority_5655 (
    .port_i (mixColumns_port_state_out_7_1_0[2:0]), //i
    .port_o (majority_5655_port_o                )  //o
  );
  Majority majority_5656 (
    .port_i (mixColumns_port_state_out_8_1_0[2:0]), //i
    .port_o (majority_5656_port_o                )  //o
  );
  Majority majority_5657 (
    .port_i (mixColumns_port_state_out_9_1_0[2:0]), //i
    .port_o (majority_5657_port_o                )  //o
  );
  Majority majority_5658 (
    .port_i (mixColumns_port_state_out_10_1_0[2:0]), //i
    .port_o (majority_5658_port_o                 )  //o
  );
  Majority majority_5659 (
    .port_i (mixColumns_port_state_out_11_1_0[2:0]), //i
    .port_o (majority_5659_port_o                 )  //o
  );
  Majority majority_5660 (
    .port_i (mixColumns_port_state_out_12_1_0[2:0]), //i
    .port_o (majority_5660_port_o                 )  //o
  );
  Majority majority_5661 (
    .port_i (mixColumns_port_state_out_13_1_0[2:0]), //i
    .port_o (majority_5661_port_o                 )  //o
  );
  Majority majority_5662 (
    .port_i (mixColumns_port_state_out_14_1_0[2:0]), //i
    .port_o (majority_5662_port_o                 )  //o
  );
  Majority majority_5663 (
    .port_i (mixColumns_port_state_out_15_1_0[2:0]), //i
    .port_o (majority_5663_port_o                 )  //o
  );
  Majority majority_5664 (
    .port_i (mixColumns_port_state_out_0_2_0[2:0]), //i
    .port_o (majority_5664_port_o                )  //o
  );
  Majority majority_5665 (
    .port_i (mixColumns_port_state_out_1_2_0[2:0]), //i
    .port_o (majority_5665_port_o                )  //o
  );
  Majority majority_5666 (
    .port_i (mixColumns_port_state_out_2_2_0[2:0]), //i
    .port_o (majority_5666_port_o                )  //o
  );
  Majority majority_5667 (
    .port_i (mixColumns_port_state_out_3_2_0[2:0]), //i
    .port_o (majority_5667_port_o                )  //o
  );
  Majority majority_5668 (
    .port_i (mixColumns_port_state_out_4_2_0[2:0]), //i
    .port_o (majority_5668_port_o                )  //o
  );
  Majority majority_5669 (
    .port_i (mixColumns_port_state_out_5_2_0[2:0]), //i
    .port_o (majority_5669_port_o                )  //o
  );
  Majority majority_5670 (
    .port_i (mixColumns_port_state_out_6_2_0[2:0]), //i
    .port_o (majority_5670_port_o                )  //o
  );
  Majority majority_5671 (
    .port_i (mixColumns_port_state_out_7_2_0[2:0]), //i
    .port_o (majority_5671_port_o                )  //o
  );
  Majority majority_5672 (
    .port_i (mixColumns_port_state_out_8_2_0[2:0]), //i
    .port_o (majority_5672_port_o                )  //o
  );
  Majority majority_5673 (
    .port_i (mixColumns_port_state_out_9_2_0[2:0]), //i
    .port_o (majority_5673_port_o                )  //o
  );
  Majority majority_5674 (
    .port_i (mixColumns_port_state_out_10_2_0[2:0]), //i
    .port_o (majority_5674_port_o                 )  //o
  );
  Majority majority_5675 (
    .port_i (mixColumns_port_state_out_11_2_0[2:0]), //i
    .port_o (majority_5675_port_o                 )  //o
  );
  Majority majority_5676 (
    .port_i (mixColumns_port_state_out_12_2_0[2:0]), //i
    .port_o (majority_5676_port_o                 )  //o
  );
  Majority majority_5677 (
    .port_i (mixColumns_port_state_out_13_2_0[2:0]), //i
    .port_o (majority_5677_port_o                 )  //o
  );
  Majority majority_5678 (
    .port_i (mixColumns_port_state_out_14_2_0[2:0]), //i
    .port_o (majority_5678_port_o                 )  //o
  );
  Majority majority_5679 (
    .port_i (mixColumns_port_state_out_15_2_0[2:0]), //i
    .port_o (majority_5679_port_o                 )  //o
  );
  Majority majority_5680 (
    .port_i (mixColumns_port_state_out_0_3_0[2:0]), //i
    .port_o (majority_5680_port_o                )  //o
  );
  Majority majority_5681 (
    .port_i (mixColumns_port_state_out_1_3_0[2:0]), //i
    .port_o (majority_5681_port_o                )  //o
  );
  Majority majority_5682 (
    .port_i (mixColumns_port_state_out_2_3_0[2:0]), //i
    .port_o (majority_5682_port_o                )  //o
  );
  Majority majority_5683 (
    .port_i (mixColumns_port_state_out_3_3_0[2:0]), //i
    .port_o (majority_5683_port_o                )  //o
  );
  Majority majority_5684 (
    .port_i (mixColumns_port_state_out_4_3_0[2:0]), //i
    .port_o (majority_5684_port_o                )  //o
  );
  Majority majority_5685 (
    .port_i (mixColumns_port_state_out_5_3_0[2:0]), //i
    .port_o (majority_5685_port_o                )  //o
  );
  Majority majority_5686 (
    .port_i (mixColumns_port_state_out_6_3_0[2:0]), //i
    .port_o (majority_5686_port_o                )  //o
  );
  Majority majority_5687 (
    .port_i (mixColumns_port_state_out_7_3_0[2:0]), //i
    .port_o (majority_5687_port_o                )  //o
  );
  Majority majority_5688 (
    .port_i (mixColumns_port_state_out_8_3_0[2:0]), //i
    .port_o (majority_5688_port_o                )  //o
  );
  Majority majority_5689 (
    .port_i (mixColumns_port_state_out_9_3_0[2:0]), //i
    .port_o (majority_5689_port_o                )  //o
  );
  Majority majority_5690 (
    .port_i (mixColumns_port_state_out_10_3_0[2:0]), //i
    .port_o (majority_5690_port_o                 )  //o
  );
  Majority majority_5691 (
    .port_i (mixColumns_port_state_out_11_3_0[2:0]), //i
    .port_o (majority_5691_port_o                 )  //o
  );
  Majority majority_5692 (
    .port_i (mixColumns_port_state_out_12_3_0[2:0]), //i
    .port_o (majority_5692_port_o                 )  //o
  );
  Majority majority_5693 (
    .port_i (mixColumns_port_state_out_13_3_0[2:0]), //i
    .port_o (majority_5693_port_o                 )  //o
  );
  Majority majority_5694 (
    .port_i (mixColumns_port_state_out_14_3_0[2:0]), //i
    .port_o (majority_5694_port_o                 )  //o
  );
  Majority majority_5695 (
    .port_i (mixColumns_port_state_out_15_3_0[2:0]), //i
    .port_o (majority_5695_port_o                 )  //o
  );
  Majority majority_5696 (
    .port_i (mixColumns_port_state_out_0_0_1[2:0]), //i
    .port_o (majority_5696_port_o                )  //o
  );
  Majority majority_5697 (
    .port_i (mixColumns_port_state_out_1_0_1[2:0]), //i
    .port_o (majority_5697_port_o                )  //o
  );
  Majority majority_5698 (
    .port_i (mixColumns_port_state_out_2_0_1[2:0]), //i
    .port_o (majority_5698_port_o                )  //o
  );
  Majority majority_5699 (
    .port_i (mixColumns_port_state_out_3_0_1[2:0]), //i
    .port_o (majority_5699_port_o                )  //o
  );
  Majority majority_5700 (
    .port_i (mixColumns_port_state_out_4_0_1[2:0]), //i
    .port_o (majority_5700_port_o                )  //o
  );
  Majority majority_5701 (
    .port_i (mixColumns_port_state_out_5_0_1[2:0]), //i
    .port_o (majority_5701_port_o                )  //o
  );
  Majority majority_5702 (
    .port_i (mixColumns_port_state_out_6_0_1[2:0]), //i
    .port_o (majority_5702_port_o                )  //o
  );
  Majority majority_5703 (
    .port_i (mixColumns_port_state_out_7_0_1[2:0]), //i
    .port_o (majority_5703_port_o                )  //o
  );
  Majority majority_5704 (
    .port_i (mixColumns_port_state_out_8_0_1[2:0]), //i
    .port_o (majority_5704_port_o                )  //o
  );
  Majority majority_5705 (
    .port_i (mixColumns_port_state_out_9_0_1[2:0]), //i
    .port_o (majority_5705_port_o                )  //o
  );
  Majority majority_5706 (
    .port_i (mixColumns_port_state_out_10_0_1[2:0]), //i
    .port_o (majority_5706_port_o                 )  //o
  );
  Majority majority_5707 (
    .port_i (mixColumns_port_state_out_11_0_1[2:0]), //i
    .port_o (majority_5707_port_o                 )  //o
  );
  Majority majority_5708 (
    .port_i (mixColumns_port_state_out_12_0_1[2:0]), //i
    .port_o (majority_5708_port_o                 )  //o
  );
  Majority majority_5709 (
    .port_i (mixColumns_port_state_out_13_0_1[2:0]), //i
    .port_o (majority_5709_port_o                 )  //o
  );
  Majority majority_5710 (
    .port_i (mixColumns_port_state_out_14_0_1[2:0]), //i
    .port_o (majority_5710_port_o                 )  //o
  );
  Majority majority_5711 (
    .port_i (mixColumns_port_state_out_15_0_1[2:0]), //i
    .port_o (majority_5711_port_o                 )  //o
  );
  Majority majority_5712 (
    .port_i (mixColumns_port_state_out_0_1_1[2:0]), //i
    .port_o (majority_5712_port_o                )  //o
  );
  Majority majority_5713 (
    .port_i (mixColumns_port_state_out_1_1_1[2:0]), //i
    .port_o (majority_5713_port_o                )  //o
  );
  Majority majority_5714 (
    .port_i (mixColumns_port_state_out_2_1_1[2:0]), //i
    .port_o (majority_5714_port_o                )  //o
  );
  Majority majority_5715 (
    .port_i (mixColumns_port_state_out_3_1_1[2:0]), //i
    .port_o (majority_5715_port_o                )  //o
  );
  Majority majority_5716 (
    .port_i (mixColumns_port_state_out_4_1_1[2:0]), //i
    .port_o (majority_5716_port_o                )  //o
  );
  Majority majority_5717 (
    .port_i (mixColumns_port_state_out_5_1_1[2:0]), //i
    .port_o (majority_5717_port_o                )  //o
  );
  Majority majority_5718 (
    .port_i (mixColumns_port_state_out_6_1_1[2:0]), //i
    .port_o (majority_5718_port_o                )  //o
  );
  Majority majority_5719 (
    .port_i (mixColumns_port_state_out_7_1_1[2:0]), //i
    .port_o (majority_5719_port_o                )  //o
  );
  Majority majority_5720 (
    .port_i (mixColumns_port_state_out_8_1_1[2:0]), //i
    .port_o (majority_5720_port_o                )  //o
  );
  Majority majority_5721 (
    .port_i (mixColumns_port_state_out_9_1_1[2:0]), //i
    .port_o (majority_5721_port_o                )  //o
  );
  Majority majority_5722 (
    .port_i (mixColumns_port_state_out_10_1_1[2:0]), //i
    .port_o (majority_5722_port_o                 )  //o
  );
  Majority majority_5723 (
    .port_i (mixColumns_port_state_out_11_1_1[2:0]), //i
    .port_o (majority_5723_port_o                 )  //o
  );
  Majority majority_5724 (
    .port_i (mixColumns_port_state_out_12_1_1[2:0]), //i
    .port_o (majority_5724_port_o                 )  //o
  );
  Majority majority_5725 (
    .port_i (mixColumns_port_state_out_13_1_1[2:0]), //i
    .port_o (majority_5725_port_o                 )  //o
  );
  Majority majority_5726 (
    .port_i (mixColumns_port_state_out_14_1_1[2:0]), //i
    .port_o (majority_5726_port_o                 )  //o
  );
  Majority majority_5727 (
    .port_i (mixColumns_port_state_out_15_1_1[2:0]), //i
    .port_o (majority_5727_port_o                 )  //o
  );
  Majority majority_5728 (
    .port_i (mixColumns_port_state_out_0_2_1[2:0]), //i
    .port_o (majority_5728_port_o                )  //o
  );
  Majority majority_5729 (
    .port_i (mixColumns_port_state_out_1_2_1[2:0]), //i
    .port_o (majority_5729_port_o                )  //o
  );
  Majority majority_5730 (
    .port_i (mixColumns_port_state_out_2_2_1[2:0]), //i
    .port_o (majority_5730_port_o                )  //o
  );
  Majority majority_5731 (
    .port_i (mixColumns_port_state_out_3_2_1[2:0]), //i
    .port_o (majority_5731_port_o                )  //o
  );
  Majority majority_5732 (
    .port_i (mixColumns_port_state_out_4_2_1[2:0]), //i
    .port_o (majority_5732_port_o                )  //o
  );
  Majority majority_5733 (
    .port_i (mixColumns_port_state_out_5_2_1[2:0]), //i
    .port_o (majority_5733_port_o                )  //o
  );
  Majority majority_5734 (
    .port_i (mixColumns_port_state_out_6_2_1[2:0]), //i
    .port_o (majority_5734_port_o                )  //o
  );
  Majority majority_5735 (
    .port_i (mixColumns_port_state_out_7_2_1[2:0]), //i
    .port_o (majority_5735_port_o                )  //o
  );
  Majority majority_5736 (
    .port_i (mixColumns_port_state_out_8_2_1[2:0]), //i
    .port_o (majority_5736_port_o                )  //o
  );
  Majority majority_5737 (
    .port_i (mixColumns_port_state_out_9_2_1[2:0]), //i
    .port_o (majority_5737_port_o                )  //o
  );
  Majority majority_5738 (
    .port_i (mixColumns_port_state_out_10_2_1[2:0]), //i
    .port_o (majority_5738_port_o                 )  //o
  );
  Majority majority_5739 (
    .port_i (mixColumns_port_state_out_11_2_1[2:0]), //i
    .port_o (majority_5739_port_o                 )  //o
  );
  Majority majority_5740 (
    .port_i (mixColumns_port_state_out_12_2_1[2:0]), //i
    .port_o (majority_5740_port_o                 )  //o
  );
  Majority majority_5741 (
    .port_i (mixColumns_port_state_out_13_2_1[2:0]), //i
    .port_o (majority_5741_port_o                 )  //o
  );
  Majority majority_5742 (
    .port_i (mixColumns_port_state_out_14_2_1[2:0]), //i
    .port_o (majority_5742_port_o                 )  //o
  );
  Majority majority_5743 (
    .port_i (mixColumns_port_state_out_15_2_1[2:0]), //i
    .port_o (majority_5743_port_o                 )  //o
  );
  Majority majority_5744 (
    .port_i (mixColumns_port_state_out_0_3_1[2:0]), //i
    .port_o (majority_5744_port_o                )  //o
  );
  Majority majority_5745 (
    .port_i (mixColumns_port_state_out_1_3_1[2:0]), //i
    .port_o (majority_5745_port_o                )  //o
  );
  Majority majority_5746 (
    .port_i (mixColumns_port_state_out_2_3_1[2:0]), //i
    .port_o (majority_5746_port_o                )  //o
  );
  Majority majority_5747 (
    .port_i (mixColumns_port_state_out_3_3_1[2:0]), //i
    .port_o (majority_5747_port_o                )  //o
  );
  Majority majority_5748 (
    .port_i (mixColumns_port_state_out_4_3_1[2:0]), //i
    .port_o (majority_5748_port_o                )  //o
  );
  Majority majority_5749 (
    .port_i (mixColumns_port_state_out_5_3_1[2:0]), //i
    .port_o (majority_5749_port_o                )  //o
  );
  Majority majority_5750 (
    .port_i (mixColumns_port_state_out_6_3_1[2:0]), //i
    .port_o (majority_5750_port_o                )  //o
  );
  Majority majority_5751 (
    .port_i (mixColumns_port_state_out_7_3_1[2:0]), //i
    .port_o (majority_5751_port_o                )  //o
  );
  Majority majority_5752 (
    .port_i (mixColumns_port_state_out_8_3_1[2:0]), //i
    .port_o (majority_5752_port_o                )  //o
  );
  Majority majority_5753 (
    .port_i (mixColumns_port_state_out_9_3_1[2:0]), //i
    .port_o (majority_5753_port_o                )  //o
  );
  Majority majority_5754 (
    .port_i (mixColumns_port_state_out_10_3_1[2:0]), //i
    .port_o (majority_5754_port_o                 )  //o
  );
  Majority majority_5755 (
    .port_i (mixColumns_port_state_out_11_3_1[2:0]), //i
    .port_o (majority_5755_port_o                 )  //o
  );
  Majority majority_5756 (
    .port_i (mixColumns_port_state_out_12_3_1[2:0]), //i
    .port_o (majority_5756_port_o                 )  //o
  );
  Majority majority_5757 (
    .port_i (mixColumns_port_state_out_13_3_1[2:0]), //i
    .port_o (majority_5757_port_o                 )  //o
  );
  Majority majority_5758 (
    .port_i (mixColumns_port_state_out_14_3_1[2:0]), //i
    .port_o (majority_5758_port_o                 )  //o
  );
  Majority majority_5759 (
    .port_i (mixColumns_port_state_out_15_3_1[2:0]), //i
    .port_o (majority_5759_port_o                 )  //o
  );
  Majority majority_5760 (
    .port_i (mixColumns_port_state_out_0_0_2[2:0]), //i
    .port_o (majority_5760_port_o                )  //o
  );
  Majority majority_5761 (
    .port_i (mixColumns_port_state_out_1_0_2[2:0]), //i
    .port_o (majority_5761_port_o                )  //o
  );
  Majority majority_5762 (
    .port_i (mixColumns_port_state_out_2_0_2[2:0]), //i
    .port_o (majority_5762_port_o                )  //o
  );
  Majority majority_5763 (
    .port_i (mixColumns_port_state_out_3_0_2[2:0]), //i
    .port_o (majority_5763_port_o                )  //o
  );
  Majority majority_5764 (
    .port_i (mixColumns_port_state_out_4_0_2[2:0]), //i
    .port_o (majority_5764_port_o                )  //o
  );
  Majority majority_5765 (
    .port_i (mixColumns_port_state_out_5_0_2[2:0]), //i
    .port_o (majority_5765_port_o                )  //o
  );
  Majority majority_5766 (
    .port_i (mixColumns_port_state_out_6_0_2[2:0]), //i
    .port_o (majority_5766_port_o                )  //o
  );
  Majority majority_5767 (
    .port_i (mixColumns_port_state_out_7_0_2[2:0]), //i
    .port_o (majority_5767_port_o                )  //o
  );
  Majority majority_5768 (
    .port_i (mixColumns_port_state_out_8_0_2[2:0]), //i
    .port_o (majority_5768_port_o                )  //o
  );
  Majority majority_5769 (
    .port_i (mixColumns_port_state_out_9_0_2[2:0]), //i
    .port_o (majority_5769_port_o                )  //o
  );
  Majority majority_5770 (
    .port_i (mixColumns_port_state_out_10_0_2[2:0]), //i
    .port_o (majority_5770_port_o                 )  //o
  );
  Majority majority_5771 (
    .port_i (mixColumns_port_state_out_11_0_2[2:0]), //i
    .port_o (majority_5771_port_o                 )  //o
  );
  Majority majority_5772 (
    .port_i (mixColumns_port_state_out_12_0_2[2:0]), //i
    .port_o (majority_5772_port_o                 )  //o
  );
  Majority majority_5773 (
    .port_i (mixColumns_port_state_out_13_0_2[2:0]), //i
    .port_o (majority_5773_port_o                 )  //o
  );
  Majority majority_5774 (
    .port_i (mixColumns_port_state_out_14_0_2[2:0]), //i
    .port_o (majority_5774_port_o                 )  //o
  );
  Majority majority_5775 (
    .port_i (mixColumns_port_state_out_15_0_2[2:0]), //i
    .port_o (majority_5775_port_o                 )  //o
  );
  Majority majority_5776 (
    .port_i (mixColumns_port_state_out_0_1_2[2:0]), //i
    .port_o (majority_5776_port_o                )  //o
  );
  Majority majority_5777 (
    .port_i (mixColumns_port_state_out_1_1_2[2:0]), //i
    .port_o (majority_5777_port_o                )  //o
  );
  Majority majority_5778 (
    .port_i (mixColumns_port_state_out_2_1_2[2:0]), //i
    .port_o (majority_5778_port_o                )  //o
  );
  Majority majority_5779 (
    .port_i (mixColumns_port_state_out_3_1_2[2:0]), //i
    .port_o (majority_5779_port_o                )  //o
  );
  Majority majority_5780 (
    .port_i (mixColumns_port_state_out_4_1_2[2:0]), //i
    .port_o (majority_5780_port_o                )  //o
  );
  Majority majority_5781 (
    .port_i (mixColumns_port_state_out_5_1_2[2:0]), //i
    .port_o (majority_5781_port_o                )  //o
  );
  Majority majority_5782 (
    .port_i (mixColumns_port_state_out_6_1_2[2:0]), //i
    .port_o (majority_5782_port_o                )  //o
  );
  Majority majority_5783 (
    .port_i (mixColumns_port_state_out_7_1_2[2:0]), //i
    .port_o (majority_5783_port_o                )  //o
  );
  Majority majority_5784 (
    .port_i (mixColumns_port_state_out_8_1_2[2:0]), //i
    .port_o (majority_5784_port_o                )  //o
  );
  Majority majority_5785 (
    .port_i (mixColumns_port_state_out_9_1_2[2:0]), //i
    .port_o (majority_5785_port_o                )  //o
  );
  Majority majority_5786 (
    .port_i (mixColumns_port_state_out_10_1_2[2:0]), //i
    .port_o (majority_5786_port_o                 )  //o
  );
  Majority majority_5787 (
    .port_i (mixColumns_port_state_out_11_1_2[2:0]), //i
    .port_o (majority_5787_port_o                 )  //o
  );
  Majority majority_5788 (
    .port_i (mixColumns_port_state_out_12_1_2[2:0]), //i
    .port_o (majority_5788_port_o                 )  //o
  );
  Majority majority_5789 (
    .port_i (mixColumns_port_state_out_13_1_2[2:0]), //i
    .port_o (majority_5789_port_o                 )  //o
  );
  Majority majority_5790 (
    .port_i (mixColumns_port_state_out_14_1_2[2:0]), //i
    .port_o (majority_5790_port_o                 )  //o
  );
  Majority majority_5791 (
    .port_i (mixColumns_port_state_out_15_1_2[2:0]), //i
    .port_o (majority_5791_port_o                 )  //o
  );
  Majority majority_5792 (
    .port_i (mixColumns_port_state_out_0_2_2[2:0]), //i
    .port_o (majority_5792_port_o                )  //o
  );
  Majority majority_5793 (
    .port_i (mixColumns_port_state_out_1_2_2[2:0]), //i
    .port_o (majority_5793_port_o                )  //o
  );
  Majority majority_5794 (
    .port_i (mixColumns_port_state_out_2_2_2[2:0]), //i
    .port_o (majority_5794_port_o                )  //o
  );
  Majority majority_5795 (
    .port_i (mixColumns_port_state_out_3_2_2[2:0]), //i
    .port_o (majority_5795_port_o                )  //o
  );
  Majority majority_5796 (
    .port_i (mixColumns_port_state_out_4_2_2[2:0]), //i
    .port_o (majority_5796_port_o                )  //o
  );
  Majority majority_5797 (
    .port_i (mixColumns_port_state_out_5_2_2[2:0]), //i
    .port_o (majority_5797_port_o                )  //o
  );
  Majority majority_5798 (
    .port_i (mixColumns_port_state_out_6_2_2[2:0]), //i
    .port_o (majority_5798_port_o                )  //o
  );
  Majority majority_5799 (
    .port_i (mixColumns_port_state_out_7_2_2[2:0]), //i
    .port_o (majority_5799_port_o                )  //o
  );
  Majority majority_5800 (
    .port_i (mixColumns_port_state_out_8_2_2[2:0]), //i
    .port_o (majority_5800_port_o                )  //o
  );
  Majority majority_5801 (
    .port_i (mixColumns_port_state_out_9_2_2[2:0]), //i
    .port_o (majority_5801_port_o                )  //o
  );
  Majority majority_5802 (
    .port_i (mixColumns_port_state_out_10_2_2[2:0]), //i
    .port_o (majority_5802_port_o                 )  //o
  );
  Majority majority_5803 (
    .port_i (mixColumns_port_state_out_11_2_2[2:0]), //i
    .port_o (majority_5803_port_o                 )  //o
  );
  Majority majority_5804 (
    .port_i (mixColumns_port_state_out_12_2_2[2:0]), //i
    .port_o (majority_5804_port_o                 )  //o
  );
  Majority majority_5805 (
    .port_i (mixColumns_port_state_out_13_2_2[2:0]), //i
    .port_o (majority_5805_port_o                 )  //o
  );
  Majority majority_5806 (
    .port_i (mixColumns_port_state_out_14_2_2[2:0]), //i
    .port_o (majority_5806_port_o                 )  //o
  );
  Majority majority_5807 (
    .port_i (mixColumns_port_state_out_15_2_2[2:0]), //i
    .port_o (majority_5807_port_o                 )  //o
  );
  Majority majority_5808 (
    .port_i (mixColumns_port_state_out_0_3_2[2:0]), //i
    .port_o (majority_5808_port_o                )  //o
  );
  Majority majority_5809 (
    .port_i (mixColumns_port_state_out_1_3_2[2:0]), //i
    .port_o (majority_5809_port_o                )  //o
  );
  Majority majority_5810 (
    .port_i (mixColumns_port_state_out_2_3_2[2:0]), //i
    .port_o (majority_5810_port_o                )  //o
  );
  Majority majority_5811 (
    .port_i (mixColumns_port_state_out_3_3_2[2:0]), //i
    .port_o (majority_5811_port_o                )  //o
  );
  Majority majority_5812 (
    .port_i (mixColumns_port_state_out_4_3_2[2:0]), //i
    .port_o (majority_5812_port_o                )  //o
  );
  Majority majority_5813 (
    .port_i (mixColumns_port_state_out_5_3_2[2:0]), //i
    .port_o (majority_5813_port_o                )  //o
  );
  Majority majority_5814 (
    .port_i (mixColumns_port_state_out_6_3_2[2:0]), //i
    .port_o (majority_5814_port_o                )  //o
  );
  Majority majority_5815 (
    .port_i (mixColumns_port_state_out_7_3_2[2:0]), //i
    .port_o (majority_5815_port_o                )  //o
  );
  Majority majority_5816 (
    .port_i (mixColumns_port_state_out_8_3_2[2:0]), //i
    .port_o (majority_5816_port_o                )  //o
  );
  Majority majority_5817 (
    .port_i (mixColumns_port_state_out_9_3_2[2:0]), //i
    .port_o (majority_5817_port_o                )  //o
  );
  Majority majority_5818 (
    .port_i (mixColumns_port_state_out_10_3_2[2:0]), //i
    .port_o (majority_5818_port_o                 )  //o
  );
  Majority majority_5819 (
    .port_i (mixColumns_port_state_out_11_3_2[2:0]), //i
    .port_o (majority_5819_port_o                 )  //o
  );
  Majority majority_5820 (
    .port_i (mixColumns_port_state_out_12_3_2[2:0]), //i
    .port_o (majority_5820_port_o                 )  //o
  );
  Majority majority_5821 (
    .port_i (mixColumns_port_state_out_13_3_2[2:0]), //i
    .port_o (majority_5821_port_o                 )  //o
  );
  Majority majority_5822 (
    .port_i (mixColumns_port_state_out_14_3_2[2:0]), //i
    .port_o (majority_5822_port_o                 )  //o
  );
  Majority majority_5823 (
    .port_i (mixColumns_port_state_out_15_3_2[2:0]), //i
    .port_o (majority_5823_port_o                 )  //o
  );
  Majority majority_5824 (
    .port_i (mixColumns_port_state_out_0_0_3[2:0]), //i
    .port_o (majority_5824_port_o                )  //o
  );
  Majority majority_5825 (
    .port_i (mixColumns_port_state_out_1_0_3[2:0]), //i
    .port_o (majority_5825_port_o                )  //o
  );
  Majority majority_5826 (
    .port_i (mixColumns_port_state_out_2_0_3[2:0]), //i
    .port_o (majority_5826_port_o                )  //o
  );
  Majority majority_5827 (
    .port_i (mixColumns_port_state_out_3_0_3[2:0]), //i
    .port_o (majority_5827_port_o                )  //o
  );
  Majority majority_5828 (
    .port_i (mixColumns_port_state_out_4_0_3[2:0]), //i
    .port_o (majority_5828_port_o                )  //o
  );
  Majority majority_5829 (
    .port_i (mixColumns_port_state_out_5_0_3[2:0]), //i
    .port_o (majority_5829_port_o                )  //o
  );
  Majority majority_5830 (
    .port_i (mixColumns_port_state_out_6_0_3[2:0]), //i
    .port_o (majority_5830_port_o                )  //o
  );
  Majority majority_5831 (
    .port_i (mixColumns_port_state_out_7_0_3[2:0]), //i
    .port_o (majority_5831_port_o                )  //o
  );
  Majority majority_5832 (
    .port_i (mixColumns_port_state_out_8_0_3[2:0]), //i
    .port_o (majority_5832_port_o                )  //o
  );
  Majority majority_5833 (
    .port_i (mixColumns_port_state_out_9_0_3[2:0]), //i
    .port_o (majority_5833_port_o                )  //o
  );
  Majority majority_5834 (
    .port_i (mixColumns_port_state_out_10_0_3[2:0]), //i
    .port_o (majority_5834_port_o                 )  //o
  );
  Majority majority_5835 (
    .port_i (mixColumns_port_state_out_11_0_3[2:0]), //i
    .port_o (majority_5835_port_o                 )  //o
  );
  Majority majority_5836 (
    .port_i (mixColumns_port_state_out_12_0_3[2:0]), //i
    .port_o (majority_5836_port_o                 )  //o
  );
  Majority majority_5837 (
    .port_i (mixColumns_port_state_out_13_0_3[2:0]), //i
    .port_o (majority_5837_port_o                 )  //o
  );
  Majority majority_5838 (
    .port_i (mixColumns_port_state_out_14_0_3[2:0]), //i
    .port_o (majority_5838_port_o                 )  //o
  );
  Majority majority_5839 (
    .port_i (mixColumns_port_state_out_15_0_3[2:0]), //i
    .port_o (majority_5839_port_o                 )  //o
  );
  Majority majority_5840 (
    .port_i (mixColumns_port_state_out_0_1_3[2:0]), //i
    .port_o (majority_5840_port_o                )  //o
  );
  Majority majority_5841 (
    .port_i (mixColumns_port_state_out_1_1_3[2:0]), //i
    .port_o (majority_5841_port_o                )  //o
  );
  Majority majority_5842 (
    .port_i (mixColumns_port_state_out_2_1_3[2:0]), //i
    .port_o (majority_5842_port_o                )  //o
  );
  Majority majority_5843 (
    .port_i (mixColumns_port_state_out_3_1_3[2:0]), //i
    .port_o (majority_5843_port_o                )  //o
  );
  Majority majority_5844 (
    .port_i (mixColumns_port_state_out_4_1_3[2:0]), //i
    .port_o (majority_5844_port_o                )  //o
  );
  Majority majority_5845 (
    .port_i (mixColumns_port_state_out_5_1_3[2:0]), //i
    .port_o (majority_5845_port_o                )  //o
  );
  Majority majority_5846 (
    .port_i (mixColumns_port_state_out_6_1_3[2:0]), //i
    .port_o (majority_5846_port_o                )  //o
  );
  Majority majority_5847 (
    .port_i (mixColumns_port_state_out_7_1_3[2:0]), //i
    .port_o (majority_5847_port_o                )  //o
  );
  Majority majority_5848 (
    .port_i (mixColumns_port_state_out_8_1_3[2:0]), //i
    .port_o (majority_5848_port_o                )  //o
  );
  Majority majority_5849 (
    .port_i (mixColumns_port_state_out_9_1_3[2:0]), //i
    .port_o (majority_5849_port_o                )  //o
  );
  Majority majority_5850 (
    .port_i (mixColumns_port_state_out_10_1_3[2:0]), //i
    .port_o (majority_5850_port_o                 )  //o
  );
  Majority majority_5851 (
    .port_i (mixColumns_port_state_out_11_1_3[2:0]), //i
    .port_o (majority_5851_port_o                 )  //o
  );
  Majority majority_5852 (
    .port_i (mixColumns_port_state_out_12_1_3[2:0]), //i
    .port_o (majority_5852_port_o                 )  //o
  );
  Majority majority_5853 (
    .port_i (mixColumns_port_state_out_13_1_3[2:0]), //i
    .port_o (majority_5853_port_o                 )  //o
  );
  Majority majority_5854 (
    .port_i (mixColumns_port_state_out_14_1_3[2:0]), //i
    .port_o (majority_5854_port_o                 )  //o
  );
  Majority majority_5855 (
    .port_i (mixColumns_port_state_out_15_1_3[2:0]), //i
    .port_o (majority_5855_port_o                 )  //o
  );
  Majority majority_5856 (
    .port_i (mixColumns_port_state_out_0_2_3[2:0]), //i
    .port_o (majority_5856_port_o                )  //o
  );
  Majority majority_5857 (
    .port_i (mixColumns_port_state_out_1_2_3[2:0]), //i
    .port_o (majority_5857_port_o                )  //o
  );
  Majority majority_5858 (
    .port_i (mixColumns_port_state_out_2_2_3[2:0]), //i
    .port_o (majority_5858_port_o                )  //o
  );
  Majority majority_5859 (
    .port_i (mixColumns_port_state_out_3_2_3[2:0]), //i
    .port_o (majority_5859_port_o                )  //o
  );
  Majority majority_5860 (
    .port_i (mixColumns_port_state_out_4_2_3[2:0]), //i
    .port_o (majority_5860_port_o                )  //o
  );
  Majority majority_5861 (
    .port_i (mixColumns_port_state_out_5_2_3[2:0]), //i
    .port_o (majority_5861_port_o                )  //o
  );
  Majority majority_5862 (
    .port_i (mixColumns_port_state_out_6_2_3[2:0]), //i
    .port_o (majority_5862_port_o                )  //o
  );
  Majority majority_5863 (
    .port_i (mixColumns_port_state_out_7_2_3[2:0]), //i
    .port_o (majority_5863_port_o                )  //o
  );
  Majority majority_5864 (
    .port_i (mixColumns_port_state_out_8_2_3[2:0]), //i
    .port_o (majority_5864_port_o                )  //o
  );
  Majority majority_5865 (
    .port_i (mixColumns_port_state_out_9_2_3[2:0]), //i
    .port_o (majority_5865_port_o                )  //o
  );
  Majority majority_5866 (
    .port_i (mixColumns_port_state_out_10_2_3[2:0]), //i
    .port_o (majority_5866_port_o                 )  //o
  );
  Majority majority_5867 (
    .port_i (mixColumns_port_state_out_11_2_3[2:0]), //i
    .port_o (majority_5867_port_o                 )  //o
  );
  Majority majority_5868 (
    .port_i (mixColumns_port_state_out_12_2_3[2:0]), //i
    .port_o (majority_5868_port_o                 )  //o
  );
  Majority majority_5869 (
    .port_i (mixColumns_port_state_out_13_2_3[2:0]), //i
    .port_o (majority_5869_port_o                 )  //o
  );
  Majority majority_5870 (
    .port_i (mixColumns_port_state_out_14_2_3[2:0]), //i
    .port_o (majority_5870_port_o                 )  //o
  );
  Majority majority_5871 (
    .port_i (mixColumns_port_state_out_15_2_3[2:0]), //i
    .port_o (majority_5871_port_o                 )  //o
  );
  Majority majority_5872 (
    .port_i (mixColumns_port_state_out_0_3_3[2:0]), //i
    .port_o (majority_5872_port_o                )  //o
  );
  Majority majority_5873 (
    .port_i (mixColumns_port_state_out_1_3_3[2:0]), //i
    .port_o (majority_5873_port_o                )  //o
  );
  Majority majority_5874 (
    .port_i (mixColumns_port_state_out_2_3_3[2:0]), //i
    .port_o (majority_5874_port_o                )  //o
  );
  Majority majority_5875 (
    .port_i (mixColumns_port_state_out_3_3_3[2:0]), //i
    .port_o (majority_5875_port_o                )  //o
  );
  Majority majority_5876 (
    .port_i (mixColumns_port_state_out_4_3_3[2:0]), //i
    .port_o (majority_5876_port_o                )  //o
  );
  Majority majority_5877 (
    .port_i (mixColumns_port_state_out_5_3_3[2:0]), //i
    .port_o (majority_5877_port_o                )  //o
  );
  Majority majority_5878 (
    .port_i (mixColumns_port_state_out_6_3_3[2:0]), //i
    .port_o (majority_5878_port_o                )  //o
  );
  Majority majority_5879 (
    .port_i (mixColumns_port_state_out_7_3_3[2:0]), //i
    .port_o (majority_5879_port_o                )  //o
  );
  Majority majority_5880 (
    .port_i (mixColumns_port_state_out_8_3_3[2:0]), //i
    .port_o (majority_5880_port_o                )  //o
  );
  Majority majority_5881 (
    .port_i (mixColumns_port_state_out_9_3_3[2:0]), //i
    .port_o (majority_5881_port_o                )  //o
  );
  Majority majority_5882 (
    .port_i (mixColumns_port_state_out_10_3_3[2:0]), //i
    .port_o (majority_5882_port_o                 )  //o
  );
  Majority majority_5883 (
    .port_i (mixColumns_port_state_out_11_3_3[2:0]), //i
    .port_o (majority_5883_port_o                 )  //o
  );
  Majority majority_5884 (
    .port_i (mixColumns_port_state_out_12_3_3[2:0]), //i
    .port_o (majority_5884_port_o                 )  //o
  );
  Majority majority_5885 (
    .port_i (mixColumns_port_state_out_13_3_3[2:0]), //i
    .port_o (majority_5885_port_o                 )  //o
  );
  Majority majority_5886 (
    .port_i (mixColumns_port_state_out_14_3_3[2:0]), //i
    .port_o (majority_5886_port_o                 )  //o
  );
  Majority majority_5887 (
    .port_i (mixColumns_port_state_out_15_3_3[2:0]), //i
    .port_o (majority_5887_port_o                 )  //o
  );
  Majority majority_5888 (
    .port_i (mixColumns_port_state_out_0_0_4[2:0]), //i
    .port_o (majority_5888_port_o                )  //o
  );
  Majority majority_5889 (
    .port_i (mixColumns_port_state_out_1_0_4[2:0]), //i
    .port_o (majority_5889_port_o                )  //o
  );
  Majority majority_5890 (
    .port_i (mixColumns_port_state_out_2_0_4[2:0]), //i
    .port_o (majority_5890_port_o                )  //o
  );
  Majority majority_5891 (
    .port_i (mixColumns_port_state_out_3_0_4[2:0]), //i
    .port_o (majority_5891_port_o                )  //o
  );
  Majority majority_5892 (
    .port_i (mixColumns_port_state_out_4_0_4[2:0]), //i
    .port_o (majority_5892_port_o                )  //o
  );
  Majority majority_5893 (
    .port_i (mixColumns_port_state_out_5_0_4[2:0]), //i
    .port_o (majority_5893_port_o                )  //o
  );
  Majority majority_5894 (
    .port_i (mixColumns_port_state_out_6_0_4[2:0]), //i
    .port_o (majority_5894_port_o                )  //o
  );
  Majority majority_5895 (
    .port_i (mixColumns_port_state_out_7_0_4[2:0]), //i
    .port_o (majority_5895_port_o                )  //o
  );
  Majority majority_5896 (
    .port_i (mixColumns_port_state_out_8_0_4[2:0]), //i
    .port_o (majority_5896_port_o                )  //o
  );
  Majority majority_5897 (
    .port_i (mixColumns_port_state_out_9_0_4[2:0]), //i
    .port_o (majority_5897_port_o                )  //o
  );
  Majority majority_5898 (
    .port_i (mixColumns_port_state_out_10_0_4[2:0]), //i
    .port_o (majority_5898_port_o                 )  //o
  );
  Majority majority_5899 (
    .port_i (mixColumns_port_state_out_11_0_4[2:0]), //i
    .port_o (majority_5899_port_o                 )  //o
  );
  Majority majority_5900 (
    .port_i (mixColumns_port_state_out_12_0_4[2:0]), //i
    .port_o (majority_5900_port_o                 )  //o
  );
  Majority majority_5901 (
    .port_i (mixColumns_port_state_out_13_0_4[2:0]), //i
    .port_o (majority_5901_port_o                 )  //o
  );
  Majority majority_5902 (
    .port_i (mixColumns_port_state_out_14_0_4[2:0]), //i
    .port_o (majority_5902_port_o                 )  //o
  );
  Majority majority_5903 (
    .port_i (mixColumns_port_state_out_15_0_4[2:0]), //i
    .port_o (majority_5903_port_o                 )  //o
  );
  Majority majority_5904 (
    .port_i (mixColumns_port_state_out_0_1_4[2:0]), //i
    .port_o (majority_5904_port_o                )  //o
  );
  Majority majority_5905 (
    .port_i (mixColumns_port_state_out_1_1_4[2:0]), //i
    .port_o (majority_5905_port_o                )  //o
  );
  Majority majority_5906 (
    .port_i (mixColumns_port_state_out_2_1_4[2:0]), //i
    .port_o (majority_5906_port_o                )  //o
  );
  Majority majority_5907 (
    .port_i (mixColumns_port_state_out_3_1_4[2:0]), //i
    .port_o (majority_5907_port_o                )  //o
  );
  Majority majority_5908 (
    .port_i (mixColumns_port_state_out_4_1_4[2:0]), //i
    .port_o (majority_5908_port_o                )  //o
  );
  Majority majority_5909 (
    .port_i (mixColumns_port_state_out_5_1_4[2:0]), //i
    .port_o (majority_5909_port_o                )  //o
  );
  Majority majority_5910 (
    .port_i (mixColumns_port_state_out_6_1_4[2:0]), //i
    .port_o (majority_5910_port_o                )  //o
  );
  Majority majority_5911 (
    .port_i (mixColumns_port_state_out_7_1_4[2:0]), //i
    .port_o (majority_5911_port_o                )  //o
  );
  Majority majority_5912 (
    .port_i (mixColumns_port_state_out_8_1_4[2:0]), //i
    .port_o (majority_5912_port_o                )  //o
  );
  Majority majority_5913 (
    .port_i (mixColumns_port_state_out_9_1_4[2:0]), //i
    .port_o (majority_5913_port_o                )  //o
  );
  Majority majority_5914 (
    .port_i (mixColumns_port_state_out_10_1_4[2:0]), //i
    .port_o (majority_5914_port_o                 )  //o
  );
  Majority majority_5915 (
    .port_i (mixColumns_port_state_out_11_1_4[2:0]), //i
    .port_o (majority_5915_port_o                 )  //o
  );
  Majority majority_5916 (
    .port_i (mixColumns_port_state_out_12_1_4[2:0]), //i
    .port_o (majority_5916_port_o                 )  //o
  );
  Majority majority_5917 (
    .port_i (mixColumns_port_state_out_13_1_4[2:0]), //i
    .port_o (majority_5917_port_o                 )  //o
  );
  Majority majority_5918 (
    .port_i (mixColumns_port_state_out_14_1_4[2:0]), //i
    .port_o (majority_5918_port_o                 )  //o
  );
  Majority majority_5919 (
    .port_i (mixColumns_port_state_out_15_1_4[2:0]), //i
    .port_o (majority_5919_port_o                 )  //o
  );
  Majority majority_5920 (
    .port_i (mixColumns_port_state_out_0_2_4[2:0]), //i
    .port_o (majority_5920_port_o                )  //o
  );
  Majority majority_5921 (
    .port_i (mixColumns_port_state_out_1_2_4[2:0]), //i
    .port_o (majority_5921_port_o                )  //o
  );
  Majority majority_5922 (
    .port_i (mixColumns_port_state_out_2_2_4[2:0]), //i
    .port_o (majority_5922_port_o                )  //o
  );
  Majority majority_5923 (
    .port_i (mixColumns_port_state_out_3_2_4[2:0]), //i
    .port_o (majority_5923_port_o                )  //o
  );
  Majority majority_5924 (
    .port_i (mixColumns_port_state_out_4_2_4[2:0]), //i
    .port_o (majority_5924_port_o                )  //o
  );
  Majority majority_5925 (
    .port_i (mixColumns_port_state_out_5_2_4[2:0]), //i
    .port_o (majority_5925_port_o                )  //o
  );
  Majority majority_5926 (
    .port_i (mixColumns_port_state_out_6_2_4[2:0]), //i
    .port_o (majority_5926_port_o                )  //o
  );
  Majority majority_5927 (
    .port_i (mixColumns_port_state_out_7_2_4[2:0]), //i
    .port_o (majority_5927_port_o                )  //o
  );
  Majority majority_5928 (
    .port_i (mixColumns_port_state_out_8_2_4[2:0]), //i
    .port_o (majority_5928_port_o                )  //o
  );
  Majority majority_5929 (
    .port_i (mixColumns_port_state_out_9_2_4[2:0]), //i
    .port_o (majority_5929_port_o                )  //o
  );
  Majority majority_5930 (
    .port_i (mixColumns_port_state_out_10_2_4[2:0]), //i
    .port_o (majority_5930_port_o                 )  //o
  );
  Majority majority_5931 (
    .port_i (mixColumns_port_state_out_11_2_4[2:0]), //i
    .port_o (majority_5931_port_o                 )  //o
  );
  Majority majority_5932 (
    .port_i (mixColumns_port_state_out_12_2_4[2:0]), //i
    .port_o (majority_5932_port_o                 )  //o
  );
  Majority majority_5933 (
    .port_i (mixColumns_port_state_out_13_2_4[2:0]), //i
    .port_o (majority_5933_port_o                 )  //o
  );
  Majority majority_5934 (
    .port_i (mixColumns_port_state_out_14_2_4[2:0]), //i
    .port_o (majority_5934_port_o                 )  //o
  );
  Majority majority_5935 (
    .port_i (mixColumns_port_state_out_15_2_4[2:0]), //i
    .port_o (majority_5935_port_o                 )  //o
  );
  Majority majority_5936 (
    .port_i (mixColumns_port_state_out_0_3_4[2:0]), //i
    .port_o (majority_5936_port_o                )  //o
  );
  Majority majority_5937 (
    .port_i (mixColumns_port_state_out_1_3_4[2:0]), //i
    .port_o (majority_5937_port_o                )  //o
  );
  Majority majority_5938 (
    .port_i (mixColumns_port_state_out_2_3_4[2:0]), //i
    .port_o (majority_5938_port_o                )  //o
  );
  Majority majority_5939 (
    .port_i (mixColumns_port_state_out_3_3_4[2:0]), //i
    .port_o (majority_5939_port_o                )  //o
  );
  Majority majority_5940 (
    .port_i (mixColumns_port_state_out_4_3_4[2:0]), //i
    .port_o (majority_5940_port_o                )  //o
  );
  Majority majority_5941 (
    .port_i (mixColumns_port_state_out_5_3_4[2:0]), //i
    .port_o (majority_5941_port_o                )  //o
  );
  Majority majority_5942 (
    .port_i (mixColumns_port_state_out_6_3_4[2:0]), //i
    .port_o (majority_5942_port_o                )  //o
  );
  Majority majority_5943 (
    .port_i (mixColumns_port_state_out_7_3_4[2:0]), //i
    .port_o (majority_5943_port_o                )  //o
  );
  Majority majority_5944 (
    .port_i (mixColumns_port_state_out_8_3_4[2:0]), //i
    .port_o (majority_5944_port_o                )  //o
  );
  Majority majority_5945 (
    .port_i (mixColumns_port_state_out_9_3_4[2:0]), //i
    .port_o (majority_5945_port_o                )  //o
  );
  Majority majority_5946 (
    .port_i (mixColumns_port_state_out_10_3_4[2:0]), //i
    .port_o (majority_5946_port_o                 )  //o
  );
  Majority majority_5947 (
    .port_i (mixColumns_port_state_out_11_3_4[2:0]), //i
    .port_o (majority_5947_port_o                 )  //o
  );
  Majority majority_5948 (
    .port_i (mixColumns_port_state_out_12_3_4[2:0]), //i
    .port_o (majority_5948_port_o                 )  //o
  );
  Majority majority_5949 (
    .port_i (mixColumns_port_state_out_13_3_4[2:0]), //i
    .port_o (majority_5949_port_o                 )  //o
  );
  Majority majority_5950 (
    .port_i (mixColumns_port_state_out_14_3_4[2:0]), //i
    .port_o (majority_5950_port_o                 )  //o
  );
  Majority majority_5951 (
    .port_i (mixColumns_port_state_out_15_3_4[2:0]), //i
    .port_o (majority_5951_port_o                 )  //o
  );
  Majority majority_5952 (
    .port_i (mixColumns_port_state_out_0_0_5[2:0]), //i
    .port_o (majority_5952_port_o                )  //o
  );
  Majority majority_5953 (
    .port_i (mixColumns_port_state_out_1_0_5[2:0]), //i
    .port_o (majority_5953_port_o                )  //o
  );
  Majority majority_5954 (
    .port_i (mixColumns_port_state_out_2_0_5[2:0]), //i
    .port_o (majority_5954_port_o                )  //o
  );
  Majority majority_5955 (
    .port_i (mixColumns_port_state_out_3_0_5[2:0]), //i
    .port_o (majority_5955_port_o                )  //o
  );
  Majority majority_5956 (
    .port_i (mixColumns_port_state_out_4_0_5[2:0]), //i
    .port_o (majority_5956_port_o                )  //o
  );
  Majority majority_5957 (
    .port_i (mixColumns_port_state_out_5_0_5[2:0]), //i
    .port_o (majority_5957_port_o                )  //o
  );
  Majority majority_5958 (
    .port_i (mixColumns_port_state_out_6_0_5[2:0]), //i
    .port_o (majority_5958_port_o                )  //o
  );
  Majority majority_5959 (
    .port_i (mixColumns_port_state_out_7_0_5[2:0]), //i
    .port_o (majority_5959_port_o                )  //o
  );
  Majority majority_5960 (
    .port_i (mixColumns_port_state_out_8_0_5[2:0]), //i
    .port_o (majority_5960_port_o                )  //o
  );
  Majority majority_5961 (
    .port_i (mixColumns_port_state_out_9_0_5[2:0]), //i
    .port_o (majority_5961_port_o                )  //o
  );
  Majority majority_5962 (
    .port_i (mixColumns_port_state_out_10_0_5[2:0]), //i
    .port_o (majority_5962_port_o                 )  //o
  );
  Majority majority_5963 (
    .port_i (mixColumns_port_state_out_11_0_5[2:0]), //i
    .port_o (majority_5963_port_o                 )  //o
  );
  Majority majority_5964 (
    .port_i (mixColumns_port_state_out_12_0_5[2:0]), //i
    .port_o (majority_5964_port_o                 )  //o
  );
  Majority majority_5965 (
    .port_i (mixColumns_port_state_out_13_0_5[2:0]), //i
    .port_o (majority_5965_port_o                 )  //o
  );
  Majority majority_5966 (
    .port_i (mixColumns_port_state_out_14_0_5[2:0]), //i
    .port_o (majority_5966_port_o                 )  //o
  );
  Majority majority_5967 (
    .port_i (mixColumns_port_state_out_15_0_5[2:0]), //i
    .port_o (majority_5967_port_o                 )  //o
  );
  Majority majority_5968 (
    .port_i (mixColumns_port_state_out_0_1_5[2:0]), //i
    .port_o (majority_5968_port_o                )  //o
  );
  Majority majority_5969 (
    .port_i (mixColumns_port_state_out_1_1_5[2:0]), //i
    .port_o (majority_5969_port_o                )  //o
  );
  Majority majority_5970 (
    .port_i (mixColumns_port_state_out_2_1_5[2:0]), //i
    .port_o (majority_5970_port_o                )  //o
  );
  Majority majority_5971 (
    .port_i (mixColumns_port_state_out_3_1_5[2:0]), //i
    .port_o (majority_5971_port_o                )  //o
  );
  Majority majority_5972 (
    .port_i (mixColumns_port_state_out_4_1_5[2:0]), //i
    .port_o (majority_5972_port_o                )  //o
  );
  Majority majority_5973 (
    .port_i (mixColumns_port_state_out_5_1_5[2:0]), //i
    .port_o (majority_5973_port_o                )  //o
  );
  Majority majority_5974 (
    .port_i (mixColumns_port_state_out_6_1_5[2:0]), //i
    .port_o (majority_5974_port_o                )  //o
  );
  Majority majority_5975 (
    .port_i (mixColumns_port_state_out_7_1_5[2:0]), //i
    .port_o (majority_5975_port_o                )  //o
  );
  Majority majority_5976 (
    .port_i (mixColumns_port_state_out_8_1_5[2:0]), //i
    .port_o (majority_5976_port_o                )  //o
  );
  Majority majority_5977 (
    .port_i (mixColumns_port_state_out_9_1_5[2:0]), //i
    .port_o (majority_5977_port_o                )  //o
  );
  Majority majority_5978 (
    .port_i (mixColumns_port_state_out_10_1_5[2:0]), //i
    .port_o (majority_5978_port_o                 )  //o
  );
  Majority majority_5979 (
    .port_i (mixColumns_port_state_out_11_1_5[2:0]), //i
    .port_o (majority_5979_port_o                 )  //o
  );
  Majority majority_5980 (
    .port_i (mixColumns_port_state_out_12_1_5[2:0]), //i
    .port_o (majority_5980_port_o                 )  //o
  );
  Majority majority_5981 (
    .port_i (mixColumns_port_state_out_13_1_5[2:0]), //i
    .port_o (majority_5981_port_o                 )  //o
  );
  Majority majority_5982 (
    .port_i (mixColumns_port_state_out_14_1_5[2:0]), //i
    .port_o (majority_5982_port_o                 )  //o
  );
  Majority majority_5983 (
    .port_i (mixColumns_port_state_out_15_1_5[2:0]), //i
    .port_o (majority_5983_port_o                 )  //o
  );
  Majority majority_5984 (
    .port_i (mixColumns_port_state_out_0_2_5[2:0]), //i
    .port_o (majority_5984_port_o                )  //o
  );
  Majority majority_5985 (
    .port_i (mixColumns_port_state_out_1_2_5[2:0]), //i
    .port_o (majority_5985_port_o                )  //o
  );
  Majority majority_5986 (
    .port_i (mixColumns_port_state_out_2_2_5[2:0]), //i
    .port_o (majority_5986_port_o                )  //o
  );
  Majority majority_5987 (
    .port_i (mixColumns_port_state_out_3_2_5[2:0]), //i
    .port_o (majority_5987_port_o                )  //o
  );
  Majority majority_5988 (
    .port_i (mixColumns_port_state_out_4_2_5[2:0]), //i
    .port_o (majority_5988_port_o                )  //o
  );
  Majority majority_5989 (
    .port_i (mixColumns_port_state_out_5_2_5[2:0]), //i
    .port_o (majority_5989_port_o                )  //o
  );
  Majority majority_5990 (
    .port_i (mixColumns_port_state_out_6_2_5[2:0]), //i
    .port_o (majority_5990_port_o                )  //o
  );
  Majority majority_5991 (
    .port_i (mixColumns_port_state_out_7_2_5[2:0]), //i
    .port_o (majority_5991_port_o                )  //o
  );
  Majority majority_5992 (
    .port_i (mixColumns_port_state_out_8_2_5[2:0]), //i
    .port_o (majority_5992_port_o                )  //o
  );
  Majority majority_5993 (
    .port_i (mixColumns_port_state_out_9_2_5[2:0]), //i
    .port_o (majority_5993_port_o                )  //o
  );
  Majority majority_5994 (
    .port_i (mixColumns_port_state_out_10_2_5[2:0]), //i
    .port_o (majority_5994_port_o                 )  //o
  );
  Majority majority_5995 (
    .port_i (mixColumns_port_state_out_11_2_5[2:0]), //i
    .port_o (majority_5995_port_o                 )  //o
  );
  Majority majority_5996 (
    .port_i (mixColumns_port_state_out_12_2_5[2:0]), //i
    .port_o (majority_5996_port_o                 )  //o
  );
  Majority majority_5997 (
    .port_i (mixColumns_port_state_out_13_2_5[2:0]), //i
    .port_o (majority_5997_port_o                 )  //o
  );
  Majority majority_5998 (
    .port_i (mixColumns_port_state_out_14_2_5[2:0]), //i
    .port_o (majority_5998_port_o                 )  //o
  );
  Majority majority_5999 (
    .port_i (mixColumns_port_state_out_15_2_5[2:0]), //i
    .port_o (majority_5999_port_o                 )  //o
  );
  Majority majority_6000 (
    .port_i (mixColumns_port_state_out_0_3_5[2:0]), //i
    .port_o (majority_6000_port_o                )  //o
  );
  Majority majority_6001 (
    .port_i (mixColumns_port_state_out_1_3_5[2:0]), //i
    .port_o (majority_6001_port_o                )  //o
  );
  Majority majority_6002 (
    .port_i (mixColumns_port_state_out_2_3_5[2:0]), //i
    .port_o (majority_6002_port_o                )  //o
  );
  Majority majority_6003 (
    .port_i (mixColumns_port_state_out_3_3_5[2:0]), //i
    .port_o (majority_6003_port_o                )  //o
  );
  Majority majority_6004 (
    .port_i (mixColumns_port_state_out_4_3_5[2:0]), //i
    .port_o (majority_6004_port_o                )  //o
  );
  Majority majority_6005 (
    .port_i (mixColumns_port_state_out_5_3_5[2:0]), //i
    .port_o (majority_6005_port_o                )  //o
  );
  Majority majority_6006 (
    .port_i (mixColumns_port_state_out_6_3_5[2:0]), //i
    .port_o (majority_6006_port_o                )  //o
  );
  Majority majority_6007 (
    .port_i (mixColumns_port_state_out_7_3_5[2:0]), //i
    .port_o (majority_6007_port_o                )  //o
  );
  Majority majority_6008 (
    .port_i (mixColumns_port_state_out_8_3_5[2:0]), //i
    .port_o (majority_6008_port_o                )  //o
  );
  Majority majority_6009 (
    .port_i (mixColumns_port_state_out_9_3_5[2:0]), //i
    .port_o (majority_6009_port_o                )  //o
  );
  Majority majority_6010 (
    .port_i (mixColumns_port_state_out_10_3_5[2:0]), //i
    .port_o (majority_6010_port_o                 )  //o
  );
  Majority majority_6011 (
    .port_i (mixColumns_port_state_out_11_3_5[2:0]), //i
    .port_o (majority_6011_port_o                 )  //o
  );
  Majority majority_6012 (
    .port_i (mixColumns_port_state_out_12_3_5[2:0]), //i
    .port_o (majority_6012_port_o                 )  //o
  );
  Majority majority_6013 (
    .port_i (mixColumns_port_state_out_13_3_5[2:0]), //i
    .port_o (majority_6013_port_o                 )  //o
  );
  Majority majority_6014 (
    .port_i (mixColumns_port_state_out_14_3_5[2:0]), //i
    .port_o (majority_6014_port_o                 )  //o
  );
  Majority majority_6015 (
    .port_i (mixColumns_port_state_out_15_3_5[2:0]), //i
    .port_o (majority_6015_port_o                 )  //o
  );
  Majority majority_6016 (
    .port_i (mixColumns_port_state_out_0_0_6[2:0]), //i
    .port_o (majority_6016_port_o                )  //o
  );
  Majority majority_6017 (
    .port_i (mixColumns_port_state_out_1_0_6[2:0]), //i
    .port_o (majority_6017_port_o                )  //o
  );
  Majority majority_6018 (
    .port_i (mixColumns_port_state_out_2_0_6[2:0]), //i
    .port_o (majority_6018_port_o                )  //o
  );
  Majority majority_6019 (
    .port_i (mixColumns_port_state_out_3_0_6[2:0]), //i
    .port_o (majority_6019_port_o                )  //o
  );
  Majority majority_6020 (
    .port_i (mixColumns_port_state_out_4_0_6[2:0]), //i
    .port_o (majority_6020_port_o                )  //o
  );
  Majority majority_6021 (
    .port_i (mixColumns_port_state_out_5_0_6[2:0]), //i
    .port_o (majority_6021_port_o                )  //o
  );
  Majority majority_6022 (
    .port_i (mixColumns_port_state_out_6_0_6[2:0]), //i
    .port_o (majority_6022_port_o                )  //o
  );
  Majority majority_6023 (
    .port_i (mixColumns_port_state_out_7_0_6[2:0]), //i
    .port_o (majority_6023_port_o                )  //o
  );
  Majority majority_6024 (
    .port_i (mixColumns_port_state_out_8_0_6[2:0]), //i
    .port_o (majority_6024_port_o                )  //o
  );
  Majority majority_6025 (
    .port_i (mixColumns_port_state_out_9_0_6[2:0]), //i
    .port_o (majority_6025_port_o                )  //o
  );
  Majority majority_6026 (
    .port_i (mixColumns_port_state_out_10_0_6[2:0]), //i
    .port_o (majority_6026_port_o                 )  //o
  );
  Majority majority_6027 (
    .port_i (mixColumns_port_state_out_11_0_6[2:0]), //i
    .port_o (majority_6027_port_o                 )  //o
  );
  Majority majority_6028 (
    .port_i (mixColumns_port_state_out_12_0_6[2:0]), //i
    .port_o (majority_6028_port_o                 )  //o
  );
  Majority majority_6029 (
    .port_i (mixColumns_port_state_out_13_0_6[2:0]), //i
    .port_o (majority_6029_port_o                 )  //o
  );
  Majority majority_6030 (
    .port_i (mixColumns_port_state_out_14_0_6[2:0]), //i
    .port_o (majority_6030_port_o                 )  //o
  );
  Majority majority_6031 (
    .port_i (mixColumns_port_state_out_15_0_6[2:0]), //i
    .port_o (majority_6031_port_o                 )  //o
  );
  Majority majority_6032 (
    .port_i (mixColumns_port_state_out_0_1_6[2:0]), //i
    .port_o (majority_6032_port_o                )  //o
  );
  Majority majority_6033 (
    .port_i (mixColumns_port_state_out_1_1_6[2:0]), //i
    .port_o (majority_6033_port_o                )  //o
  );
  Majority majority_6034 (
    .port_i (mixColumns_port_state_out_2_1_6[2:0]), //i
    .port_o (majority_6034_port_o                )  //o
  );
  Majority majority_6035 (
    .port_i (mixColumns_port_state_out_3_1_6[2:0]), //i
    .port_o (majority_6035_port_o                )  //o
  );
  Majority majority_6036 (
    .port_i (mixColumns_port_state_out_4_1_6[2:0]), //i
    .port_o (majority_6036_port_o                )  //o
  );
  Majority majority_6037 (
    .port_i (mixColumns_port_state_out_5_1_6[2:0]), //i
    .port_o (majority_6037_port_o                )  //o
  );
  Majority majority_6038 (
    .port_i (mixColumns_port_state_out_6_1_6[2:0]), //i
    .port_o (majority_6038_port_o                )  //o
  );
  Majority majority_6039 (
    .port_i (mixColumns_port_state_out_7_1_6[2:0]), //i
    .port_o (majority_6039_port_o                )  //o
  );
  Majority majority_6040 (
    .port_i (mixColumns_port_state_out_8_1_6[2:0]), //i
    .port_o (majority_6040_port_o                )  //o
  );
  Majority majority_6041 (
    .port_i (mixColumns_port_state_out_9_1_6[2:0]), //i
    .port_o (majority_6041_port_o                )  //o
  );
  Majority majority_6042 (
    .port_i (mixColumns_port_state_out_10_1_6[2:0]), //i
    .port_o (majority_6042_port_o                 )  //o
  );
  Majority majority_6043 (
    .port_i (mixColumns_port_state_out_11_1_6[2:0]), //i
    .port_o (majority_6043_port_o                 )  //o
  );
  Majority majority_6044 (
    .port_i (mixColumns_port_state_out_12_1_6[2:0]), //i
    .port_o (majority_6044_port_o                 )  //o
  );
  Majority majority_6045 (
    .port_i (mixColumns_port_state_out_13_1_6[2:0]), //i
    .port_o (majority_6045_port_o                 )  //o
  );
  Majority majority_6046 (
    .port_i (mixColumns_port_state_out_14_1_6[2:0]), //i
    .port_o (majority_6046_port_o                 )  //o
  );
  Majority majority_6047 (
    .port_i (mixColumns_port_state_out_15_1_6[2:0]), //i
    .port_o (majority_6047_port_o                 )  //o
  );
  Majority majority_6048 (
    .port_i (mixColumns_port_state_out_0_2_6[2:0]), //i
    .port_o (majority_6048_port_o                )  //o
  );
  Majority majority_6049 (
    .port_i (mixColumns_port_state_out_1_2_6[2:0]), //i
    .port_o (majority_6049_port_o                )  //o
  );
  Majority majority_6050 (
    .port_i (mixColumns_port_state_out_2_2_6[2:0]), //i
    .port_o (majority_6050_port_o                )  //o
  );
  Majority majority_6051 (
    .port_i (mixColumns_port_state_out_3_2_6[2:0]), //i
    .port_o (majority_6051_port_o                )  //o
  );
  Majority majority_6052 (
    .port_i (mixColumns_port_state_out_4_2_6[2:0]), //i
    .port_o (majority_6052_port_o                )  //o
  );
  Majority majority_6053 (
    .port_i (mixColumns_port_state_out_5_2_6[2:0]), //i
    .port_o (majority_6053_port_o                )  //o
  );
  Majority majority_6054 (
    .port_i (mixColumns_port_state_out_6_2_6[2:0]), //i
    .port_o (majority_6054_port_o                )  //o
  );
  Majority majority_6055 (
    .port_i (mixColumns_port_state_out_7_2_6[2:0]), //i
    .port_o (majority_6055_port_o                )  //o
  );
  Majority majority_6056 (
    .port_i (mixColumns_port_state_out_8_2_6[2:0]), //i
    .port_o (majority_6056_port_o                )  //o
  );
  Majority majority_6057 (
    .port_i (mixColumns_port_state_out_9_2_6[2:0]), //i
    .port_o (majority_6057_port_o                )  //o
  );
  Majority majority_6058 (
    .port_i (mixColumns_port_state_out_10_2_6[2:0]), //i
    .port_o (majority_6058_port_o                 )  //o
  );
  Majority majority_6059 (
    .port_i (mixColumns_port_state_out_11_2_6[2:0]), //i
    .port_o (majority_6059_port_o                 )  //o
  );
  Majority majority_6060 (
    .port_i (mixColumns_port_state_out_12_2_6[2:0]), //i
    .port_o (majority_6060_port_o                 )  //o
  );
  Majority majority_6061 (
    .port_i (mixColumns_port_state_out_13_2_6[2:0]), //i
    .port_o (majority_6061_port_o                 )  //o
  );
  Majority majority_6062 (
    .port_i (mixColumns_port_state_out_14_2_6[2:0]), //i
    .port_o (majority_6062_port_o                 )  //o
  );
  Majority majority_6063 (
    .port_i (mixColumns_port_state_out_15_2_6[2:0]), //i
    .port_o (majority_6063_port_o                 )  //o
  );
  Majority majority_6064 (
    .port_i (mixColumns_port_state_out_0_3_6[2:0]), //i
    .port_o (majority_6064_port_o                )  //o
  );
  Majority majority_6065 (
    .port_i (mixColumns_port_state_out_1_3_6[2:0]), //i
    .port_o (majority_6065_port_o                )  //o
  );
  Majority majority_6066 (
    .port_i (mixColumns_port_state_out_2_3_6[2:0]), //i
    .port_o (majority_6066_port_o                )  //o
  );
  Majority majority_6067 (
    .port_i (mixColumns_port_state_out_3_3_6[2:0]), //i
    .port_o (majority_6067_port_o                )  //o
  );
  Majority majority_6068 (
    .port_i (mixColumns_port_state_out_4_3_6[2:0]), //i
    .port_o (majority_6068_port_o                )  //o
  );
  Majority majority_6069 (
    .port_i (mixColumns_port_state_out_5_3_6[2:0]), //i
    .port_o (majority_6069_port_o                )  //o
  );
  Majority majority_6070 (
    .port_i (mixColumns_port_state_out_6_3_6[2:0]), //i
    .port_o (majority_6070_port_o                )  //o
  );
  Majority majority_6071 (
    .port_i (mixColumns_port_state_out_7_3_6[2:0]), //i
    .port_o (majority_6071_port_o                )  //o
  );
  Majority majority_6072 (
    .port_i (mixColumns_port_state_out_8_3_6[2:0]), //i
    .port_o (majority_6072_port_o                )  //o
  );
  Majority majority_6073 (
    .port_i (mixColumns_port_state_out_9_3_6[2:0]), //i
    .port_o (majority_6073_port_o                )  //o
  );
  Majority majority_6074 (
    .port_i (mixColumns_port_state_out_10_3_6[2:0]), //i
    .port_o (majority_6074_port_o                 )  //o
  );
  Majority majority_6075 (
    .port_i (mixColumns_port_state_out_11_3_6[2:0]), //i
    .port_o (majority_6075_port_o                 )  //o
  );
  Majority majority_6076 (
    .port_i (mixColumns_port_state_out_12_3_6[2:0]), //i
    .port_o (majority_6076_port_o                 )  //o
  );
  Majority majority_6077 (
    .port_i (mixColumns_port_state_out_13_3_6[2:0]), //i
    .port_o (majority_6077_port_o                 )  //o
  );
  Majority majority_6078 (
    .port_i (mixColumns_port_state_out_14_3_6[2:0]), //i
    .port_o (majority_6078_port_o                 )  //o
  );
  Majority majority_6079 (
    .port_i (mixColumns_port_state_out_15_3_6[2:0]), //i
    .port_o (majority_6079_port_o                 )  //o
  );
  Majority majority_6080 (
    .port_i (mixColumns_port_state_out_0_0_7[2:0]), //i
    .port_o (majority_6080_port_o                )  //o
  );
  Majority majority_6081 (
    .port_i (mixColumns_port_state_out_1_0_7[2:0]), //i
    .port_o (majority_6081_port_o                )  //o
  );
  Majority majority_6082 (
    .port_i (mixColumns_port_state_out_2_0_7[2:0]), //i
    .port_o (majority_6082_port_o                )  //o
  );
  Majority majority_6083 (
    .port_i (mixColumns_port_state_out_3_0_7[2:0]), //i
    .port_o (majority_6083_port_o                )  //o
  );
  Majority majority_6084 (
    .port_i (mixColumns_port_state_out_4_0_7[2:0]), //i
    .port_o (majority_6084_port_o                )  //o
  );
  Majority majority_6085 (
    .port_i (mixColumns_port_state_out_5_0_7[2:0]), //i
    .port_o (majority_6085_port_o                )  //o
  );
  Majority majority_6086 (
    .port_i (mixColumns_port_state_out_6_0_7[2:0]), //i
    .port_o (majority_6086_port_o                )  //o
  );
  Majority majority_6087 (
    .port_i (mixColumns_port_state_out_7_0_7[2:0]), //i
    .port_o (majority_6087_port_o                )  //o
  );
  Majority majority_6088 (
    .port_i (mixColumns_port_state_out_8_0_7[2:0]), //i
    .port_o (majority_6088_port_o                )  //o
  );
  Majority majority_6089 (
    .port_i (mixColumns_port_state_out_9_0_7[2:0]), //i
    .port_o (majority_6089_port_o                )  //o
  );
  Majority majority_6090 (
    .port_i (mixColumns_port_state_out_10_0_7[2:0]), //i
    .port_o (majority_6090_port_o                 )  //o
  );
  Majority majority_6091 (
    .port_i (mixColumns_port_state_out_11_0_7[2:0]), //i
    .port_o (majority_6091_port_o                 )  //o
  );
  Majority majority_6092 (
    .port_i (mixColumns_port_state_out_12_0_7[2:0]), //i
    .port_o (majority_6092_port_o                 )  //o
  );
  Majority majority_6093 (
    .port_i (mixColumns_port_state_out_13_0_7[2:0]), //i
    .port_o (majority_6093_port_o                 )  //o
  );
  Majority majority_6094 (
    .port_i (mixColumns_port_state_out_14_0_7[2:0]), //i
    .port_o (majority_6094_port_o                 )  //o
  );
  Majority majority_6095 (
    .port_i (mixColumns_port_state_out_15_0_7[2:0]), //i
    .port_o (majority_6095_port_o                 )  //o
  );
  Majority majority_6096 (
    .port_i (mixColumns_port_state_out_0_1_7[2:0]), //i
    .port_o (majority_6096_port_o                )  //o
  );
  Majority majority_6097 (
    .port_i (mixColumns_port_state_out_1_1_7[2:0]), //i
    .port_o (majority_6097_port_o                )  //o
  );
  Majority majority_6098 (
    .port_i (mixColumns_port_state_out_2_1_7[2:0]), //i
    .port_o (majority_6098_port_o                )  //o
  );
  Majority majority_6099 (
    .port_i (mixColumns_port_state_out_3_1_7[2:0]), //i
    .port_o (majority_6099_port_o                )  //o
  );
  Majority majority_6100 (
    .port_i (mixColumns_port_state_out_4_1_7[2:0]), //i
    .port_o (majority_6100_port_o                )  //o
  );
  Majority majority_6101 (
    .port_i (mixColumns_port_state_out_5_1_7[2:0]), //i
    .port_o (majority_6101_port_o                )  //o
  );
  Majority majority_6102 (
    .port_i (mixColumns_port_state_out_6_1_7[2:0]), //i
    .port_o (majority_6102_port_o                )  //o
  );
  Majority majority_6103 (
    .port_i (mixColumns_port_state_out_7_1_7[2:0]), //i
    .port_o (majority_6103_port_o                )  //o
  );
  Majority majority_6104 (
    .port_i (mixColumns_port_state_out_8_1_7[2:0]), //i
    .port_o (majority_6104_port_o                )  //o
  );
  Majority majority_6105 (
    .port_i (mixColumns_port_state_out_9_1_7[2:0]), //i
    .port_o (majority_6105_port_o                )  //o
  );
  Majority majority_6106 (
    .port_i (mixColumns_port_state_out_10_1_7[2:0]), //i
    .port_o (majority_6106_port_o                 )  //o
  );
  Majority majority_6107 (
    .port_i (mixColumns_port_state_out_11_1_7[2:0]), //i
    .port_o (majority_6107_port_o                 )  //o
  );
  Majority majority_6108 (
    .port_i (mixColumns_port_state_out_12_1_7[2:0]), //i
    .port_o (majority_6108_port_o                 )  //o
  );
  Majority majority_6109 (
    .port_i (mixColumns_port_state_out_13_1_7[2:0]), //i
    .port_o (majority_6109_port_o                 )  //o
  );
  Majority majority_6110 (
    .port_i (mixColumns_port_state_out_14_1_7[2:0]), //i
    .port_o (majority_6110_port_o                 )  //o
  );
  Majority majority_6111 (
    .port_i (mixColumns_port_state_out_15_1_7[2:0]), //i
    .port_o (majority_6111_port_o                 )  //o
  );
  Majority majority_6112 (
    .port_i (mixColumns_port_state_out_0_2_7[2:0]), //i
    .port_o (majority_6112_port_o                )  //o
  );
  Majority majority_6113 (
    .port_i (mixColumns_port_state_out_1_2_7[2:0]), //i
    .port_o (majority_6113_port_o                )  //o
  );
  Majority majority_6114 (
    .port_i (mixColumns_port_state_out_2_2_7[2:0]), //i
    .port_o (majority_6114_port_o                )  //o
  );
  Majority majority_6115 (
    .port_i (mixColumns_port_state_out_3_2_7[2:0]), //i
    .port_o (majority_6115_port_o                )  //o
  );
  Majority majority_6116 (
    .port_i (mixColumns_port_state_out_4_2_7[2:0]), //i
    .port_o (majority_6116_port_o                )  //o
  );
  Majority majority_6117 (
    .port_i (mixColumns_port_state_out_5_2_7[2:0]), //i
    .port_o (majority_6117_port_o                )  //o
  );
  Majority majority_6118 (
    .port_i (mixColumns_port_state_out_6_2_7[2:0]), //i
    .port_o (majority_6118_port_o                )  //o
  );
  Majority majority_6119 (
    .port_i (mixColumns_port_state_out_7_2_7[2:0]), //i
    .port_o (majority_6119_port_o                )  //o
  );
  Majority majority_6120 (
    .port_i (mixColumns_port_state_out_8_2_7[2:0]), //i
    .port_o (majority_6120_port_o                )  //o
  );
  Majority majority_6121 (
    .port_i (mixColumns_port_state_out_9_2_7[2:0]), //i
    .port_o (majority_6121_port_o                )  //o
  );
  Majority majority_6122 (
    .port_i (mixColumns_port_state_out_10_2_7[2:0]), //i
    .port_o (majority_6122_port_o                 )  //o
  );
  Majority majority_6123 (
    .port_i (mixColumns_port_state_out_11_2_7[2:0]), //i
    .port_o (majority_6123_port_o                 )  //o
  );
  Majority majority_6124 (
    .port_i (mixColumns_port_state_out_12_2_7[2:0]), //i
    .port_o (majority_6124_port_o                 )  //o
  );
  Majority majority_6125 (
    .port_i (mixColumns_port_state_out_13_2_7[2:0]), //i
    .port_o (majority_6125_port_o                 )  //o
  );
  Majority majority_6126 (
    .port_i (mixColumns_port_state_out_14_2_7[2:0]), //i
    .port_o (majority_6126_port_o                 )  //o
  );
  Majority majority_6127 (
    .port_i (mixColumns_port_state_out_15_2_7[2:0]), //i
    .port_o (majority_6127_port_o                 )  //o
  );
  Majority majority_6128 (
    .port_i (mixColumns_port_state_out_0_3_7[2:0]), //i
    .port_o (majority_6128_port_o                )  //o
  );
  Majority majority_6129 (
    .port_i (mixColumns_port_state_out_1_3_7[2:0]), //i
    .port_o (majority_6129_port_o                )  //o
  );
  Majority majority_6130 (
    .port_i (mixColumns_port_state_out_2_3_7[2:0]), //i
    .port_o (majority_6130_port_o                )  //o
  );
  Majority majority_6131 (
    .port_i (mixColumns_port_state_out_3_3_7[2:0]), //i
    .port_o (majority_6131_port_o                )  //o
  );
  Majority majority_6132 (
    .port_i (mixColumns_port_state_out_4_3_7[2:0]), //i
    .port_o (majority_6132_port_o                )  //o
  );
  Majority majority_6133 (
    .port_i (mixColumns_port_state_out_5_3_7[2:0]), //i
    .port_o (majority_6133_port_o                )  //o
  );
  Majority majority_6134 (
    .port_i (mixColumns_port_state_out_6_3_7[2:0]), //i
    .port_o (majority_6134_port_o                )  //o
  );
  Majority majority_6135 (
    .port_i (mixColumns_port_state_out_7_3_7[2:0]), //i
    .port_o (majority_6135_port_o                )  //o
  );
  Majority majority_6136 (
    .port_i (mixColumns_port_state_out_8_3_7[2:0]), //i
    .port_o (majority_6136_port_o                )  //o
  );
  Majority majority_6137 (
    .port_i (mixColumns_port_state_out_9_3_7[2:0]), //i
    .port_o (majority_6137_port_o                )  //o
  );
  Majority majority_6138 (
    .port_i (mixColumns_port_state_out_10_3_7[2:0]), //i
    .port_o (majority_6138_port_o                 )  //o
  );
  Majority majority_6139 (
    .port_i (mixColumns_port_state_out_11_3_7[2:0]), //i
    .port_o (majority_6139_port_o                 )  //o
  );
  Majority majority_6140 (
    .port_i (mixColumns_port_state_out_12_3_7[2:0]), //i
    .port_o (majority_6140_port_o                 )  //o
  );
  Majority majority_6141 (
    .port_i (mixColumns_port_state_out_13_3_7[2:0]), //i
    .port_o (majority_6141_port_o                 )  //o
  );
  Majority majority_6142 (
    .port_i (mixColumns_port_state_out_14_3_7[2:0]), //i
    .port_o (majority_6142_port_o                 )  //o
  );
  Majority majority_6143 (
    .port_i (mixColumns_port_state_out_15_3_7[2:0]), //i
    .port_o (majority_6143_port_o                 )  //o
  );
  assign subBytes_out_0_0_0 = sbox_AES_BoyarPeralta_16_port_o_0_0;
  assign subBytes_out_0_0_1 = sbox_AES_BoyarPeralta_16_port_o_0_1;
  assign subBytes_out_0_0_2 = sbox_AES_BoyarPeralta_16_port_o_0_2;
  assign subBytes_out_0_0_3 = sbox_AES_BoyarPeralta_16_port_o_0_3;
  assign subBytes_out_0_0_4 = sbox_AES_BoyarPeralta_16_port_o_0_4;
  assign subBytes_out_0_0_5 = sbox_AES_BoyarPeralta_16_port_o_0_5;
  assign subBytes_out_0_0_6 = sbox_AES_BoyarPeralta_16_port_o_0_6;
  assign subBytes_out_0_0_7 = sbox_AES_BoyarPeralta_16_port_o_0_7;
  assign subBytes_out_0_1_0 = sbox_AES_BoyarPeralta_16_port_o_1_0;
  assign subBytes_out_0_1_1 = sbox_AES_BoyarPeralta_16_port_o_1_1;
  assign subBytes_out_0_1_2 = sbox_AES_BoyarPeralta_16_port_o_1_2;
  assign subBytes_out_0_1_3 = sbox_AES_BoyarPeralta_16_port_o_1_3;
  assign subBytes_out_0_1_4 = sbox_AES_BoyarPeralta_16_port_o_1_4;
  assign subBytes_out_0_1_5 = sbox_AES_BoyarPeralta_16_port_o_1_5;
  assign subBytes_out_0_1_6 = sbox_AES_BoyarPeralta_16_port_o_1_6;
  assign subBytes_out_0_1_7 = sbox_AES_BoyarPeralta_16_port_o_1_7;
  assign subBytes_out_0_2_0 = sbox_AES_BoyarPeralta_16_port_o_2_0;
  assign subBytes_out_0_2_1 = sbox_AES_BoyarPeralta_16_port_o_2_1;
  assign subBytes_out_0_2_2 = sbox_AES_BoyarPeralta_16_port_o_2_2;
  assign subBytes_out_0_2_3 = sbox_AES_BoyarPeralta_16_port_o_2_3;
  assign subBytes_out_0_2_4 = sbox_AES_BoyarPeralta_16_port_o_2_4;
  assign subBytes_out_0_2_5 = sbox_AES_BoyarPeralta_16_port_o_2_5;
  assign subBytes_out_0_2_6 = sbox_AES_BoyarPeralta_16_port_o_2_6;
  assign subBytes_out_0_2_7 = sbox_AES_BoyarPeralta_16_port_o_2_7;
  assign subBytes_out_0_3_0 = sbox_AES_BoyarPeralta_16_port_o_3_0;
  assign subBytes_out_0_3_1 = sbox_AES_BoyarPeralta_16_port_o_3_1;
  assign subBytes_out_0_3_2 = sbox_AES_BoyarPeralta_16_port_o_3_2;
  assign subBytes_out_0_3_3 = sbox_AES_BoyarPeralta_16_port_o_3_3;
  assign subBytes_out_0_3_4 = sbox_AES_BoyarPeralta_16_port_o_3_4;
  assign subBytes_out_0_3_5 = sbox_AES_BoyarPeralta_16_port_o_3_5;
  assign subBytes_out_0_3_6 = sbox_AES_BoyarPeralta_16_port_o_3_6;
  assign subBytes_out_0_3_7 = sbox_AES_BoyarPeralta_16_port_o_3_7;
  assign subBytes_out_1_0_0 = sbox_AES_BoyarPeralta_17_port_o_0_0;
  assign subBytes_out_1_0_1 = sbox_AES_BoyarPeralta_17_port_o_0_1;
  assign subBytes_out_1_0_2 = sbox_AES_BoyarPeralta_17_port_o_0_2;
  assign subBytes_out_1_0_3 = sbox_AES_BoyarPeralta_17_port_o_0_3;
  assign subBytes_out_1_0_4 = sbox_AES_BoyarPeralta_17_port_o_0_4;
  assign subBytes_out_1_0_5 = sbox_AES_BoyarPeralta_17_port_o_0_5;
  assign subBytes_out_1_0_6 = sbox_AES_BoyarPeralta_17_port_o_0_6;
  assign subBytes_out_1_0_7 = sbox_AES_BoyarPeralta_17_port_o_0_7;
  assign subBytes_out_1_1_0 = sbox_AES_BoyarPeralta_17_port_o_1_0;
  assign subBytes_out_1_1_1 = sbox_AES_BoyarPeralta_17_port_o_1_1;
  assign subBytes_out_1_1_2 = sbox_AES_BoyarPeralta_17_port_o_1_2;
  assign subBytes_out_1_1_3 = sbox_AES_BoyarPeralta_17_port_o_1_3;
  assign subBytes_out_1_1_4 = sbox_AES_BoyarPeralta_17_port_o_1_4;
  assign subBytes_out_1_1_5 = sbox_AES_BoyarPeralta_17_port_o_1_5;
  assign subBytes_out_1_1_6 = sbox_AES_BoyarPeralta_17_port_o_1_6;
  assign subBytes_out_1_1_7 = sbox_AES_BoyarPeralta_17_port_o_1_7;
  assign subBytes_out_1_2_0 = sbox_AES_BoyarPeralta_17_port_o_2_0;
  assign subBytes_out_1_2_1 = sbox_AES_BoyarPeralta_17_port_o_2_1;
  assign subBytes_out_1_2_2 = sbox_AES_BoyarPeralta_17_port_o_2_2;
  assign subBytes_out_1_2_3 = sbox_AES_BoyarPeralta_17_port_o_2_3;
  assign subBytes_out_1_2_4 = sbox_AES_BoyarPeralta_17_port_o_2_4;
  assign subBytes_out_1_2_5 = sbox_AES_BoyarPeralta_17_port_o_2_5;
  assign subBytes_out_1_2_6 = sbox_AES_BoyarPeralta_17_port_o_2_6;
  assign subBytes_out_1_2_7 = sbox_AES_BoyarPeralta_17_port_o_2_7;
  assign subBytes_out_1_3_0 = sbox_AES_BoyarPeralta_17_port_o_3_0;
  assign subBytes_out_1_3_1 = sbox_AES_BoyarPeralta_17_port_o_3_1;
  assign subBytes_out_1_3_2 = sbox_AES_BoyarPeralta_17_port_o_3_2;
  assign subBytes_out_1_3_3 = sbox_AES_BoyarPeralta_17_port_o_3_3;
  assign subBytes_out_1_3_4 = sbox_AES_BoyarPeralta_17_port_o_3_4;
  assign subBytes_out_1_3_5 = sbox_AES_BoyarPeralta_17_port_o_3_5;
  assign subBytes_out_1_3_6 = sbox_AES_BoyarPeralta_17_port_o_3_6;
  assign subBytes_out_1_3_7 = sbox_AES_BoyarPeralta_17_port_o_3_7;
  assign subBytes_out_2_0_0 = sbox_AES_BoyarPeralta_18_port_o_0_0;
  assign subBytes_out_2_0_1 = sbox_AES_BoyarPeralta_18_port_o_0_1;
  assign subBytes_out_2_0_2 = sbox_AES_BoyarPeralta_18_port_o_0_2;
  assign subBytes_out_2_0_3 = sbox_AES_BoyarPeralta_18_port_o_0_3;
  assign subBytes_out_2_0_4 = sbox_AES_BoyarPeralta_18_port_o_0_4;
  assign subBytes_out_2_0_5 = sbox_AES_BoyarPeralta_18_port_o_0_5;
  assign subBytes_out_2_0_6 = sbox_AES_BoyarPeralta_18_port_o_0_6;
  assign subBytes_out_2_0_7 = sbox_AES_BoyarPeralta_18_port_o_0_7;
  assign subBytes_out_2_1_0 = sbox_AES_BoyarPeralta_18_port_o_1_0;
  assign subBytes_out_2_1_1 = sbox_AES_BoyarPeralta_18_port_o_1_1;
  assign subBytes_out_2_1_2 = sbox_AES_BoyarPeralta_18_port_o_1_2;
  assign subBytes_out_2_1_3 = sbox_AES_BoyarPeralta_18_port_o_1_3;
  assign subBytes_out_2_1_4 = sbox_AES_BoyarPeralta_18_port_o_1_4;
  assign subBytes_out_2_1_5 = sbox_AES_BoyarPeralta_18_port_o_1_5;
  assign subBytes_out_2_1_6 = sbox_AES_BoyarPeralta_18_port_o_1_6;
  assign subBytes_out_2_1_7 = sbox_AES_BoyarPeralta_18_port_o_1_7;
  assign subBytes_out_2_2_0 = sbox_AES_BoyarPeralta_18_port_o_2_0;
  assign subBytes_out_2_2_1 = sbox_AES_BoyarPeralta_18_port_o_2_1;
  assign subBytes_out_2_2_2 = sbox_AES_BoyarPeralta_18_port_o_2_2;
  assign subBytes_out_2_2_3 = sbox_AES_BoyarPeralta_18_port_o_2_3;
  assign subBytes_out_2_2_4 = sbox_AES_BoyarPeralta_18_port_o_2_4;
  assign subBytes_out_2_2_5 = sbox_AES_BoyarPeralta_18_port_o_2_5;
  assign subBytes_out_2_2_6 = sbox_AES_BoyarPeralta_18_port_o_2_6;
  assign subBytes_out_2_2_7 = sbox_AES_BoyarPeralta_18_port_o_2_7;
  assign subBytes_out_2_3_0 = sbox_AES_BoyarPeralta_18_port_o_3_0;
  assign subBytes_out_2_3_1 = sbox_AES_BoyarPeralta_18_port_o_3_1;
  assign subBytes_out_2_3_2 = sbox_AES_BoyarPeralta_18_port_o_3_2;
  assign subBytes_out_2_3_3 = sbox_AES_BoyarPeralta_18_port_o_3_3;
  assign subBytes_out_2_3_4 = sbox_AES_BoyarPeralta_18_port_o_3_4;
  assign subBytes_out_2_3_5 = sbox_AES_BoyarPeralta_18_port_o_3_5;
  assign subBytes_out_2_3_6 = sbox_AES_BoyarPeralta_18_port_o_3_6;
  assign subBytes_out_2_3_7 = sbox_AES_BoyarPeralta_18_port_o_3_7;
  assign subBytes_out_3_0_0 = sbox_AES_BoyarPeralta_19_port_o_0_0;
  assign subBytes_out_3_0_1 = sbox_AES_BoyarPeralta_19_port_o_0_1;
  assign subBytes_out_3_0_2 = sbox_AES_BoyarPeralta_19_port_o_0_2;
  assign subBytes_out_3_0_3 = sbox_AES_BoyarPeralta_19_port_o_0_3;
  assign subBytes_out_3_0_4 = sbox_AES_BoyarPeralta_19_port_o_0_4;
  assign subBytes_out_3_0_5 = sbox_AES_BoyarPeralta_19_port_o_0_5;
  assign subBytes_out_3_0_6 = sbox_AES_BoyarPeralta_19_port_o_0_6;
  assign subBytes_out_3_0_7 = sbox_AES_BoyarPeralta_19_port_o_0_7;
  assign subBytes_out_3_1_0 = sbox_AES_BoyarPeralta_19_port_o_1_0;
  assign subBytes_out_3_1_1 = sbox_AES_BoyarPeralta_19_port_o_1_1;
  assign subBytes_out_3_1_2 = sbox_AES_BoyarPeralta_19_port_o_1_2;
  assign subBytes_out_3_1_3 = sbox_AES_BoyarPeralta_19_port_o_1_3;
  assign subBytes_out_3_1_4 = sbox_AES_BoyarPeralta_19_port_o_1_4;
  assign subBytes_out_3_1_5 = sbox_AES_BoyarPeralta_19_port_o_1_5;
  assign subBytes_out_3_1_6 = sbox_AES_BoyarPeralta_19_port_o_1_6;
  assign subBytes_out_3_1_7 = sbox_AES_BoyarPeralta_19_port_o_1_7;
  assign subBytes_out_3_2_0 = sbox_AES_BoyarPeralta_19_port_o_2_0;
  assign subBytes_out_3_2_1 = sbox_AES_BoyarPeralta_19_port_o_2_1;
  assign subBytes_out_3_2_2 = sbox_AES_BoyarPeralta_19_port_o_2_2;
  assign subBytes_out_3_2_3 = sbox_AES_BoyarPeralta_19_port_o_2_3;
  assign subBytes_out_3_2_4 = sbox_AES_BoyarPeralta_19_port_o_2_4;
  assign subBytes_out_3_2_5 = sbox_AES_BoyarPeralta_19_port_o_2_5;
  assign subBytes_out_3_2_6 = sbox_AES_BoyarPeralta_19_port_o_2_6;
  assign subBytes_out_3_2_7 = sbox_AES_BoyarPeralta_19_port_o_2_7;
  assign subBytes_out_3_3_0 = sbox_AES_BoyarPeralta_19_port_o_3_0;
  assign subBytes_out_3_3_1 = sbox_AES_BoyarPeralta_19_port_o_3_1;
  assign subBytes_out_3_3_2 = sbox_AES_BoyarPeralta_19_port_o_3_2;
  assign subBytes_out_3_3_3 = sbox_AES_BoyarPeralta_19_port_o_3_3;
  assign subBytes_out_3_3_4 = sbox_AES_BoyarPeralta_19_port_o_3_4;
  assign subBytes_out_3_3_5 = sbox_AES_BoyarPeralta_19_port_o_3_5;
  assign subBytes_out_3_3_6 = sbox_AES_BoyarPeralta_19_port_o_3_6;
  assign subBytes_out_3_3_7 = sbox_AES_BoyarPeralta_19_port_o_3_7;
  assign subBytes_out_4_0_0 = sbox_AES_BoyarPeralta_20_port_o_0_0;
  assign subBytes_out_4_0_1 = sbox_AES_BoyarPeralta_20_port_o_0_1;
  assign subBytes_out_4_0_2 = sbox_AES_BoyarPeralta_20_port_o_0_2;
  assign subBytes_out_4_0_3 = sbox_AES_BoyarPeralta_20_port_o_0_3;
  assign subBytes_out_4_0_4 = sbox_AES_BoyarPeralta_20_port_o_0_4;
  assign subBytes_out_4_0_5 = sbox_AES_BoyarPeralta_20_port_o_0_5;
  assign subBytes_out_4_0_6 = sbox_AES_BoyarPeralta_20_port_o_0_6;
  assign subBytes_out_4_0_7 = sbox_AES_BoyarPeralta_20_port_o_0_7;
  assign subBytes_out_4_1_0 = sbox_AES_BoyarPeralta_20_port_o_1_0;
  assign subBytes_out_4_1_1 = sbox_AES_BoyarPeralta_20_port_o_1_1;
  assign subBytes_out_4_1_2 = sbox_AES_BoyarPeralta_20_port_o_1_2;
  assign subBytes_out_4_1_3 = sbox_AES_BoyarPeralta_20_port_o_1_3;
  assign subBytes_out_4_1_4 = sbox_AES_BoyarPeralta_20_port_o_1_4;
  assign subBytes_out_4_1_5 = sbox_AES_BoyarPeralta_20_port_o_1_5;
  assign subBytes_out_4_1_6 = sbox_AES_BoyarPeralta_20_port_o_1_6;
  assign subBytes_out_4_1_7 = sbox_AES_BoyarPeralta_20_port_o_1_7;
  assign subBytes_out_4_2_0 = sbox_AES_BoyarPeralta_20_port_o_2_0;
  assign subBytes_out_4_2_1 = sbox_AES_BoyarPeralta_20_port_o_2_1;
  assign subBytes_out_4_2_2 = sbox_AES_BoyarPeralta_20_port_o_2_2;
  assign subBytes_out_4_2_3 = sbox_AES_BoyarPeralta_20_port_o_2_3;
  assign subBytes_out_4_2_4 = sbox_AES_BoyarPeralta_20_port_o_2_4;
  assign subBytes_out_4_2_5 = sbox_AES_BoyarPeralta_20_port_o_2_5;
  assign subBytes_out_4_2_6 = sbox_AES_BoyarPeralta_20_port_o_2_6;
  assign subBytes_out_4_2_7 = sbox_AES_BoyarPeralta_20_port_o_2_7;
  assign subBytes_out_4_3_0 = sbox_AES_BoyarPeralta_20_port_o_3_0;
  assign subBytes_out_4_3_1 = sbox_AES_BoyarPeralta_20_port_o_3_1;
  assign subBytes_out_4_3_2 = sbox_AES_BoyarPeralta_20_port_o_3_2;
  assign subBytes_out_4_3_3 = sbox_AES_BoyarPeralta_20_port_o_3_3;
  assign subBytes_out_4_3_4 = sbox_AES_BoyarPeralta_20_port_o_3_4;
  assign subBytes_out_4_3_5 = sbox_AES_BoyarPeralta_20_port_o_3_5;
  assign subBytes_out_4_3_6 = sbox_AES_BoyarPeralta_20_port_o_3_6;
  assign subBytes_out_4_3_7 = sbox_AES_BoyarPeralta_20_port_o_3_7;
  assign subBytes_out_5_0_0 = sbox_AES_BoyarPeralta_21_port_o_0_0;
  assign subBytes_out_5_0_1 = sbox_AES_BoyarPeralta_21_port_o_0_1;
  assign subBytes_out_5_0_2 = sbox_AES_BoyarPeralta_21_port_o_0_2;
  assign subBytes_out_5_0_3 = sbox_AES_BoyarPeralta_21_port_o_0_3;
  assign subBytes_out_5_0_4 = sbox_AES_BoyarPeralta_21_port_o_0_4;
  assign subBytes_out_5_0_5 = sbox_AES_BoyarPeralta_21_port_o_0_5;
  assign subBytes_out_5_0_6 = sbox_AES_BoyarPeralta_21_port_o_0_6;
  assign subBytes_out_5_0_7 = sbox_AES_BoyarPeralta_21_port_o_0_7;
  assign subBytes_out_5_1_0 = sbox_AES_BoyarPeralta_21_port_o_1_0;
  assign subBytes_out_5_1_1 = sbox_AES_BoyarPeralta_21_port_o_1_1;
  assign subBytes_out_5_1_2 = sbox_AES_BoyarPeralta_21_port_o_1_2;
  assign subBytes_out_5_1_3 = sbox_AES_BoyarPeralta_21_port_o_1_3;
  assign subBytes_out_5_1_4 = sbox_AES_BoyarPeralta_21_port_o_1_4;
  assign subBytes_out_5_1_5 = sbox_AES_BoyarPeralta_21_port_o_1_5;
  assign subBytes_out_5_1_6 = sbox_AES_BoyarPeralta_21_port_o_1_6;
  assign subBytes_out_5_1_7 = sbox_AES_BoyarPeralta_21_port_o_1_7;
  assign subBytes_out_5_2_0 = sbox_AES_BoyarPeralta_21_port_o_2_0;
  assign subBytes_out_5_2_1 = sbox_AES_BoyarPeralta_21_port_o_2_1;
  assign subBytes_out_5_2_2 = sbox_AES_BoyarPeralta_21_port_o_2_2;
  assign subBytes_out_5_2_3 = sbox_AES_BoyarPeralta_21_port_o_2_3;
  assign subBytes_out_5_2_4 = sbox_AES_BoyarPeralta_21_port_o_2_4;
  assign subBytes_out_5_2_5 = sbox_AES_BoyarPeralta_21_port_o_2_5;
  assign subBytes_out_5_2_6 = sbox_AES_BoyarPeralta_21_port_o_2_6;
  assign subBytes_out_5_2_7 = sbox_AES_BoyarPeralta_21_port_o_2_7;
  assign subBytes_out_5_3_0 = sbox_AES_BoyarPeralta_21_port_o_3_0;
  assign subBytes_out_5_3_1 = sbox_AES_BoyarPeralta_21_port_o_3_1;
  assign subBytes_out_5_3_2 = sbox_AES_BoyarPeralta_21_port_o_3_2;
  assign subBytes_out_5_3_3 = sbox_AES_BoyarPeralta_21_port_o_3_3;
  assign subBytes_out_5_3_4 = sbox_AES_BoyarPeralta_21_port_o_3_4;
  assign subBytes_out_5_3_5 = sbox_AES_BoyarPeralta_21_port_o_3_5;
  assign subBytes_out_5_3_6 = sbox_AES_BoyarPeralta_21_port_o_3_6;
  assign subBytes_out_5_3_7 = sbox_AES_BoyarPeralta_21_port_o_3_7;
  assign subBytes_out_6_0_0 = sbox_AES_BoyarPeralta_22_port_o_0_0;
  assign subBytes_out_6_0_1 = sbox_AES_BoyarPeralta_22_port_o_0_1;
  assign subBytes_out_6_0_2 = sbox_AES_BoyarPeralta_22_port_o_0_2;
  assign subBytes_out_6_0_3 = sbox_AES_BoyarPeralta_22_port_o_0_3;
  assign subBytes_out_6_0_4 = sbox_AES_BoyarPeralta_22_port_o_0_4;
  assign subBytes_out_6_0_5 = sbox_AES_BoyarPeralta_22_port_o_0_5;
  assign subBytes_out_6_0_6 = sbox_AES_BoyarPeralta_22_port_o_0_6;
  assign subBytes_out_6_0_7 = sbox_AES_BoyarPeralta_22_port_o_0_7;
  assign subBytes_out_6_1_0 = sbox_AES_BoyarPeralta_22_port_o_1_0;
  assign subBytes_out_6_1_1 = sbox_AES_BoyarPeralta_22_port_o_1_1;
  assign subBytes_out_6_1_2 = sbox_AES_BoyarPeralta_22_port_o_1_2;
  assign subBytes_out_6_1_3 = sbox_AES_BoyarPeralta_22_port_o_1_3;
  assign subBytes_out_6_1_4 = sbox_AES_BoyarPeralta_22_port_o_1_4;
  assign subBytes_out_6_1_5 = sbox_AES_BoyarPeralta_22_port_o_1_5;
  assign subBytes_out_6_1_6 = sbox_AES_BoyarPeralta_22_port_o_1_6;
  assign subBytes_out_6_1_7 = sbox_AES_BoyarPeralta_22_port_o_1_7;
  assign subBytes_out_6_2_0 = sbox_AES_BoyarPeralta_22_port_o_2_0;
  assign subBytes_out_6_2_1 = sbox_AES_BoyarPeralta_22_port_o_2_1;
  assign subBytes_out_6_2_2 = sbox_AES_BoyarPeralta_22_port_o_2_2;
  assign subBytes_out_6_2_3 = sbox_AES_BoyarPeralta_22_port_o_2_3;
  assign subBytes_out_6_2_4 = sbox_AES_BoyarPeralta_22_port_o_2_4;
  assign subBytes_out_6_2_5 = sbox_AES_BoyarPeralta_22_port_o_2_5;
  assign subBytes_out_6_2_6 = sbox_AES_BoyarPeralta_22_port_o_2_6;
  assign subBytes_out_6_2_7 = sbox_AES_BoyarPeralta_22_port_o_2_7;
  assign subBytes_out_6_3_0 = sbox_AES_BoyarPeralta_22_port_o_3_0;
  assign subBytes_out_6_3_1 = sbox_AES_BoyarPeralta_22_port_o_3_1;
  assign subBytes_out_6_3_2 = sbox_AES_BoyarPeralta_22_port_o_3_2;
  assign subBytes_out_6_3_3 = sbox_AES_BoyarPeralta_22_port_o_3_3;
  assign subBytes_out_6_3_4 = sbox_AES_BoyarPeralta_22_port_o_3_4;
  assign subBytes_out_6_3_5 = sbox_AES_BoyarPeralta_22_port_o_3_5;
  assign subBytes_out_6_3_6 = sbox_AES_BoyarPeralta_22_port_o_3_6;
  assign subBytes_out_6_3_7 = sbox_AES_BoyarPeralta_22_port_o_3_7;
  assign subBytes_out_7_0_0 = sbox_AES_BoyarPeralta_23_port_o_0_0;
  assign subBytes_out_7_0_1 = sbox_AES_BoyarPeralta_23_port_o_0_1;
  assign subBytes_out_7_0_2 = sbox_AES_BoyarPeralta_23_port_o_0_2;
  assign subBytes_out_7_0_3 = sbox_AES_BoyarPeralta_23_port_o_0_3;
  assign subBytes_out_7_0_4 = sbox_AES_BoyarPeralta_23_port_o_0_4;
  assign subBytes_out_7_0_5 = sbox_AES_BoyarPeralta_23_port_o_0_5;
  assign subBytes_out_7_0_6 = sbox_AES_BoyarPeralta_23_port_o_0_6;
  assign subBytes_out_7_0_7 = sbox_AES_BoyarPeralta_23_port_o_0_7;
  assign subBytes_out_7_1_0 = sbox_AES_BoyarPeralta_23_port_o_1_0;
  assign subBytes_out_7_1_1 = sbox_AES_BoyarPeralta_23_port_o_1_1;
  assign subBytes_out_7_1_2 = sbox_AES_BoyarPeralta_23_port_o_1_2;
  assign subBytes_out_7_1_3 = sbox_AES_BoyarPeralta_23_port_o_1_3;
  assign subBytes_out_7_1_4 = sbox_AES_BoyarPeralta_23_port_o_1_4;
  assign subBytes_out_7_1_5 = sbox_AES_BoyarPeralta_23_port_o_1_5;
  assign subBytes_out_7_1_6 = sbox_AES_BoyarPeralta_23_port_o_1_6;
  assign subBytes_out_7_1_7 = sbox_AES_BoyarPeralta_23_port_o_1_7;
  assign subBytes_out_7_2_0 = sbox_AES_BoyarPeralta_23_port_o_2_0;
  assign subBytes_out_7_2_1 = sbox_AES_BoyarPeralta_23_port_o_2_1;
  assign subBytes_out_7_2_2 = sbox_AES_BoyarPeralta_23_port_o_2_2;
  assign subBytes_out_7_2_3 = sbox_AES_BoyarPeralta_23_port_o_2_3;
  assign subBytes_out_7_2_4 = sbox_AES_BoyarPeralta_23_port_o_2_4;
  assign subBytes_out_7_2_5 = sbox_AES_BoyarPeralta_23_port_o_2_5;
  assign subBytes_out_7_2_6 = sbox_AES_BoyarPeralta_23_port_o_2_6;
  assign subBytes_out_7_2_7 = sbox_AES_BoyarPeralta_23_port_o_2_7;
  assign subBytes_out_7_3_0 = sbox_AES_BoyarPeralta_23_port_o_3_0;
  assign subBytes_out_7_3_1 = sbox_AES_BoyarPeralta_23_port_o_3_1;
  assign subBytes_out_7_3_2 = sbox_AES_BoyarPeralta_23_port_o_3_2;
  assign subBytes_out_7_3_3 = sbox_AES_BoyarPeralta_23_port_o_3_3;
  assign subBytes_out_7_3_4 = sbox_AES_BoyarPeralta_23_port_o_3_4;
  assign subBytes_out_7_3_5 = sbox_AES_BoyarPeralta_23_port_o_3_5;
  assign subBytes_out_7_3_6 = sbox_AES_BoyarPeralta_23_port_o_3_6;
  assign subBytes_out_7_3_7 = sbox_AES_BoyarPeralta_23_port_o_3_7;
  assign subBytes_out_8_0_0 = sbox_AES_BoyarPeralta_24_port_o_0_0;
  assign subBytes_out_8_0_1 = sbox_AES_BoyarPeralta_24_port_o_0_1;
  assign subBytes_out_8_0_2 = sbox_AES_BoyarPeralta_24_port_o_0_2;
  assign subBytes_out_8_0_3 = sbox_AES_BoyarPeralta_24_port_o_0_3;
  assign subBytes_out_8_0_4 = sbox_AES_BoyarPeralta_24_port_o_0_4;
  assign subBytes_out_8_0_5 = sbox_AES_BoyarPeralta_24_port_o_0_5;
  assign subBytes_out_8_0_6 = sbox_AES_BoyarPeralta_24_port_o_0_6;
  assign subBytes_out_8_0_7 = sbox_AES_BoyarPeralta_24_port_o_0_7;
  assign subBytes_out_8_1_0 = sbox_AES_BoyarPeralta_24_port_o_1_0;
  assign subBytes_out_8_1_1 = sbox_AES_BoyarPeralta_24_port_o_1_1;
  assign subBytes_out_8_1_2 = sbox_AES_BoyarPeralta_24_port_o_1_2;
  assign subBytes_out_8_1_3 = sbox_AES_BoyarPeralta_24_port_o_1_3;
  assign subBytes_out_8_1_4 = sbox_AES_BoyarPeralta_24_port_o_1_4;
  assign subBytes_out_8_1_5 = sbox_AES_BoyarPeralta_24_port_o_1_5;
  assign subBytes_out_8_1_6 = sbox_AES_BoyarPeralta_24_port_o_1_6;
  assign subBytes_out_8_1_7 = sbox_AES_BoyarPeralta_24_port_o_1_7;
  assign subBytes_out_8_2_0 = sbox_AES_BoyarPeralta_24_port_o_2_0;
  assign subBytes_out_8_2_1 = sbox_AES_BoyarPeralta_24_port_o_2_1;
  assign subBytes_out_8_2_2 = sbox_AES_BoyarPeralta_24_port_o_2_2;
  assign subBytes_out_8_2_3 = sbox_AES_BoyarPeralta_24_port_o_2_3;
  assign subBytes_out_8_2_4 = sbox_AES_BoyarPeralta_24_port_o_2_4;
  assign subBytes_out_8_2_5 = sbox_AES_BoyarPeralta_24_port_o_2_5;
  assign subBytes_out_8_2_6 = sbox_AES_BoyarPeralta_24_port_o_2_6;
  assign subBytes_out_8_2_7 = sbox_AES_BoyarPeralta_24_port_o_2_7;
  assign subBytes_out_8_3_0 = sbox_AES_BoyarPeralta_24_port_o_3_0;
  assign subBytes_out_8_3_1 = sbox_AES_BoyarPeralta_24_port_o_3_1;
  assign subBytes_out_8_3_2 = sbox_AES_BoyarPeralta_24_port_o_3_2;
  assign subBytes_out_8_3_3 = sbox_AES_BoyarPeralta_24_port_o_3_3;
  assign subBytes_out_8_3_4 = sbox_AES_BoyarPeralta_24_port_o_3_4;
  assign subBytes_out_8_3_5 = sbox_AES_BoyarPeralta_24_port_o_3_5;
  assign subBytes_out_8_3_6 = sbox_AES_BoyarPeralta_24_port_o_3_6;
  assign subBytes_out_8_3_7 = sbox_AES_BoyarPeralta_24_port_o_3_7;
  assign subBytes_out_9_0_0 = sbox_AES_BoyarPeralta_25_port_o_0_0;
  assign subBytes_out_9_0_1 = sbox_AES_BoyarPeralta_25_port_o_0_1;
  assign subBytes_out_9_0_2 = sbox_AES_BoyarPeralta_25_port_o_0_2;
  assign subBytes_out_9_0_3 = sbox_AES_BoyarPeralta_25_port_o_0_3;
  assign subBytes_out_9_0_4 = sbox_AES_BoyarPeralta_25_port_o_0_4;
  assign subBytes_out_9_0_5 = sbox_AES_BoyarPeralta_25_port_o_0_5;
  assign subBytes_out_9_0_6 = sbox_AES_BoyarPeralta_25_port_o_0_6;
  assign subBytes_out_9_0_7 = sbox_AES_BoyarPeralta_25_port_o_0_7;
  assign subBytes_out_9_1_0 = sbox_AES_BoyarPeralta_25_port_o_1_0;
  assign subBytes_out_9_1_1 = sbox_AES_BoyarPeralta_25_port_o_1_1;
  assign subBytes_out_9_1_2 = sbox_AES_BoyarPeralta_25_port_o_1_2;
  assign subBytes_out_9_1_3 = sbox_AES_BoyarPeralta_25_port_o_1_3;
  assign subBytes_out_9_1_4 = sbox_AES_BoyarPeralta_25_port_o_1_4;
  assign subBytes_out_9_1_5 = sbox_AES_BoyarPeralta_25_port_o_1_5;
  assign subBytes_out_9_1_6 = sbox_AES_BoyarPeralta_25_port_o_1_6;
  assign subBytes_out_9_1_7 = sbox_AES_BoyarPeralta_25_port_o_1_7;
  assign subBytes_out_9_2_0 = sbox_AES_BoyarPeralta_25_port_o_2_0;
  assign subBytes_out_9_2_1 = sbox_AES_BoyarPeralta_25_port_o_2_1;
  assign subBytes_out_9_2_2 = sbox_AES_BoyarPeralta_25_port_o_2_2;
  assign subBytes_out_9_2_3 = sbox_AES_BoyarPeralta_25_port_o_2_3;
  assign subBytes_out_9_2_4 = sbox_AES_BoyarPeralta_25_port_o_2_4;
  assign subBytes_out_9_2_5 = sbox_AES_BoyarPeralta_25_port_o_2_5;
  assign subBytes_out_9_2_6 = sbox_AES_BoyarPeralta_25_port_o_2_6;
  assign subBytes_out_9_2_7 = sbox_AES_BoyarPeralta_25_port_o_2_7;
  assign subBytes_out_9_3_0 = sbox_AES_BoyarPeralta_25_port_o_3_0;
  assign subBytes_out_9_3_1 = sbox_AES_BoyarPeralta_25_port_o_3_1;
  assign subBytes_out_9_3_2 = sbox_AES_BoyarPeralta_25_port_o_3_2;
  assign subBytes_out_9_3_3 = sbox_AES_BoyarPeralta_25_port_o_3_3;
  assign subBytes_out_9_3_4 = sbox_AES_BoyarPeralta_25_port_o_3_4;
  assign subBytes_out_9_3_5 = sbox_AES_BoyarPeralta_25_port_o_3_5;
  assign subBytes_out_9_3_6 = sbox_AES_BoyarPeralta_25_port_o_3_6;
  assign subBytes_out_9_3_7 = sbox_AES_BoyarPeralta_25_port_o_3_7;
  assign subBytes_out_10_0_0 = sbox_AES_BoyarPeralta_26_port_o_0_0;
  assign subBytes_out_10_0_1 = sbox_AES_BoyarPeralta_26_port_o_0_1;
  assign subBytes_out_10_0_2 = sbox_AES_BoyarPeralta_26_port_o_0_2;
  assign subBytes_out_10_0_3 = sbox_AES_BoyarPeralta_26_port_o_0_3;
  assign subBytes_out_10_0_4 = sbox_AES_BoyarPeralta_26_port_o_0_4;
  assign subBytes_out_10_0_5 = sbox_AES_BoyarPeralta_26_port_o_0_5;
  assign subBytes_out_10_0_6 = sbox_AES_BoyarPeralta_26_port_o_0_6;
  assign subBytes_out_10_0_7 = sbox_AES_BoyarPeralta_26_port_o_0_7;
  assign subBytes_out_10_1_0 = sbox_AES_BoyarPeralta_26_port_o_1_0;
  assign subBytes_out_10_1_1 = sbox_AES_BoyarPeralta_26_port_o_1_1;
  assign subBytes_out_10_1_2 = sbox_AES_BoyarPeralta_26_port_o_1_2;
  assign subBytes_out_10_1_3 = sbox_AES_BoyarPeralta_26_port_o_1_3;
  assign subBytes_out_10_1_4 = sbox_AES_BoyarPeralta_26_port_o_1_4;
  assign subBytes_out_10_1_5 = sbox_AES_BoyarPeralta_26_port_o_1_5;
  assign subBytes_out_10_1_6 = sbox_AES_BoyarPeralta_26_port_o_1_6;
  assign subBytes_out_10_1_7 = sbox_AES_BoyarPeralta_26_port_o_1_7;
  assign subBytes_out_10_2_0 = sbox_AES_BoyarPeralta_26_port_o_2_0;
  assign subBytes_out_10_2_1 = sbox_AES_BoyarPeralta_26_port_o_2_1;
  assign subBytes_out_10_2_2 = sbox_AES_BoyarPeralta_26_port_o_2_2;
  assign subBytes_out_10_2_3 = sbox_AES_BoyarPeralta_26_port_o_2_3;
  assign subBytes_out_10_2_4 = sbox_AES_BoyarPeralta_26_port_o_2_4;
  assign subBytes_out_10_2_5 = sbox_AES_BoyarPeralta_26_port_o_2_5;
  assign subBytes_out_10_2_6 = sbox_AES_BoyarPeralta_26_port_o_2_6;
  assign subBytes_out_10_2_7 = sbox_AES_BoyarPeralta_26_port_o_2_7;
  assign subBytes_out_10_3_0 = sbox_AES_BoyarPeralta_26_port_o_3_0;
  assign subBytes_out_10_3_1 = sbox_AES_BoyarPeralta_26_port_o_3_1;
  assign subBytes_out_10_3_2 = sbox_AES_BoyarPeralta_26_port_o_3_2;
  assign subBytes_out_10_3_3 = sbox_AES_BoyarPeralta_26_port_o_3_3;
  assign subBytes_out_10_3_4 = sbox_AES_BoyarPeralta_26_port_o_3_4;
  assign subBytes_out_10_3_5 = sbox_AES_BoyarPeralta_26_port_o_3_5;
  assign subBytes_out_10_3_6 = sbox_AES_BoyarPeralta_26_port_o_3_6;
  assign subBytes_out_10_3_7 = sbox_AES_BoyarPeralta_26_port_o_3_7;
  assign subBytes_out_11_0_0 = sbox_AES_BoyarPeralta_27_port_o_0_0;
  assign subBytes_out_11_0_1 = sbox_AES_BoyarPeralta_27_port_o_0_1;
  assign subBytes_out_11_0_2 = sbox_AES_BoyarPeralta_27_port_o_0_2;
  assign subBytes_out_11_0_3 = sbox_AES_BoyarPeralta_27_port_o_0_3;
  assign subBytes_out_11_0_4 = sbox_AES_BoyarPeralta_27_port_o_0_4;
  assign subBytes_out_11_0_5 = sbox_AES_BoyarPeralta_27_port_o_0_5;
  assign subBytes_out_11_0_6 = sbox_AES_BoyarPeralta_27_port_o_0_6;
  assign subBytes_out_11_0_7 = sbox_AES_BoyarPeralta_27_port_o_0_7;
  assign subBytes_out_11_1_0 = sbox_AES_BoyarPeralta_27_port_o_1_0;
  assign subBytes_out_11_1_1 = sbox_AES_BoyarPeralta_27_port_o_1_1;
  assign subBytes_out_11_1_2 = sbox_AES_BoyarPeralta_27_port_o_1_2;
  assign subBytes_out_11_1_3 = sbox_AES_BoyarPeralta_27_port_o_1_3;
  assign subBytes_out_11_1_4 = sbox_AES_BoyarPeralta_27_port_o_1_4;
  assign subBytes_out_11_1_5 = sbox_AES_BoyarPeralta_27_port_o_1_5;
  assign subBytes_out_11_1_6 = sbox_AES_BoyarPeralta_27_port_o_1_6;
  assign subBytes_out_11_1_7 = sbox_AES_BoyarPeralta_27_port_o_1_7;
  assign subBytes_out_11_2_0 = sbox_AES_BoyarPeralta_27_port_o_2_0;
  assign subBytes_out_11_2_1 = sbox_AES_BoyarPeralta_27_port_o_2_1;
  assign subBytes_out_11_2_2 = sbox_AES_BoyarPeralta_27_port_o_2_2;
  assign subBytes_out_11_2_3 = sbox_AES_BoyarPeralta_27_port_o_2_3;
  assign subBytes_out_11_2_4 = sbox_AES_BoyarPeralta_27_port_o_2_4;
  assign subBytes_out_11_2_5 = sbox_AES_BoyarPeralta_27_port_o_2_5;
  assign subBytes_out_11_2_6 = sbox_AES_BoyarPeralta_27_port_o_2_6;
  assign subBytes_out_11_2_7 = sbox_AES_BoyarPeralta_27_port_o_2_7;
  assign subBytes_out_11_3_0 = sbox_AES_BoyarPeralta_27_port_o_3_0;
  assign subBytes_out_11_3_1 = sbox_AES_BoyarPeralta_27_port_o_3_1;
  assign subBytes_out_11_3_2 = sbox_AES_BoyarPeralta_27_port_o_3_2;
  assign subBytes_out_11_3_3 = sbox_AES_BoyarPeralta_27_port_o_3_3;
  assign subBytes_out_11_3_4 = sbox_AES_BoyarPeralta_27_port_o_3_4;
  assign subBytes_out_11_3_5 = sbox_AES_BoyarPeralta_27_port_o_3_5;
  assign subBytes_out_11_3_6 = sbox_AES_BoyarPeralta_27_port_o_3_6;
  assign subBytes_out_11_3_7 = sbox_AES_BoyarPeralta_27_port_o_3_7;
  assign subBytes_out_12_0_0 = sbox_AES_BoyarPeralta_28_port_o_0_0;
  assign subBytes_out_12_0_1 = sbox_AES_BoyarPeralta_28_port_o_0_1;
  assign subBytes_out_12_0_2 = sbox_AES_BoyarPeralta_28_port_o_0_2;
  assign subBytes_out_12_0_3 = sbox_AES_BoyarPeralta_28_port_o_0_3;
  assign subBytes_out_12_0_4 = sbox_AES_BoyarPeralta_28_port_o_0_4;
  assign subBytes_out_12_0_5 = sbox_AES_BoyarPeralta_28_port_o_0_5;
  assign subBytes_out_12_0_6 = sbox_AES_BoyarPeralta_28_port_o_0_6;
  assign subBytes_out_12_0_7 = sbox_AES_BoyarPeralta_28_port_o_0_7;
  assign subBytes_out_12_1_0 = sbox_AES_BoyarPeralta_28_port_o_1_0;
  assign subBytes_out_12_1_1 = sbox_AES_BoyarPeralta_28_port_o_1_1;
  assign subBytes_out_12_1_2 = sbox_AES_BoyarPeralta_28_port_o_1_2;
  assign subBytes_out_12_1_3 = sbox_AES_BoyarPeralta_28_port_o_1_3;
  assign subBytes_out_12_1_4 = sbox_AES_BoyarPeralta_28_port_o_1_4;
  assign subBytes_out_12_1_5 = sbox_AES_BoyarPeralta_28_port_o_1_5;
  assign subBytes_out_12_1_6 = sbox_AES_BoyarPeralta_28_port_o_1_6;
  assign subBytes_out_12_1_7 = sbox_AES_BoyarPeralta_28_port_o_1_7;
  assign subBytes_out_12_2_0 = sbox_AES_BoyarPeralta_28_port_o_2_0;
  assign subBytes_out_12_2_1 = sbox_AES_BoyarPeralta_28_port_o_2_1;
  assign subBytes_out_12_2_2 = sbox_AES_BoyarPeralta_28_port_o_2_2;
  assign subBytes_out_12_2_3 = sbox_AES_BoyarPeralta_28_port_o_2_3;
  assign subBytes_out_12_2_4 = sbox_AES_BoyarPeralta_28_port_o_2_4;
  assign subBytes_out_12_2_5 = sbox_AES_BoyarPeralta_28_port_o_2_5;
  assign subBytes_out_12_2_6 = sbox_AES_BoyarPeralta_28_port_o_2_6;
  assign subBytes_out_12_2_7 = sbox_AES_BoyarPeralta_28_port_o_2_7;
  assign subBytes_out_12_3_0 = sbox_AES_BoyarPeralta_28_port_o_3_0;
  assign subBytes_out_12_3_1 = sbox_AES_BoyarPeralta_28_port_o_3_1;
  assign subBytes_out_12_3_2 = sbox_AES_BoyarPeralta_28_port_o_3_2;
  assign subBytes_out_12_3_3 = sbox_AES_BoyarPeralta_28_port_o_3_3;
  assign subBytes_out_12_3_4 = sbox_AES_BoyarPeralta_28_port_o_3_4;
  assign subBytes_out_12_3_5 = sbox_AES_BoyarPeralta_28_port_o_3_5;
  assign subBytes_out_12_3_6 = sbox_AES_BoyarPeralta_28_port_o_3_6;
  assign subBytes_out_12_3_7 = sbox_AES_BoyarPeralta_28_port_o_3_7;
  assign subBytes_out_13_0_0 = sbox_AES_BoyarPeralta_29_port_o_0_0;
  assign subBytes_out_13_0_1 = sbox_AES_BoyarPeralta_29_port_o_0_1;
  assign subBytes_out_13_0_2 = sbox_AES_BoyarPeralta_29_port_o_0_2;
  assign subBytes_out_13_0_3 = sbox_AES_BoyarPeralta_29_port_o_0_3;
  assign subBytes_out_13_0_4 = sbox_AES_BoyarPeralta_29_port_o_0_4;
  assign subBytes_out_13_0_5 = sbox_AES_BoyarPeralta_29_port_o_0_5;
  assign subBytes_out_13_0_6 = sbox_AES_BoyarPeralta_29_port_o_0_6;
  assign subBytes_out_13_0_7 = sbox_AES_BoyarPeralta_29_port_o_0_7;
  assign subBytes_out_13_1_0 = sbox_AES_BoyarPeralta_29_port_o_1_0;
  assign subBytes_out_13_1_1 = sbox_AES_BoyarPeralta_29_port_o_1_1;
  assign subBytes_out_13_1_2 = sbox_AES_BoyarPeralta_29_port_o_1_2;
  assign subBytes_out_13_1_3 = sbox_AES_BoyarPeralta_29_port_o_1_3;
  assign subBytes_out_13_1_4 = sbox_AES_BoyarPeralta_29_port_o_1_4;
  assign subBytes_out_13_1_5 = sbox_AES_BoyarPeralta_29_port_o_1_5;
  assign subBytes_out_13_1_6 = sbox_AES_BoyarPeralta_29_port_o_1_6;
  assign subBytes_out_13_1_7 = sbox_AES_BoyarPeralta_29_port_o_1_7;
  assign subBytes_out_13_2_0 = sbox_AES_BoyarPeralta_29_port_o_2_0;
  assign subBytes_out_13_2_1 = sbox_AES_BoyarPeralta_29_port_o_2_1;
  assign subBytes_out_13_2_2 = sbox_AES_BoyarPeralta_29_port_o_2_2;
  assign subBytes_out_13_2_3 = sbox_AES_BoyarPeralta_29_port_o_2_3;
  assign subBytes_out_13_2_4 = sbox_AES_BoyarPeralta_29_port_o_2_4;
  assign subBytes_out_13_2_5 = sbox_AES_BoyarPeralta_29_port_o_2_5;
  assign subBytes_out_13_2_6 = sbox_AES_BoyarPeralta_29_port_o_2_6;
  assign subBytes_out_13_2_7 = sbox_AES_BoyarPeralta_29_port_o_2_7;
  assign subBytes_out_13_3_0 = sbox_AES_BoyarPeralta_29_port_o_3_0;
  assign subBytes_out_13_3_1 = sbox_AES_BoyarPeralta_29_port_o_3_1;
  assign subBytes_out_13_3_2 = sbox_AES_BoyarPeralta_29_port_o_3_2;
  assign subBytes_out_13_3_3 = sbox_AES_BoyarPeralta_29_port_o_3_3;
  assign subBytes_out_13_3_4 = sbox_AES_BoyarPeralta_29_port_o_3_4;
  assign subBytes_out_13_3_5 = sbox_AES_BoyarPeralta_29_port_o_3_5;
  assign subBytes_out_13_3_6 = sbox_AES_BoyarPeralta_29_port_o_3_6;
  assign subBytes_out_13_3_7 = sbox_AES_BoyarPeralta_29_port_o_3_7;
  assign subBytes_out_14_0_0 = sbox_AES_BoyarPeralta_30_port_o_0_0;
  assign subBytes_out_14_0_1 = sbox_AES_BoyarPeralta_30_port_o_0_1;
  assign subBytes_out_14_0_2 = sbox_AES_BoyarPeralta_30_port_o_0_2;
  assign subBytes_out_14_0_3 = sbox_AES_BoyarPeralta_30_port_o_0_3;
  assign subBytes_out_14_0_4 = sbox_AES_BoyarPeralta_30_port_o_0_4;
  assign subBytes_out_14_0_5 = sbox_AES_BoyarPeralta_30_port_o_0_5;
  assign subBytes_out_14_0_6 = sbox_AES_BoyarPeralta_30_port_o_0_6;
  assign subBytes_out_14_0_7 = sbox_AES_BoyarPeralta_30_port_o_0_7;
  assign subBytes_out_14_1_0 = sbox_AES_BoyarPeralta_30_port_o_1_0;
  assign subBytes_out_14_1_1 = sbox_AES_BoyarPeralta_30_port_o_1_1;
  assign subBytes_out_14_1_2 = sbox_AES_BoyarPeralta_30_port_o_1_2;
  assign subBytes_out_14_1_3 = sbox_AES_BoyarPeralta_30_port_o_1_3;
  assign subBytes_out_14_1_4 = sbox_AES_BoyarPeralta_30_port_o_1_4;
  assign subBytes_out_14_1_5 = sbox_AES_BoyarPeralta_30_port_o_1_5;
  assign subBytes_out_14_1_6 = sbox_AES_BoyarPeralta_30_port_o_1_6;
  assign subBytes_out_14_1_7 = sbox_AES_BoyarPeralta_30_port_o_1_7;
  assign subBytes_out_14_2_0 = sbox_AES_BoyarPeralta_30_port_o_2_0;
  assign subBytes_out_14_2_1 = sbox_AES_BoyarPeralta_30_port_o_2_1;
  assign subBytes_out_14_2_2 = sbox_AES_BoyarPeralta_30_port_o_2_2;
  assign subBytes_out_14_2_3 = sbox_AES_BoyarPeralta_30_port_o_2_3;
  assign subBytes_out_14_2_4 = sbox_AES_BoyarPeralta_30_port_o_2_4;
  assign subBytes_out_14_2_5 = sbox_AES_BoyarPeralta_30_port_o_2_5;
  assign subBytes_out_14_2_6 = sbox_AES_BoyarPeralta_30_port_o_2_6;
  assign subBytes_out_14_2_7 = sbox_AES_BoyarPeralta_30_port_o_2_7;
  assign subBytes_out_14_3_0 = sbox_AES_BoyarPeralta_30_port_o_3_0;
  assign subBytes_out_14_3_1 = sbox_AES_BoyarPeralta_30_port_o_3_1;
  assign subBytes_out_14_3_2 = sbox_AES_BoyarPeralta_30_port_o_3_2;
  assign subBytes_out_14_3_3 = sbox_AES_BoyarPeralta_30_port_o_3_3;
  assign subBytes_out_14_3_4 = sbox_AES_BoyarPeralta_30_port_o_3_4;
  assign subBytes_out_14_3_5 = sbox_AES_BoyarPeralta_30_port_o_3_5;
  assign subBytes_out_14_3_6 = sbox_AES_BoyarPeralta_30_port_o_3_6;
  assign subBytes_out_14_3_7 = sbox_AES_BoyarPeralta_30_port_o_3_7;
  assign subBytes_out_15_0_0 = sbox_AES_BoyarPeralta_31_port_o_0_0;
  assign subBytes_out_15_0_1 = sbox_AES_BoyarPeralta_31_port_o_0_1;
  assign subBytes_out_15_0_2 = sbox_AES_BoyarPeralta_31_port_o_0_2;
  assign subBytes_out_15_0_3 = sbox_AES_BoyarPeralta_31_port_o_0_3;
  assign subBytes_out_15_0_4 = sbox_AES_BoyarPeralta_31_port_o_0_4;
  assign subBytes_out_15_0_5 = sbox_AES_BoyarPeralta_31_port_o_0_5;
  assign subBytes_out_15_0_6 = sbox_AES_BoyarPeralta_31_port_o_0_6;
  assign subBytes_out_15_0_7 = sbox_AES_BoyarPeralta_31_port_o_0_7;
  assign subBytes_out_15_1_0 = sbox_AES_BoyarPeralta_31_port_o_1_0;
  assign subBytes_out_15_1_1 = sbox_AES_BoyarPeralta_31_port_o_1_1;
  assign subBytes_out_15_1_2 = sbox_AES_BoyarPeralta_31_port_o_1_2;
  assign subBytes_out_15_1_3 = sbox_AES_BoyarPeralta_31_port_o_1_3;
  assign subBytes_out_15_1_4 = sbox_AES_BoyarPeralta_31_port_o_1_4;
  assign subBytes_out_15_1_5 = sbox_AES_BoyarPeralta_31_port_o_1_5;
  assign subBytes_out_15_1_6 = sbox_AES_BoyarPeralta_31_port_o_1_6;
  assign subBytes_out_15_1_7 = sbox_AES_BoyarPeralta_31_port_o_1_7;
  assign subBytes_out_15_2_0 = sbox_AES_BoyarPeralta_31_port_o_2_0;
  assign subBytes_out_15_2_1 = sbox_AES_BoyarPeralta_31_port_o_2_1;
  assign subBytes_out_15_2_2 = sbox_AES_BoyarPeralta_31_port_o_2_2;
  assign subBytes_out_15_2_3 = sbox_AES_BoyarPeralta_31_port_o_2_3;
  assign subBytes_out_15_2_4 = sbox_AES_BoyarPeralta_31_port_o_2_4;
  assign subBytes_out_15_2_5 = sbox_AES_BoyarPeralta_31_port_o_2_5;
  assign subBytes_out_15_2_6 = sbox_AES_BoyarPeralta_31_port_o_2_6;
  assign subBytes_out_15_2_7 = sbox_AES_BoyarPeralta_31_port_o_2_7;
  assign subBytes_out_15_3_0 = sbox_AES_BoyarPeralta_31_port_o_3_0;
  assign subBytes_out_15_3_1 = sbox_AES_BoyarPeralta_31_port_o_3_1;
  assign subBytes_out_15_3_2 = sbox_AES_BoyarPeralta_31_port_o_3_2;
  assign subBytes_out_15_3_3 = sbox_AES_BoyarPeralta_31_port_o_3_3;
  assign subBytes_out_15_3_4 = sbox_AES_BoyarPeralta_31_port_o_3_4;
  assign subBytes_out_15_3_5 = sbox_AES_BoyarPeralta_31_port_o_3_5;
  assign subBytes_out_15_3_6 = sbox_AES_BoyarPeralta_31_port_o_3_6;
  assign subBytes_out_15_3_7 = sbox_AES_BoyarPeralta_31_port_o_3_7;
  assign port_state_out_0_0_0 = roundReg_0_0_0;
  assign port_state_out_0_0_1 = roundReg_0_0_1;
  assign port_state_out_0_0_2 = roundReg_0_0_2;
  assign port_state_out_0_0_3 = roundReg_0_0_3;
  assign port_state_out_0_0_4 = roundReg_0_0_4;
  assign port_state_out_0_0_5 = roundReg_0_0_5;
  assign port_state_out_0_0_6 = roundReg_0_0_6;
  assign port_state_out_0_0_7 = roundReg_0_0_7;
  assign port_state_out_0_1_0 = roundReg_0_1_0;
  assign port_state_out_0_1_1 = roundReg_0_1_1;
  assign port_state_out_0_1_2 = roundReg_0_1_2;
  assign port_state_out_0_1_3 = roundReg_0_1_3;
  assign port_state_out_0_1_4 = roundReg_0_1_4;
  assign port_state_out_0_1_5 = roundReg_0_1_5;
  assign port_state_out_0_1_6 = roundReg_0_1_6;
  assign port_state_out_0_1_7 = roundReg_0_1_7;
  assign port_state_out_0_2_0 = roundReg_0_2_0;
  assign port_state_out_0_2_1 = roundReg_0_2_1;
  assign port_state_out_0_2_2 = roundReg_0_2_2;
  assign port_state_out_0_2_3 = roundReg_0_2_3;
  assign port_state_out_0_2_4 = roundReg_0_2_4;
  assign port_state_out_0_2_5 = roundReg_0_2_5;
  assign port_state_out_0_2_6 = roundReg_0_2_6;
  assign port_state_out_0_2_7 = roundReg_0_2_7;
  assign port_state_out_0_3_0 = roundReg_0_3_0;
  assign port_state_out_0_3_1 = roundReg_0_3_1;
  assign port_state_out_0_3_2 = roundReg_0_3_2;
  assign port_state_out_0_3_3 = roundReg_0_3_3;
  assign port_state_out_0_3_4 = roundReg_0_3_4;
  assign port_state_out_0_3_5 = roundReg_0_3_5;
  assign port_state_out_0_3_6 = roundReg_0_3_6;
  assign port_state_out_0_3_7 = roundReg_0_3_7;
  assign port_state_out_1_0_0 = roundReg_1_0_0;
  assign port_state_out_1_0_1 = roundReg_1_0_1;
  assign port_state_out_1_0_2 = roundReg_1_0_2;
  assign port_state_out_1_0_3 = roundReg_1_0_3;
  assign port_state_out_1_0_4 = roundReg_1_0_4;
  assign port_state_out_1_0_5 = roundReg_1_0_5;
  assign port_state_out_1_0_6 = roundReg_1_0_6;
  assign port_state_out_1_0_7 = roundReg_1_0_7;
  assign port_state_out_1_1_0 = roundReg_1_1_0;
  assign port_state_out_1_1_1 = roundReg_1_1_1;
  assign port_state_out_1_1_2 = roundReg_1_1_2;
  assign port_state_out_1_1_3 = roundReg_1_1_3;
  assign port_state_out_1_1_4 = roundReg_1_1_4;
  assign port_state_out_1_1_5 = roundReg_1_1_5;
  assign port_state_out_1_1_6 = roundReg_1_1_6;
  assign port_state_out_1_1_7 = roundReg_1_1_7;
  assign port_state_out_1_2_0 = roundReg_1_2_0;
  assign port_state_out_1_2_1 = roundReg_1_2_1;
  assign port_state_out_1_2_2 = roundReg_1_2_2;
  assign port_state_out_1_2_3 = roundReg_1_2_3;
  assign port_state_out_1_2_4 = roundReg_1_2_4;
  assign port_state_out_1_2_5 = roundReg_1_2_5;
  assign port_state_out_1_2_6 = roundReg_1_2_6;
  assign port_state_out_1_2_7 = roundReg_1_2_7;
  assign port_state_out_1_3_0 = roundReg_1_3_0;
  assign port_state_out_1_3_1 = roundReg_1_3_1;
  assign port_state_out_1_3_2 = roundReg_1_3_2;
  assign port_state_out_1_3_3 = roundReg_1_3_3;
  assign port_state_out_1_3_4 = roundReg_1_3_4;
  assign port_state_out_1_3_5 = roundReg_1_3_5;
  assign port_state_out_1_3_6 = roundReg_1_3_6;
  assign port_state_out_1_3_7 = roundReg_1_3_7;
  assign port_state_out_2_0_0 = roundReg_2_0_0;
  assign port_state_out_2_0_1 = roundReg_2_0_1;
  assign port_state_out_2_0_2 = roundReg_2_0_2;
  assign port_state_out_2_0_3 = roundReg_2_0_3;
  assign port_state_out_2_0_4 = roundReg_2_0_4;
  assign port_state_out_2_0_5 = roundReg_2_0_5;
  assign port_state_out_2_0_6 = roundReg_2_0_6;
  assign port_state_out_2_0_7 = roundReg_2_0_7;
  assign port_state_out_2_1_0 = roundReg_2_1_0;
  assign port_state_out_2_1_1 = roundReg_2_1_1;
  assign port_state_out_2_1_2 = roundReg_2_1_2;
  assign port_state_out_2_1_3 = roundReg_2_1_3;
  assign port_state_out_2_1_4 = roundReg_2_1_4;
  assign port_state_out_2_1_5 = roundReg_2_1_5;
  assign port_state_out_2_1_6 = roundReg_2_1_6;
  assign port_state_out_2_1_7 = roundReg_2_1_7;
  assign port_state_out_2_2_0 = roundReg_2_2_0;
  assign port_state_out_2_2_1 = roundReg_2_2_1;
  assign port_state_out_2_2_2 = roundReg_2_2_2;
  assign port_state_out_2_2_3 = roundReg_2_2_3;
  assign port_state_out_2_2_4 = roundReg_2_2_4;
  assign port_state_out_2_2_5 = roundReg_2_2_5;
  assign port_state_out_2_2_6 = roundReg_2_2_6;
  assign port_state_out_2_2_7 = roundReg_2_2_7;
  assign port_state_out_2_3_0 = roundReg_2_3_0;
  assign port_state_out_2_3_1 = roundReg_2_3_1;
  assign port_state_out_2_3_2 = roundReg_2_3_2;
  assign port_state_out_2_3_3 = roundReg_2_3_3;
  assign port_state_out_2_3_4 = roundReg_2_3_4;
  assign port_state_out_2_3_5 = roundReg_2_3_5;
  assign port_state_out_2_3_6 = roundReg_2_3_6;
  assign port_state_out_2_3_7 = roundReg_2_3_7;
  assign port_state_out_3_0_0 = roundReg_3_0_0;
  assign port_state_out_3_0_1 = roundReg_3_0_1;
  assign port_state_out_3_0_2 = roundReg_3_0_2;
  assign port_state_out_3_0_3 = roundReg_3_0_3;
  assign port_state_out_3_0_4 = roundReg_3_0_4;
  assign port_state_out_3_0_5 = roundReg_3_0_5;
  assign port_state_out_3_0_6 = roundReg_3_0_6;
  assign port_state_out_3_0_7 = roundReg_3_0_7;
  assign port_state_out_3_1_0 = roundReg_3_1_0;
  assign port_state_out_3_1_1 = roundReg_3_1_1;
  assign port_state_out_3_1_2 = roundReg_3_1_2;
  assign port_state_out_3_1_3 = roundReg_3_1_3;
  assign port_state_out_3_1_4 = roundReg_3_1_4;
  assign port_state_out_3_1_5 = roundReg_3_1_5;
  assign port_state_out_3_1_6 = roundReg_3_1_6;
  assign port_state_out_3_1_7 = roundReg_3_1_7;
  assign port_state_out_3_2_0 = roundReg_3_2_0;
  assign port_state_out_3_2_1 = roundReg_3_2_1;
  assign port_state_out_3_2_2 = roundReg_3_2_2;
  assign port_state_out_3_2_3 = roundReg_3_2_3;
  assign port_state_out_3_2_4 = roundReg_3_2_4;
  assign port_state_out_3_2_5 = roundReg_3_2_5;
  assign port_state_out_3_2_6 = roundReg_3_2_6;
  assign port_state_out_3_2_7 = roundReg_3_2_7;
  assign port_state_out_3_3_0 = roundReg_3_3_0;
  assign port_state_out_3_3_1 = roundReg_3_3_1;
  assign port_state_out_3_3_2 = roundReg_3_3_2;
  assign port_state_out_3_3_3 = roundReg_3_3_3;
  assign port_state_out_3_3_4 = roundReg_3_3_4;
  assign port_state_out_3_3_5 = roundReg_3_3_5;
  assign port_state_out_3_3_6 = roundReg_3_3_6;
  assign port_state_out_3_3_7 = roundReg_3_3_7;
  assign port_state_out_4_0_0 = roundReg_4_0_0;
  assign port_state_out_4_0_1 = roundReg_4_0_1;
  assign port_state_out_4_0_2 = roundReg_4_0_2;
  assign port_state_out_4_0_3 = roundReg_4_0_3;
  assign port_state_out_4_0_4 = roundReg_4_0_4;
  assign port_state_out_4_0_5 = roundReg_4_0_5;
  assign port_state_out_4_0_6 = roundReg_4_0_6;
  assign port_state_out_4_0_7 = roundReg_4_0_7;
  assign port_state_out_4_1_0 = roundReg_4_1_0;
  assign port_state_out_4_1_1 = roundReg_4_1_1;
  assign port_state_out_4_1_2 = roundReg_4_1_2;
  assign port_state_out_4_1_3 = roundReg_4_1_3;
  assign port_state_out_4_1_4 = roundReg_4_1_4;
  assign port_state_out_4_1_5 = roundReg_4_1_5;
  assign port_state_out_4_1_6 = roundReg_4_1_6;
  assign port_state_out_4_1_7 = roundReg_4_1_7;
  assign port_state_out_4_2_0 = roundReg_4_2_0;
  assign port_state_out_4_2_1 = roundReg_4_2_1;
  assign port_state_out_4_2_2 = roundReg_4_2_2;
  assign port_state_out_4_2_3 = roundReg_4_2_3;
  assign port_state_out_4_2_4 = roundReg_4_2_4;
  assign port_state_out_4_2_5 = roundReg_4_2_5;
  assign port_state_out_4_2_6 = roundReg_4_2_6;
  assign port_state_out_4_2_7 = roundReg_4_2_7;
  assign port_state_out_4_3_0 = roundReg_4_3_0;
  assign port_state_out_4_3_1 = roundReg_4_3_1;
  assign port_state_out_4_3_2 = roundReg_4_3_2;
  assign port_state_out_4_3_3 = roundReg_4_3_3;
  assign port_state_out_4_3_4 = roundReg_4_3_4;
  assign port_state_out_4_3_5 = roundReg_4_3_5;
  assign port_state_out_4_3_6 = roundReg_4_3_6;
  assign port_state_out_4_3_7 = roundReg_4_3_7;
  assign port_state_out_5_0_0 = roundReg_5_0_0;
  assign port_state_out_5_0_1 = roundReg_5_0_1;
  assign port_state_out_5_0_2 = roundReg_5_0_2;
  assign port_state_out_5_0_3 = roundReg_5_0_3;
  assign port_state_out_5_0_4 = roundReg_5_0_4;
  assign port_state_out_5_0_5 = roundReg_5_0_5;
  assign port_state_out_5_0_6 = roundReg_5_0_6;
  assign port_state_out_5_0_7 = roundReg_5_0_7;
  assign port_state_out_5_1_0 = roundReg_5_1_0;
  assign port_state_out_5_1_1 = roundReg_5_1_1;
  assign port_state_out_5_1_2 = roundReg_5_1_2;
  assign port_state_out_5_1_3 = roundReg_5_1_3;
  assign port_state_out_5_1_4 = roundReg_5_1_4;
  assign port_state_out_5_1_5 = roundReg_5_1_5;
  assign port_state_out_5_1_6 = roundReg_5_1_6;
  assign port_state_out_5_1_7 = roundReg_5_1_7;
  assign port_state_out_5_2_0 = roundReg_5_2_0;
  assign port_state_out_5_2_1 = roundReg_5_2_1;
  assign port_state_out_5_2_2 = roundReg_5_2_2;
  assign port_state_out_5_2_3 = roundReg_5_2_3;
  assign port_state_out_5_2_4 = roundReg_5_2_4;
  assign port_state_out_5_2_5 = roundReg_5_2_5;
  assign port_state_out_5_2_6 = roundReg_5_2_6;
  assign port_state_out_5_2_7 = roundReg_5_2_7;
  assign port_state_out_5_3_0 = roundReg_5_3_0;
  assign port_state_out_5_3_1 = roundReg_5_3_1;
  assign port_state_out_5_3_2 = roundReg_5_3_2;
  assign port_state_out_5_3_3 = roundReg_5_3_3;
  assign port_state_out_5_3_4 = roundReg_5_3_4;
  assign port_state_out_5_3_5 = roundReg_5_3_5;
  assign port_state_out_5_3_6 = roundReg_5_3_6;
  assign port_state_out_5_3_7 = roundReg_5_3_7;
  assign port_state_out_6_0_0 = roundReg_6_0_0;
  assign port_state_out_6_0_1 = roundReg_6_0_1;
  assign port_state_out_6_0_2 = roundReg_6_0_2;
  assign port_state_out_6_0_3 = roundReg_6_0_3;
  assign port_state_out_6_0_4 = roundReg_6_0_4;
  assign port_state_out_6_0_5 = roundReg_6_0_5;
  assign port_state_out_6_0_6 = roundReg_6_0_6;
  assign port_state_out_6_0_7 = roundReg_6_0_7;
  assign port_state_out_6_1_0 = roundReg_6_1_0;
  assign port_state_out_6_1_1 = roundReg_6_1_1;
  assign port_state_out_6_1_2 = roundReg_6_1_2;
  assign port_state_out_6_1_3 = roundReg_6_1_3;
  assign port_state_out_6_1_4 = roundReg_6_1_4;
  assign port_state_out_6_1_5 = roundReg_6_1_5;
  assign port_state_out_6_1_6 = roundReg_6_1_6;
  assign port_state_out_6_1_7 = roundReg_6_1_7;
  assign port_state_out_6_2_0 = roundReg_6_2_0;
  assign port_state_out_6_2_1 = roundReg_6_2_1;
  assign port_state_out_6_2_2 = roundReg_6_2_2;
  assign port_state_out_6_2_3 = roundReg_6_2_3;
  assign port_state_out_6_2_4 = roundReg_6_2_4;
  assign port_state_out_6_2_5 = roundReg_6_2_5;
  assign port_state_out_6_2_6 = roundReg_6_2_6;
  assign port_state_out_6_2_7 = roundReg_6_2_7;
  assign port_state_out_6_3_0 = roundReg_6_3_0;
  assign port_state_out_6_3_1 = roundReg_6_3_1;
  assign port_state_out_6_3_2 = roundReg_6_3_2;
  assign port_state_out_6_3_3 = roundReg_6_3_3;
  assign port_state_out_6_3_4 = roundReg_6_3_4;
  assign port_state_out_6_3_5 = roundReg_6_3_5;
  assign port_state_out_6_3_6 = roundReg_6_3_6;
  assign port_state_out_6_3_7 = roundReg_6_3_7;
  assign port_state_out_7_0_0 = roundReg_7_0_0;
  assign port_state_out_7_0_1 = roundReg_7_0_1;
  assign port_state_out_7_0_2 = roundReg_7_0_2;
  assign port_state_out_7_0_3 = roundReg_7_0_3;
  assign port_state_out_7_0_4 = roundReg_7_0_4;
  assign port_state_out_7_0_5 = roundReg_7_0_5;
  assign port_state_out_7_0_6 = roundReg_7_0_6;
  assign port_state_out_7_0_7 = roundReg_7_0_7;
  assign port_state_out_7_1_0 = roundReg_7_1_0;
  assign port_state_out_7_1_1 = roundReg_7_1_1;
  assign port_state_out_7_1_2 = roundReg_7_1_2;
  assign port_state_out_7_1_3 = roundReg_7_1_3;
  assign port_state_out_7_1_4 = roundReg_7_1_4;
  assign port_state_out_7_1_5 = roundReg_7_1_5;
  assign port_state_out_7_1_6 = roundReg_7_1_6;
  assign port_state_out_7_1_7 = roundReg_7_1_7;
  assign port_state_out_7_2_0 = roundReg_7_2_0;
  assign port_state_out_7_2_1 = roundReg_7_2_1;
  assign port_state_out_7_2_2 = roundReg_7_2_2;
  assign port_state_out_7_2_3 = roundReg_7_2_3;
  assign port_state_out_7_2_4 = roundReg_7_2_4;
  assign port_state_out_7_2_5 = roundReg_7_2_5;
  assign port_state_out_7_2_6 = roundReg_7_2_6;
  assign port_state_out_7_2_7 = roundReg_7_2_7;
  assign port_state_out_7_3_0 = roundReg_7_3_0;
  assign port_state_out_7_3_1 = roundReg_7_3_1;
  assign port_state_out_7_3_2 = roundReg_7_3_2;
  assign port_state_out_7_3_3 = roundReg_7_3_3;
  assign port_state_out_7_3_4 = roundReg_7_3_4;
  assign port_state_out_7_3_5 = roundReg_7_3_5;
  assign port_state_out_7_3_6 = roundReg_7_3_6;
  assign port_state_out_7_3_7 = roundReg_7_3_7;
  assign port_state_out_8_0_0 = roundReg_8_0_0;
  assign port_state_out_8_0_1 = roundReg_8_0_1;
  assign port_state_out_8_0_2 = roundReg_8_0_2;
  assign port_state_out_8_0_3 = roundReg_8_0_3;
  assign port_state_out_8_0_4 = roundReg_8_0_4;
  assign port_state_out_8_0_5 = roundReg_8_0_5;
  assign port_state_out_8_0_6 = roundReg_8_0_6;
  assign port_state_out_8_0_7 = roundReg_8_0_7;
  assign port_state_out_8_1_0 = roundReg_8_1_0;
  assign port_state_out_8_1_1 = roundReg_8_1_1;
  assign port_state_out_8_1_2 = roundReg_8_1_2;
  assign port_state_out_8_1_3 = roundReg_8_1_3;
  assign port_state_out_8_1_4 = roundReg_8_1_4;
  assign port_state_out_8_1_5 = roundReg_8_1_5;
  assign port_state_out_8_1_6 = roundReg_8_1_6;
  assign port_state_out_8_1_7 = roundReg_8_1_7;
  assign port_state_out_8_2_0 = roundReg_8_2_0;
  assign port_state_out_8_2_1 = roundReg_8_2_1;
  assign port_state_out_8_2_2 = roundReg_8_2_2;
  assign port_state_out_8_2_3 = roundReg_8_2_3;
  assign port_state_out_8_2_4 = roundReg_8_2_4;
  assign port_state_out_8_2_5 = roundReg_8_2_5;
  assign port_state_out_8_2_6 = roundReg_8_2_6;
  assign port_state_out_8_2_7 = roundReg_8_2_7;
  assign port_state_out_8_3_0 = roundReg_8_3_0;
  assign port_state_out_8_3_1 = roundReg_8_3_1;
  assign port_state_out_8_3_2 = roundReg_8_3_2;
  assign port_state_out_8_3_3 = roundReg_8_3_3;
  assign port_state_out_8_3_4 = roundReg_8_3_4;
  assign port_state_out_8_3_5 = roundReg_8_3_5;
  assign port_state_out_8_3_6 = roundReg_8_3_6;
  assign port_state_out_8_3_7 = roundReg_8_3_7;
  assign port_state_out_9_0_0 = roundReg_9_0_0;
  assign port_state_out_9_0_1 = roundReg_9_0_1;
  assign port_state_out_9_0_2 = roundReg_9_0_2;
  assign port_state_out_9_0_3 = roundReg_9_0_3;
  assign port_state_out_9_0_4 = roundReg_9_0_4;
  assign port_state_out_9_0_5 = roundReg_9_0_5;
  assign port_state_out_9_0_6 = roundReg_9_0_6;
  assign port_state_out_9_0_7 = roundReg_9_0_7;
  assign port_state_out_9_1_0 = roundReg_9_1_0;
  assign port_state_out_9_1_1 = roundReg_9_1_1;
  assign port_state_out_9_1_2 = roundReg_9_1_2;
  assign port_state_out_9_1_3 = roundReg_9_1_3;
  assign port_state_out_9_1_4 = roundReg_9_1_4;
  assign port_state_out_9_1_5 = roundReg_9_1_5;
  assign port_state_out_9_1_6 = roundReg_9_1_6;
  assign port_state_out_9_1_7 = roundReg_9_1_7;
  assign port_state_out_9_2_0 = roundReg_9_2_0;
  assign port_state_out_9_2_1 = roundReg_9_2_1;
  assign port_state_out_9_2_2 = roundReg_9_2_2;
  assign port_state_out_9_2_3 = roundReg_9_2_3;
  assign port_state_out_9_2_4 = roundReg_9_2_4;
  assign port_state_out_9_2_5 = roundReg_9_2_5;
  assign port_state_out_9_2_6 = roundReg_9_2_6;
  assign port_state_out_9_2_7 = roundReg_9_2_7;
  assign port_state_out_9_3_0 = roundReg_9_3_0;
  assign port_state_out_9_3_1 = roundReg_9_3_1;
  assign port_state_out_9_3_2 = roundReg_9_3_2;
  assign port_state_out_9_3_3 = roundReg_9_3_3;
  assign port_state_out_9_3_4 = roundReg_9_3_4;
  assign port_state_out_9_3_5 = roundReg_9_3_5;
  assign port_state_out_9_3_6 = roundReg_9_3_6;
  assign port_state_out_9_3_7 = roundReg_9_3_7;
  assign port_state_out_10_0_0 = roundReg_10_0_0;
  assign port_state_out_10_0_1 = roundReg_10_0_1;
  assign port_state_out_10_0_2 = roundReg_10_0_2;
  assign port_state_out_10_0_3 = roundReg_10_0_3;
  assign port_state_out_10_0_4 = roundReg_10_0_4;
  assign port_state_out_10_0_5 = roundReg_10_0_5;
  assign port_state_out_10_0_6 = roundReg_10_0_6;
  assign port_state_out_10_0_7 = roundReg_10_0_7;
  assign port_state_out_10_1_0 = roundReg_10_1_0;
  assign port_state_out_10_1_1 = roundReg_10_1_1;
  assign port_state_out_10_1_2 = roundReg_10_1_2;
  assign port_state_out_10_1_3 = roundReg_10_1_3;
  assign port_state_out_10_1_4 = roundReg_10_1_4;
  assign port_state_out_10_1_5 = roundReg_10_1_5;
  assign port_state_out_10_1_6 = roundReg_10_1_6;
  assign port_state_out_10_1_7 = roundReg_10_1_7;
  assign port_state_out_10_2_0 = roundReg_10_2_0;
  assign port_state_out_10_2_1 = roundReg_10_2_1;
  assign port_state_out_10_2_2 = roundReg_10_2_2;
  assign port_state_out_10_2_3 = roundReg_10_2_3;
  assign port_state_out_10_2_4 = roundReg_10_2_4;
  assign port_state_out_10_2_5 = roundReg_10_2_5;
  assign port_state_out_10_2_6 = roundReg_10_2_6;
  assign port_state_out_10_2_7 = roundReg_10_2_7;
  assign port_state_out_10_3_0 = roundReg_10_3_0;
  assign port_state_out_10_3_1 = roundReg_10_3_1;
  assign port_state_out_10_3_2 = roundReg_10_3_2;
  assign port_state_out_10_3_3 = roundReg_10_3_3;
  assign port_state_out_10_3_4 = roundReg_10_3_4;
  assign port_state_out_10_3_5 = roundReg_10_3_5;
  assign port_state_out_10_3_6 = roundReg_10_3_6;
  assign port_state_out_10_3_7 = roundReg_10_3_7;
  assign port_state_out_11_0_0 = roundReg_11_0_0;
  assign port_state_out_11_0_1 = roundReg_11_0_1;
  assign port_state_out_11_0_2 = roundReg_11_0_2;
  assign port_state_out_11_0_3 = roundReg_11_0_3;
  assign port_state_out_11_0_4 = roundReg_11_0_4;
  assign port_state_out_11_0_5 = roundReg_11_0_5;
  assign port_state_out_11_0_6 = roundReg_11_0_6;
  assign port_state_out_11_0_7 = roundReg_11_0_7;
  assign port_state_out_11_1_0 = roundReg_11_1_0;
  assign port_state_out_11_1_1 = roundReg_11_1_1;
  assign port_state_out_11_1_2 = roundReg_11_1_2;
  assign port_state_out_11_1_3 = roundReg_11_1_3;
  assign port_state_out_11_1_4 = roundReg_11_1_4;
  assign port_state_out_11_1_5 = roundReg_11_1_5;
  assign port_state_out_11_1_6 = roundReg_11_1_6;
  assign port_state_out_11_1_7 = roundReg_11_1_7;
  assign port_state_out_11_2_0 = roundReg_11_2_0;
  assign port_state_out_11_2_1 = roundReg_11_2_1;
  assign port_state_out_11_2_2 = roundReg_11_2_2;
  assign port_state_out_11_2_3 = roundReg_11_2_3;
  assign port_state_out_11_2_4 = roundReg_11_2_4;
  assign port_state_out_11_2_5 = roundReg_11_2_5;
  assign port_state_out_11_2_6 = roundReg_11_2_6;
  assign port_state_out_11_2_7 = roundReg_11_2_7;
  assign port_state_out_11_3_0 = roundReg_11_3_0;
  assign port_state_out_11_3_1 = roundReg_11_3_1;
  assign port_state_out_11_3_2 = roundReg_11_3_2;
  assign port_state_out_11_3_3 = roundReg_11_3_3;
  assign port_state_out_11_3_4 = roundReg_11_3_4;
  assign port_state_out_11_3_5 = roundReg_11_3_5;
  assign port_state_out_11_3_6 = roundReg_11_3_6;
  assign port_state_out_11_3_7 = roundReg_11_3_7;
  assign port_state_out_12_0_0 = roundReg_12_0_0;
  assign port_state_out_12_0_1 = roundReg_12_0_1;
  assign port_state_out_12_0_2 = roundReg_12_0_2;
  assign port_state_out_12_0_3 = roundReg_12_0_3;
  assign port_state_out_12_0_4 = roundReg_12_0_4;
  assign port_state_out_12_0_5 = roundReg_12_0_5;
  assign port_state_out_12_0_6 = roundReg_12_0_6;
  assign port_state_out_12_0_7 = roundReg_12_0_7;
  assign port_state_out_12_1_0 = roundReg_12_1_0;
  assign port_state_out_12_1_1 = roundReg_12_1_1;
  assign port_state_out_12_1_2 = roundReg_12_1_2;
  assign port_state_out_12_1_3 = roundReg_12_1_3;
  assign port_state_out_12_1_4 = roundReg_12_1_4;
  assign port_state_out_12_1_5 = roundReg_12_1_5;
  assign port_state_out_12_1_6 = roundReg_12_1_6;
  assign port_state_out_12_1_7 = roundReg_12_1_7;
  assign port_state_out_12_2_0 = roundReg_12_2_0;
  assign port_state_out_12_2_1 = roundReg_12_2_1;
  assign port_state_out_12_2_2 = roundReg_12_2_2;
  assign port_state_out_12_2_3 = roundReg_12_2_3;
  assign port_state_out_12_2_4 = roundReg_12_2_4;
  assign port_state_out_12_2_5 = roundReg_12_2_5;
  assign port_state_out_12_2_6 = roundReg_12_2_6;
  assign port_state_out_12_2_7 = roundReg_12_2_7;
  assign port_state_out_12_3_0 = roundReg_12_3_0;
  assign port_state_out_12_3_1 = roundReg_12_3_1;
  assign port_state_out_12_3_2 = roundReg_12_3_2;
  assign port_state_out_12_3_3 = roundReg_12_3_3;
  assign port_state_out_12_3_4 = roundReg_12_3_4;
  assign port_state_out_12_3_5 = roundReg_12_3_5;
  assign port_state_out_12_3_6 = roundReg_12_3_6;
  assign port_state_out_12_3_7 = roundReg_12_3_7;
  assign port_state_out_13_0_0 = roundReg_13_0_0;
  assign port_state_out_13_0_1 = roundReg_13_0_1;
  assign port_state_out_13_0_2 = roundReg_13_0_2;
  assign port_state_out_13_0_3 = roundReg_13_0_3;
  assign port_state_out_13_0_4 = roundReg_13_0_4;
  assign port_state_out_13_0_5 = roundReg_13_0_5;
  assign port_state_out_13_0_6 = roundReg_13_0_6;
  assign port_state_out_13_0_7 = roundReg_13_0_7;
  assign port_state_out_13_1_0 = roundReg_13_1_0;
  assign port_state_out_13_1_1 = roundReg_13_1_1;
  assign port_state_out_13_1_2 = roundReg_13_1_2;
  assign port_state_out_13_1_3 = roundReg_13_1_3;
  assign port_state_out_13_1_4 = roundReg_13_1_4;
  assign port_state_out_13_1_5 = roundReg_13_1_5;
  assign port_state_out_13_1_6 = roundReg_13_1_6;
  assign port_state_out_13_1_7 = roundReg_13_1_7;
  assign port_state_out_13_2_0 = roundReg_13_2_0;
  assign port_state_out_13_2_1 = roundReg_13_2_1;
  assign port_state_out_13_2_2 = roundReg_13_2_2;
  assign port_state_out_13_2_3 = roundReg_13_2_3;
  assign port_state_out_13_2_4 = roundReg_13_2_4;
  assign port_state_out_13_2_5 = roundReg_13_2_5;
  assign port_state_out_13_2_6 = roundReg_13_2_6;
  assign port_state_out_13_2_7 = roundReg_13_2_7;
  assign port_state_out_13_3_0 = roundReg_13_3_0;
  assign port_state_out_13_3_1 = roundReg_13_3_1;
  assign port_state_out_13_3_2 = roundReg_13_3_2;
  assign port_state_out_13_3_3 = roundReg_13_3_3;
  assign port_state_out_13_3_4 = roundReg_13_3_4;
  assign port_state_out_13_3_5 = roundReg_13_3_5;
  assign port_state_out_13_3_6 = roundReg_13_3_6;
  assign port_state_out_13_3_7 = roundReg_13_3_7;
  assign port_state_out_14_0_0 = roundReg_14_0_0;
  assign port_state_out_14_0_1 = roundReg_14_0_1;
  assign port_state_out_14_0_2 = roundReg_14_0_2;
  assign port_state_out_14_0_3 = roundReg_14_0_3;
  assign port_state_out_14_0_4 = roundReg_14_0_4;
  assign port_state_out_14_0_5 = roundReg_14_0_5;
  assign port_state_out_14_0_6 = roundReg_14_0_6;
  assign port_state_out_14_0_7 = roundReg_14_0_7;
  assign port_state_out_14_1_0 = roundReg_14_1_0;
  assign port_state_out_14_1_1 = roundReg_14_1_1;
  assign port_state_out_14_1_2 = roundReg_14_1_2;
  assign port_state_out_14_1_3 = roundReg_14_1_3;
  assign port_state_out_14_1_4 = roundReg_14_1_4;
  assign port_state_out_14_1_5 = roundReg_14_1_5;
  assign port_state_out_14_1_6 = roundReg_14_1_6;
  assign port_state_out_14_1_7 = roundReg_14_1_7;
  assign port_state_out_14_2_0 = roundReg_14_2_0;
  assign port_state_out_14_2_1 = roundReg_14_2_1;
  assign port_state_out_14_2_2 = roundReg_14_2_2;
  assign port_state_out_14_2_3 = roundReg_14_2_3;
  assign port_state_out_14_2_4 = roundReg_14_2_4;
  assign port_state_out_14_2_5 = roundReg_14_2_5;
  assign port_state_out_14_2_6 = roundReg_14_2_6;
  assign port_state_out_14_2_7 = roundReg_14_2_7;
  assign port_state_out_14_3_0 = roundReg_14_3_0;
  assign port_state_out_14_3_1 = roundReg_14_3_1;
  assign port_state_out_14_3_2 = roundReg_14_3_2;
  assign port_state_out_14_3_3 = roundReg_14_3_3;
  assign port_state_out_14_3_4 = roundReg_14_3_4;
  assign port_state_out_14_3_5 = roundReg_14_3_5;
  assign port_state_out_14_3_6 = roundReg_14_3_6;
  assign port_state_out_14_3_7 = roundReg_14_3_7;
  assign port_state_out_15_0_0 = roundReg_15_0_0;
  assign port_state_out_15_0_1 = roundReg_15_0_1;
  assign port_state_out_15_0_2 = roundReg_15_0_2;
  assign port_state_out_15_0_3 = roundReg_15_0_3;
  assign port_state_out_15_0_4 = roundReg_15_0_4;
  assign port_state_out_15_0_5 = roundReg_15_0_5;
  assign port_state_out_15_0_6 = roundReg_15_0_6;
  assign port_state_out_15_0_7 = roundReg_15_0_7;
  assign port_state_out_15_1_0 = roundReg_15_1_0;
  assign port_state_out_15_1_1 = roundReg_15_1_1;
  assign port_state_out_15_1_2 = roundReg_15_1_2;
  assign port_state_out_15_1_3 = roundReg_15_1_3;
  assign port_state_out_15_1_4 = roundReg_15_1_4;
  assign port_state_out_15_1_5 = roundReg_15_1_5;
  assign port_state_out_15_1_6 = roundReg_15_1_6;
  assign port_state_out_15_1_7 = roundReg_15_1_7;
  assign port_state_out_15_2_0 = roundReg_15_2_0;
  assign port_state_out_15_2_1 = roundReg_15_2_1;
  assign port_state_out_15_2_2 = roundReg_15_2_2;
  assign port_state_out_15_2_3 = roundReg_15_2_3;
  assign port_state_out_15_2_4 = roundReg_15_2_4;
  assign port_state_out_15_2_5 = roundReg_15_2_5;
  assign port_state_out_15_2_6 = roundReg_15_2_6;
  assign port_state_out_15_2_7 = roundReg_15_2_7;
  assign port_state_out_15_3_0 = roundReg_15_3_0;
  assign port_state_out_15_3_1 = roundReg_15_3_1;
  assign port_state_out_15_3_2 = roundReg_15_3_2;
  assign port_state_out_15_3_3 = roundReg_15_3_3;
  assign port_state_out_15_3_4 = roundReg_15_3_4;
  assign port_state_out_15_3_5 = roundReg_15_3_5;
  assign port_state_out_15_3_6 = roundReg_15_3_6;
  assign port_state_out_15_3_7 = roundReg_15_3_7;
  always @(posedge clk) begin
    roundReg_0_0_0[0] <= majority_4608_port_o;
    roundReg_1_0_0[0] <= majority_4609_port_o;
    roundReg_2_0_0[0] <= majority_4610_port_o;
    roundReg_3_0_0[0] <= majority_4611_port_o;
    roundReg_4_0_0[0] <= majority_4612_port_o;
    roundReg_5_0_0[0] <= majority_4613_port_o;
    roundReg_6_0_0[0] <= majority_4614_port_o;
    roundReg_7_0_0[0] <= majority_4615_port_o;
    roundReg_8_0_0[0] <= majority_4616_port_o;
    roundReg_9_0_0[0] <= majority_4617_port_o;
    roundReg_10_0_0[0] <= majority_4618_port_o;
    roundReg_11_0_0[0] <= majority_4619_port_o;
    roundReg_12_0_0[0] <= majority_4620_port_o;
    roundReg_13_0_0[0] <= majority_4621_port_o;
    roundReg_14_0_0[0] <= majority_4622_port_o;
    roundReg_15_0_0[0] <= majority_4623_port_o;
    roundReg_0_1_0[0] <= majority_4624_port_o;
    roundReg_1_1_0[0] <= majority_4625_port_o;
    roundReg_2_1_0[0] <= majority_4626_port_o;
    roundReg_3_1_0[0] <= majority_4627_port_o;
    roundReg_4_1_0[0] <= majority_4628_port_o;
    roundReg_5_1_0[0] <= majority_4629_port_o;
    roundReg_6_1_0[0] <= majority_4630_port_o;
    roundReg_7_1_0[0] <= majority_4631_port_o;
    roundReg_8_1_0[0] <= majority_4632_port_o;
    roundReg_9_1_0[0] <= majority_4633_port_o;
    roundReg_10_1_0[0] <= majority_4634_port_o;
    roundReg_11_1_0[0] <= majority_4635_port_o;
    roundReg_12_1_0[0] <= majority_4636_port_o;
    roundReg_13_1_0[0] <= majority_4637_port_o;
    roundReg_14_1_0[0] <= majority_4638_port_o;
    roundReg_15_1_0[0] <= majority_4639_port_o;
    roundReg_0_2_0[0] <= majority_4640_port_o;
    roundReg_1_2_0[0] <= majority_4641_port_o;
    roundReg_2_2_0[0] <= majority_4642_port_o;
    roundReg_3_2_0[0] <= majority_4643_port_o;
    roundReg_4_2_0[0] <= majority_4644_port_o;
    roundReg_5_2_0[0] <= majority_4645_port_o;
    roundReg_6_2_0[0] <= majority_4646_port_o;
    roundReg_7_2_0[0] <= majority_4647_port_o;
    roundReg_8_2_0[0] <= majority_4648_port_o;
    roundReg_9_2_0[0] <= majority_4649_port_o;
    roundReg_10_2_0[0] <= majority_4650_port_o;
    roundReg_11_2_0[0] <= majority_4651_port_o;
    roundReg_12_2_0[0] <= majority_4652_port_o;
    roundReg_13_2_0[0] <= majority_4653_port_o;
    roundReg_14_2_0[0] <= majority_4654_port_o;
    roundReg_15_2_0[0] <= majority_4655_port_o;
    roundReg_0_3_0[0] <= majority_4656_port_o;
    roundReg_1_3_0[0] <= majority_4657_port_o;
    roundReg_2_3_0[0] <= majority_4658_port_o;
    roundReg_3_3_0[0] <= majority_4659_port_o;
    roundReg_4_3_0[0] <= majority_4660_port_o;
    roundReg_5_3_0[0] <= majority_4661_port_o;
    roundReg_6_3_0[0] <= majority_4662_port_o;
    roundReg_7_3_0[0] <= majority_4663_port_o;
    roundReg_8_3_0[0] <= majority_4664_port_o;
    roundReg_9_3_0[0] <= majority_4665_port_o;
    roundReg_10_3_0[0] <= majority_4666_port_o;
    roundReg_11_3_0[0] <= majority_4667_port_o;
    roundReg_12_3_0[0] <= majority_4668_port_o;
    roundReg_13_3_0[0] <= majority_4669_port_o;
    roundReg_14_3_0[0] <= majority_4670_port_o;
    roundReg_15_3_0[0] <= majority_4671_port_o;
    roundReg_0_0_1[0] <= majority_4672_port_o;
    roundReg_1_0_1[0] <= majority_4673_port_o;
    roundReg_2_0_1[0] <= majority_4674_port_o;
    roundReg_3_0_1[0] <= majority_4675_port_o;
    roundReg_4_0_1[0] <= majority_4676_port_o;
    roundReg_5_0_1[0] <= majority_4677_port_o;
    roundReg_6_0_1[0] <= majority_4678_port_o;
    roundReg_7_0_1[0] <= majority_4679_port_o;
    roundReg_8_0_1[0] <= majority_4680_port_o;
    roundReg_9_0_1[0] <= majority_4681_port_o;
    roundReg_10_0_1[0] <= majority_4682_port_o;
    roundReg_11_0_1[0] <= majority_4683_port_o;
    roundReg_12_0_1[0] <= majority_4684_port_o;
    roundReg_13_0_1[0] <= majority_4685_port_o;
    roundReg_14_0_1[0] <= majority_4686_port_o;
    roundReg_15_0_1[0] <= majority_4687_port_o;
    roundReg_0_1_1[0] <= majority_4688_port_o;
    roundReg_1_1_1[0] <= majority_4689_port_o;
    roundReg_2_1_1[0] <= majority_4690_port_o;
    roundReg_3_1_1[0] <= majority_4691_port_o;
    roundReg_4_1_1[0] <= majority_4692_port_o;
    roundReg_5_1_1[0] <= majority_4693_port_o;
    roundReg_6_1_1[0] <= majority_4694_port_o;
    roundReg_7_1_1[0] <= majority_4695_port_o;
    roundReg_8_1_1[0] <= majority_4696_port_o;
    roundReg_9_1_1[0] <= majority_4697_port_o;
    roundReg_10_1_1[0] <= majority_4698_port_o;
    roundReg_11_1_1[0] <= majority_4699_port_o;
    roundReg_12_1_1[0] <= majority_4700_port_o;
    roundReg_13_1_1[0] <= majority_4701_port_o;
    roundReg_14_1_1[0] <= majority_4702_port_o;
    roundReg_15_1_1[0] <= majority_4703_port_o;
    roundReg_0_2_1[0] <= majority_4704_port_o;
    roundReg_1_2_1[0] <= majority_4705_port_o;
    roundReg_2_2_1[0] <= majority_4706_port_o;
    roundReg_3_2_1[0] <= majority_4707_port_o;
    roundReg_4_2_1[0] <= majority_4708_port_o;
    roundReg_5_2_1[0] <= majority_4709_port_o;
    roundReg_6_2_1[0] <= majority_4710_port_o;
    roundReg_7_2_1[0] <= majority_4711_port_o;
    roundReg_8_2_1[0] <= majority_4712_port_o;
    roundReg_9_2_1[0] <= majority_4713_port_o;
    roundReg_10_2_1[0] <= majority_4714_port_o;
    roundReg_11_2_1[0] <= majority_4715_port_o;
    roundReg_12_2_1[0] <= majority_4716_port_o;
    roundReg_13_2_1[0] <= majority_4717_port_o;
    roundReg_14_2_1[0] <= majority_4718_port_o;
    roundReg_15_2_1[0] <= majority_4719_port_o;
    roundReg_0_3_1[0] <= majority_4720_port_o;
    roundReg_1_3_1[0] <= majority_4721_port_o;
    roundReg_2_3_1[0] <= majority_4722_port_o;
    roundReg_3_3_1[0] <= majority_4723_port_o;
    roundReg_4_3_1[0] <= majority_4724_port_o;
    roundReg_5_3_1[0] <= majority_4725_port_o;
    roundReg_6_3_1[0] <= majority_4726_port_o;
    roundReg_7_3_1[0] <= majority_4727_port_o;
    roundReg_8_3_1[0] <= majority_4728_port_o;
    roundReg_9_3_1[0] <= majority_4729_port_o;
    roundReg_10_3_1[0] <= majority_4730_port_o;
    roundReg_11_3_1[0] <= majority_4731_port_o;
    roundReg_12_3_1[0] <= majority_4732_port_o;
    roundReg_13_3_1[0] <= majority_4733_port_o;
    roundReg_14_3_1[0] <= majority_4734_port_o;
    roundReg_15_3_1[0] <= majority_4735_port_o;
    roundReg_0_0_2[0] <= majority_4736_port_o;
    roundReg_1_0_2[0] <= majority_4737_port_o;
    roundReg_2_0_2[0] <= majority_4738_port_o;
    roundReg_3_0_2[0] <= majority_4739_port_o;
    roundReg_4_0_2[0] <= majority_4740_port_o;
    roundReg_5_0_2[0] <= majority_4741_port_o;
    roundReg_6_0_2[0] <= majority_4742_port_o;
    roundReg_7_0_2[0] <= majority_4743_port_o;
    roundReg_8_0_2[0] <= majority_4744_port_o;
    roundReg_9_0_2[0] <= majority_4745_port_o;
    roundReg_10_0_2[0] <= majority_4746_port_o;
    roundReg_11_0_2[0] <= majority_4747_port_o;
    roundReg_12_0_2[0] <= majority_4748_port_o;
    roundReg_13_0_2[0] <= majority_4749_port_o;
    roundReg_14_0_2[0] <= majority_4750_port_o;
    roundReg_15_0_2[0] <= majority_4751_port_o;
    roundReg_0_1_2[0] <= majority_4752_port_o;
    roundReg_1_1_2[0] <= majority_4753_port_o;
    roundReg_2_1_2[0] <= majority_4754_port_o;
    roundReg_3_1_2[0] <= majority_4755_port_o;
    roundReg_4_1_2[0] <= majority_4756_port_o;
    roundReg_5_1_2[0] <= majority_4757_port_o;
    roundReg_6_1_2[0] <= majority_4758_port_o;
    roundReg_7_1_2[0] <= majority_4759_port_o;
    roundReg_8_1_2[0] <= majority_4760_port_o;
    roundReg_9_1_2[0] <= majority_4761_port_o;
    roundReg_10_1_2[0] <= majority_4762_port_o;
    roundReg_11_1_2[0] <= majority_4763_port_o;
    roundReg_12_1_2[0] <= majority_4764_port_o;
    roundReg_13_1_2[0] <= majority_4765_port_o;
    roundReg_14_1_2[0] <= majority_4766_port_o;
    roundReg_15_1_2[0] <= majority_4767_port_o;
    roundReg_0_2_2[0] <= majority_4768_port_o;
    roundReg_1_2_2[0] <= majority_4769_port_o;
    roundReg_2_2_2[0] <= majority_4770_port_o;
    roundReg_3_2_2[0] <= majority_4771_port_o;
    roundReg_4_2_2[0] <= majority_4772_port_o;
    roundReg_5_2_2[0] <= majority_4773_port_o;
    roundReg_6_2_2[0] <= majority_4774_port_o;
    roundReg_7_2_2[0] <= majority_4775_port_o;
    roundReg_8_2_2[0] <= majority_4776_port_o;
    roundReg_9_2_2[0] <= majority_4777_port_o;
    roundReg_10_2_2[0] <= majority_4778_port_o;
    roundReg_11_2_2[0] <= majority_4779_port_o;
    roundReg_12_2_2[0] <= majority_4780_port_o;
    roundReg_13_2_2[0] <= majority_4781_port_o;
    roundReg_14_2_2[0] <= majority_4782_port_o;
    roundReg_15_2_2[0] <= majority_4783_port_o;
    roundReg_0_3_2[0] <= majority_4784_port_o;
    roundReg_1_3_2[0] <= majority_4785_port_o;
    roundReg_2_3_2[0] <= majority_4786_port_o;
    roundReg_3_3_2[0] <= majority_4787_port_o;
    roundReg_4_3_2[0] <= majority_4788_port_o;
    roundReg_5_3_2[0] <= majority_4789_port_o;
    roundReg_6_3_2[0] <= majority_4790_port_o;
    roundReg_7_3_2[0] <= majority_4791_port_o;
    roundReg_8_3_2[0] <= majority_4792_port_o;
    roundReg_9_3_2[0] <= majority_4793_port_o;
    roundReg_10_3_2[0] <= majority_4794_port_o;
    roundReg_11_3_2[0] <= majority_4795_port_o;
    roundReg_12_3_2[0] <= majority_4796_port_o;
    roundReg_13_3_2[0] <= majority_4797_port_o;
    roundReg_14_3_2[0] <= majority_4798_port_o;
    roundReg_15_3_2[0] <= majority_4799_port_o;
    roundReg_0_0_3[0] <= majority_4800_port_o;
    roundReg_1_0_3[0] <= majority_4801_port_o;
    roundReg_2_0_3[0] <= majority_4802_port_o;
    roundReg_3_0_3[0] <= majority_4803_port_o;
    roundReg_4_0_3[0] <= majority_4804_port_o;
    roundReg_5_0_3[0] <= majority_4805_port_o;
    roundReg_6_0_3[0] <= majority_4806_port_o;
    roundReg_7_0_3[0] <= majority_4807_port_o;
    roundReg_8_0_3[0] <= majority_4808_port_o;
    roundReg_9_0_3[0] <= majority_4809_port_o;
    roundReg_10_0_3[0] <= majority_4810_port_o;
    roundReg_11_0_3[0] <= majority_4811_port_o;
    roundReg_12_0_3[0] <= majority_4812_port_o;
    roundReg_13_0_3[0] <= majority_4813_port_o;
    roundReg_14_0_3[0] <= majority_4814_port_o;
    roundReg_15_0_3[0] <= majority_4815_port_o;
    roundReg_0_1_3[0] <= majority_4816_port_o;
    roundReg_1_1_3[0] <= majority_4817_port_o;
    roundReg_2_1_3[0] <= majority_4818_port_o;
    roundReg_3_1_3[0] <= majority_4819_port_o;
    roundReg_4_1_3[0] <= majority_4820_port_o;
    roundReg_5_1_3[0] <= majority_4821_port_o;
    roundReg_6_1_3[0] <= majority_4822_port_o;
    roundReg_7_1_3[0] <= majority_4823_port_o;
    roundReg_8_1_3[0] <= majority_4824_port_o;
    roundReg_9_1_3[0] <= majority_4825_port_o;
    roundReg_10_1_3[0] <= majority_4826_port_o;
    roundReg_11_1_3[0] <= majority_4827_port_o;
    roundReg_12_1_3[0] <= majority_4828_port_o;
    roundReg_13_1_3[0] <= majority_4829_port_o;
    roundReg_14_1_3[0] <= majority_4830_port_o;
    roundReg_15_1_3[0] <= majority_4831_port_o;
    roundReg_0_2_3[0] <= majority_4832_port_o;
    roundReg_1_2_3[0] <= majority_4833_port_o;
    roundReg_2_2_3[0] <= majority_4834_port_o;
    roundReg_3_2_3[0] <= majority_4835_port_o;
    roundReg_4_2_3[0] <= majority_4836_port_o;
    roundReg_5_2_3[0] <= majority_4837_port_o;
    roundReg_6_2_3[0] <= majority_4838_port_o;
    roundReg_7_2_3[0] <= majority_4839_port_o;
    roundReg_8_2_3[0] <= majority_4840_port_o;
    roundReg_9_2_3[0] <= majority_4841_port_o;
    roundReg_10_2_3[0] <= majority_4842_port_o;
    roundReg_11_2_3[0] <= majority_4843_port_o;
    roundReg_12_2_3[0] <= majority_4844_port_o;
    roundReg_13_2_3[0] <= majority_4845_port_o;
    roundReg_14_2_3[0] <= majority_4846_port_o;
    roundReg_15_2_3[0] <= majority_4847_port_o;
    roundReg_0_3_3[0] <= majority_4848_port_o;
    roundReg_1_3_3[0] <= majority_4849_port_o;
    roundReg_2_3_3[0] <= majority_4850_port_o;
    roundReg_3_3_3[0] <= majority_4851_port_o;
    roundReg_4_3_3[0] <= majority_4852_port_o;
    roundReg_5_3_3[0] <= majority_4853_port_o;
    roundReg_6_3_3[0] <= majority_4854_port_o;
    roundReg_7_3_3[0] <= majority_4855_port_o;
    roundReg_8_3_3[0] <= majority_4856_port_o;
    roundReg_9_3_3[0] <= majority_4857_port_o;
    roundReg_10_3_3[0] <= majority_4858_port_o;
    roundReg_11_3_3[0] <= majority_4859_port_o;
    roundReg_12_3_3[0] <= majority_4860_port_o;
    roundReg_13_3_3[0] <= majority_4861_port_o;
    roundReg_14_3_3[0] <= majority_4862_port_o;
    roundReg_15_3_3[0] <= majority_4863_port_o;
    roundReg_0_0_4[0] <= majority_4864_port_o;
    roundReg_1_0_4[0] <= majority_4865_port_o;
    roundReg_2_0_4[0] <= majority_4866_port_o;
    roundReg_3_0_4[0] <= majority_4867_port_o;
    roundReg_4_0_4[0] <= majority_4868_port_o;
    roundReg_5_0_4[0] <= majority_4869_port_o;
    roundReg_6_0_4[0] <= majority_4870_port_o;
    roundReg_7_0_4[0] <= majority_4871_port_o;
    roundReg_8_0_4[0] <= majority_4872_port_o;
    roundReg_9_0_4[0] <= majority_4873_port_o;
    roundReg_10_0_4[0] <= majority_4874_port_o;
    roundReg_11_0_4[0] <= majority_4875_port_o;
    roundReg_12_0_4[0] <= majority_4876_port_o;
    roundReg_13_0_4[0] <= majority_4877_port_o;
    roundReg_14_0_4[0] <= majority_4878_port_o;
    roundReg_15_0_4[0] <= majority_4879_port_o;
    roundReg_0_1_4[0] <= majority_4880_port_o;
    roundReg_1_1_4[0] <= majority_4881_port_o;
    roundReg_2_1_4[0] <= majority_4882_port_o;
    roundReg_3_1_4[0] <= majority_4883_port_o;
    roundReg_4_1_4[0] <= majority_4884_port_o;
    roundReg_5_1_4[0] <= majority_4885_port_o;
    roundReg_6_1_4[0] <= majority_4886_port_o;
    roundReg_7_1_4[0] <= majority_4887_port_o;
    roundReg_8_1_4[0] <= majority_4888_port_o;
    roundReg_9_1_4[0] <= majority_4889_port_o;
    roundReg_10_1_4[0] <= majority_4890_port_o;
    roundReg_11_1_4[0] <= majority_4891_port_o;
    roundReg_12_1_4[0] <= majority_4892_port_o;
    roundReg_13_1_4[0] <= majority_4893_port_o;
    roundReg_14_1_4[0] <= majority_4894_port_o;
    roundReg_15_1_4[0] <= majority_4895_port_o;
    roundReg_0_2_4[0] <= majority_4896_port_o;
    roundReg_1_2_4[0] <= majority_4897_port_o;
    roundReg_2_2_4[0] <= majority_4898_port_o;
    roundReg_3_2_4[0] <= majority_4899_port_o;
    roundReg_4_2_4[0] <= majority_4900_port_o;
    roundReg_5_2_4[0] <= majority_4901_port_o;
    roundReg_6_2_4[0] <= majority_4902_port_o;
    roundReg_7_2_4[0] <= majority_4903_port_o;
    roundReg_8_2_4[0] <= majority_4904_port_o;
    roundReg_9_2_4[0] <= majority_4905_port_o;
    roundReg_10_2_4[0] <= majority_4906_port_o;
    roundReg_11_2_4[0] <= majority_4907_port_o;
    roundReg_12_2_4[0] <= majority_4908_port_o;
    roundReg_13_2_4[0] <= majority_4909_port_o;
    roundReg_14_2_4[0] <= majority_4910_port_o;
    roundReg_15_2_4[0] <= majority_4911_port_o;
    roundReg_0_3_4[0] <= majority_4912_port_o;
    roundReg_1_3_4[0] <= majority_4913_port_o;
    roundReg_2_3_4[0] <= majority_4914_port_o;
    roundReg_3_3_4[0] <= majority_4915_port_o;
    roundReg_4_3_4[0] <= majority_4916_port_o;
    roundReg_5_3_4[0] <= majority_4917_port_o;
    roundReg_6_3_4[0] <= majority_4918_port_o;
    roundReg_7_3_4[0] <= majority_4919_port_o;
    roundReg_8_3_4[0] <= majority_4920_port_o;
    roundReg_9_3_4[0] <= majority_4921_port_o;
    roundReg_10_3_4[0] <= majority_4922_port_o;
    roundReg_11_3_4[0] <= majority_4923_port_o;
    roundReg_12_3_4[0] <= majority_4924_port_o;
    roundReg_13_3_4[0] <= majority_4925_port_o;
    roundReg_14_3_4[0] <= majority_4926_port_o;
    roundReg_15_3_4[0] <= majority_4927_port_o;
    roundReg_0_0_5[0] <= majority_4928_port_o;
    roundReg_1_0_5[0] <= majority_4929_port_o;
    roundReg_2_0_5[0] <= majority_4930_port_o;
    roundReg_3_0_5[0] <= majority_4931_port_o;
    roundReg_4_0_5[0] <= majority_4932_port_o;
    roundReg_5_0_5[0] <= majority_4933_port_o;
    roundReg_6_0_5[0] <= majority_4934_port_o;
    roundReg_7_0_5[0] <= majority_4935_port_o;
    roundReg_8_0_5[0] <= majority_4936_port_o;
    roundReg_9_0_5[0] <= majority_4937_port_o;
    roundReg_10_0_5[0] <= majority_4938_port_o;
    roundReg_11_0_5[0] <= majority_4939_port_o;
    roundReg_12_0_5[0] <= majority_4940_port_o;
    roundReg_13_0_5[0] <= majority_4941_port_o;
    roundReg_14_0_5[0] <= majority_4942_port_o;
    roundReg_15_0_5[0] <= majority_4943_port_o;
    roundReg_0_1_5[0] <= majority_4944_port_o;
    roundReg_1_1_5[0] <= majority_4945_port_o;
    roundReg_2_1_5[0] <= majority_4946_port_o;
    roundReg_3_1_5[0] <= majority_4947_port_o;
    roundReg_4_1_5[0] <= majority_4948_port_o;
    roundReg_5_1_5[0] <= majority_4949_port_o;
    roundReg_6_1_5[0] <= majority_4950_port_o;
    roundReg_7_1_5[0] <= majority_4951_port_o;
    roundReg_8_1_5[0] <= majority_4952_port_o;
    roundReg_9_1_5[0] <= majority_4953_port_o;
    roundReg_10_1_5[0] <= majority_4954_port_o;
    roundReg_11_1_5[0] <= majority_4955_port_o;
    roundReg_12_1_5[0] <= majority_4956_port_o;
    roundReg_13_1_5[0] <= majority_4957_port_o;
    roundReg_14_1_5[0] <= majority_4958_port_o;
    roundReg_15_1_5[0] <= majority_4959_port_o;
    roundReg_0_2_5[0] <= majority_4960_port_o;
    roundReg_1_2_5[0] <= majority_4961_port_o;
    roundReg_2_2_5[0] <= majority_4962_port_o;
    roundReg_3_2_5[0] <= majority_4963_port_o;
    roundReg_4_2_5[0] <= majority_4964_port_o;
    roundReg_5_2_5[0] <= majority_4965_port_o;
    roundReg_6_2_5[0] <= majority_4966_port_o;
    roundReg_7_2_5[0] <= majority_4967_port_o;
    roundReg_8_2_5[0] <= majority_4968_port_o;
    roundReg_9_2_5[0] <= majority_4969_port_o;
    roundReg_10_2_5[0] <= majority_4970_port_o;
    roundReg_11_2_5[0] <= majority_4971_port_o;
    roundReg_12_2_5[0] <= majority_4972_port_o;
    roundReg_13_2_5[0] <= majority_4973_port_o;
    roundReg_14_2_5[0] <= majority_4974_port_o;
    roundReg_15_2_5[0] <= majority_4975_port_o;
    roundReg_0_3_5[0] <= majority_4976_port_o;
    roundReg_1_3_5[0] <= majority_4977_port_o;
    roundReg_2_3_5[0] <= majority_4978_port_o;
    roundReg_3_3_5[0] <= majority_4979_port_o;
    roundReg_4_3_5[0] <= majority_4980_port_o;
    roundReg_5_3_5[0] <= majority_4981_port_o;
    roundReg_6_3_5[0] <= majority_4982_port_o;
    roundReg_7_3_5[0] <= majority_4983_port_o;
    roundReg_8_3_5[0] <= majority_4984_port_o;
    roundReg_9_3_5[0] <= majority_4985_port_o;
    roundReg_10_3_5[0] <= majority_4986_port_o;
    roundReg_11_3_5[0] <= majority_4987_port_o;
    roundReg_12_3_5[0] <= majority_4988_port_o;
    roundReg_13_3_5[0] <= majority_4989_port_o;
    roundReg_14_3_5[0] <= majority_4990_port_o;
    roundReg_15_3_5[0] <= majority_4991_port_o;
    roundReg_0_0_6[0] <= majority_4992_port_o;
    roundReg_1_0_6[0] <= majority_4993_port_o;
    roundReg_2_0_6[0] <= majority_4994_port_o;
    roundReg_3_0_6[0] <= majority_4995_port_o;
    roundReg_4_0_6[0] <= majority_4996_port_o;
    roundReg_5_0_6[0] <= majority_4997_port_o;
    roundReg_6_0_6[0] <= majority_4998_port_o;
    roundReg_7_0_6[0] <= majority_4999_port_o;
    roundReg_8_0_6[0] <= majority_5000_port_o;
    roundReg_9_0_6[0] <= majority_5001_port_o;
    roundReg_10_0_6[0] <= majority_5002_port_o;
    roundReg_11_0_6[0] <= majority_5003_port_o;
    roundReg_12_0_6[0] <= majority_5004_port_o;
    roundReg_13_0_6[0] <= majority_5005_port_o;
    roundReg_14_0_6[0] <= majority_5006_port_o;
    roundReg_15_0_6[0] <= majority_5007_port_o;
    roundReg_0_1_6[0] <= majority_5008_port_o;
    roundReg_1_1_6[0] <= majority_5009_port_o;
    roundReg_2_1_6[0] <= majority_5010_port_o;
    roundReg_3_1_6[0] <= majority_5011_port_o;
    roundReg_4_1_6[0] <= majority_5012_port_o;
    roundReg_5_1_6[0] <= majority_5013_port_o;
    roundReg_6_1_6[0] <= majority_5014_port_o;
    roundReg_7_1_6[0] <= majority_5015_port_o;
    roundReg_8_1_6[0] <= majority_5016_port_o;
    roundReg_9_1_6[0] <= majority_5017_port_o;
    roundReg_10_1_6[0] <= majority_5018_port_o;
    roundReg_11_1_6[0] <= majority_5019_port_o;
    roundReg_12_1_6[0] <= majority_5020_port_o;
    roundReg_13_1_6[0] <= majority_5021_port_o;
    roundReg_14_1_6[0] <= majority_5022_port_o;
    roundReg_15_1_6[0] <= majority_5023_port_o;
    roundReg_0_2_6[0] <= majority_5024_port_o;
    roundReg_1_2_6[0] <= majority_5025_port_o;
    roundReg_2_2_6[0] <= majority_5026_port_o;
    roundReg_3_2_6[0] <= majority_5027_port_o;
    roundReg_4_2_6[0] <= majority_5028_port_o;
    roundReg_5_2_6[0] <= majority_5029_port_o;
    roundReg_6_2_6[0] <= majority_5030_port_o;
    roundReg_7_2_6[0] <= majority_5031_port_o;
    roundReg_8_2_6[0] <= majority_5032_port_o;
    roundReg_9_2_6[0] <= majority_5033_port_o;
    roundReg_10_2_6[0] <= majority_5034_port_o;
    roundReg_11_2_6[0] <= majority_5035_port_o;
    roundReg_12_2_6[0] <= majority_5036_port_o;
    roundReg_13_2_6[0] <= majority_5037_port_o;
    roundReg_14_2_6[0] <= majority_5038_port_o;
    roundReg_15_2_6[0] <= majority_5039_port_o;
    roundReg_0_3_6[0] <= majority_5040_port_o;
    roundReg_1_3_6[0] <= majority_5041_port_o;
    roundReg_2_3_6[0] <= majority_5042_port_o;
    roundReg_3_3_6[0] <= majority_5043_port_o;
    roundReg_4_3_6[0] <= majority_5044_port_o;
    roundReg_5_3_6[0] <= majority_5045_port_o;
    roundReg_6_3_6[0] <= majority_5046_port_o;
    roundReg_7_3_6[0] <= majority_5047_port_o;
    roundReg_8_3_6[0] <= majority_5048_port_o;
    roundReg_9_3_6[0] <= majority_5049_port_o;
    roundReg_10_3_6[0] <= majority_5050_port_o;
    roundReg_11_3_6[0] <= majority_5051_port_o;
    roundReg_12_3_6[0] <= majority_5052_port_o;
    roundReg_13_3_6[0] <= majority_5053_port_o;
    roundReg_14_3_6[0] <= majority_5054_port_o;
    roundReg_15_3_6[0] <= majority_5055_port_o;
    roundReg_0_0_7[0] <= majority_5056_port_o;
    roundReg_1_0_7[0] <= majority_5057_port_o;
    roundReg_2_0_7[0] <= majority_5058_port_o;
    roundReg_3_0_7[0] <= majority_5059_port_o;
    roundReg_4_0_7[0] <= majority_5060_port_o;
    roundReg_5_0_7[0] <= majority_5061_port_o;
    roundReg_6_0_7[0] <= majority_5062_port_o;
    roundReg_7_0_7[0] <= majority_5063_port_o;
    roundReg_8_0_7[0] <= majority_5064_port_o;
    roundReg_9_0_7[0] <= majority_5065_port_o;
    roundReg_10_0_7[0] <= majority_5066_port_o;
    roundReg_11_0_7[0] <= majority_5067_port_o;
    roundReg_12_0_7[0] <= majority_5068_port_o;
    roundReg_13_0_7[0] <= majority_5069_port_o;
    roundReg_14_0_7[0] <= majority_5070_port_o;
    roundReg_15_0_7[0] <= majority_5071_port_o;
    roundReg_0_1_7[0] <= majority_5072_port_o;
    roundReg_1_1_7[0] <= majority_5073_port_o;
    roundReg_2_1_7[0] <= majority_5074_port_o;
    roundReg_3_1_7[0] <= majority_5075_port_o;
    roundReg_4_1_7[0] <= majority_5076_port_o;
    roundReg_5_1_7[0] <= majority_5077_port_o;
    roundReg_6_1_7[0] <= majority_5078_port_o;
    roundReg_7_1_7[0] <= majority_5079_port_o;
    roundReg_8_1_7[0] <= majority_5080_port_o;
    roundReg_9_1_7[0] <= majority_5081_port_o;
    roundReg_10_1_7[0] <= majority_5082_port_o;
    roundReg_11_1_7[0] <= majority_5083_port_o;
    roundReg_12_1_7[0] <= majority_5084_port_o;
    roundReg_13_1_7[0] <= majority_5085_port_o;
    roundReg_14_1_7[0] <= majority_5086_port_o;
    roundReg_15_1_7[0] <= majority_5087_port_o;
    roundReg_0_2_7[0] <= majority_5088_port_o;
    roundReg_1_2_7[0] <= majority_5089_port_o;
    roundReg_2_2_7[0] <= majority_5090_port_o;
    roundReg_3_2_7[0] <= majority_5091_port_o;
    roundReg_4_2_7[0] <= majority_5092_port_o;
    roundReg_5_2_7[0] <= majority_5093_port_o;
    roundReg_6_2_7[0] <= majority_5094_port_o;
    roundReg_7_2_7[0] <= majority_5095_port_o;
    roundReg_8_2_7[0] <= majority_5096_port_o;
    roundReg_9_2_7[0] <= majority_5097_port_o;
    roundReg_10_2_7[0] <= majority_5098_port_o;
    roundReg_11_2_7[0] <= majority_5099_port_o;
    roundReg_12_2_7[0] <= majority_5100_port_o;
    roundReg_13_2_7[0] <= majority_5101_port_o;
    roundReg_14_2_7[0] <= majority_5102_port_o;
    roundReg_15_2_7[0] <= majority_5103_port_o;
    roundReg_0_3_7[0] <= majority_5104_port_o;
    roundReg_1_3_7[0] <= majority_5105_port_o;
    roundReg_2_3_7[0] <= majority_5106_port_o;
    roundReg_3_3_7[0] <= majority_5107_port_o;
    roundReg_4_3_7[0] <= majority_5108_port_o;
    roundReg_5_3_7[0] <= majority_5109_port_o;
    roundReg_6_3_7[0] <= majority_5110_port_o;
    roundReg_7_3_7[0] <= majority_5111_port_o;
    roundReg_8_3_7[0] <= majority_5112_port_o;
    roundReg_9_3_7[0] <= majority_5113_port_o;
    roundReg_10_3_7[0] <= majority_5114_port_o;
    roundReg_11_3_7[0] <= majority_5115_port_o;
    roundReg_12_3_7[0] <= majority_5116_port_o;
    roundReg_13_3_7[0] <= majority_5117_port_o;
    roundReg_14_3_7[0] <= majority_5118_port_o;
    roundReg_15_3_7[0] <= majority_5119_port_o;
    roundReg_0_0_0[1] <= majority_5120_port_o;
    roundReg_1_0_0[1] <= majority_5121_port_o;
    roundReg_2_0_0[1] <= majority_5122_port_o;
    roundReg_3_0_0[1] <= majority_5123_port_o;
    roundReg_4_0_0[1] <= majority_5124_port_o;
    roundReg_5_0_0[1] <= majority_5125_port_o;
    roundReg_6_0_0[1] <= majority_5126_port_o;
    roundReg_7_0_0[1] <= majority_5127_port_o;
    roundReg_8_0_0[1] <= majority_5128_port_o;
    roundReg_9_0_0[1] <= majority_5129_port_o;
    roundReg_10_0_0[1] <= majority_5130_port_o;
    roundReg_11_0_0[1] <= majority_5131_port_o;
    roundReg_12_0_0[1] <= majority_5132_port_o;
    roundReg_13_0_0[1] <= majority_5133_port_o;
    roundReg_14_0_0[1] <= majority_5134_port_o;
    roundReg_15_0_0[1] <= majority_5135_port_o;
    roundReg_0_1_0[1] <= majority_5136_port_o;
    roundReg_1_1_0[1] <= majority_5137_port_o;
    roundReg_2_1_0[1] <= majority_5138_port_o;
    roundReg_3_1_0[1] <= majority_5139_port_o;
    roundReg_4_1_0[1] <= majority_5140_port_o;
    roundReg_5_1_0[1] <= majority_5141_port_o;
    roundReg_6_1_0[1] <= majority_5142_port_o;
    roundReg_7_1_0[1] <= majority_5143_port_o;
    roundReg_8_1_0[1] <= majority_5144_port_o;
    roundReg_9_1_0[1] <= majority_5145_port_o;
    roundReg_10_1_0[1] <= majority_5146_port_o;
    roundReg_11_1_0[1] <= majority_5147_port_o;
    roundReg_12_1_0[1] <= majority_5148_port_o;
    roundReg_13_1_0[1] <= majority_5149_port_o;
    roundReg_14_1_0[1] <= majority_5150_port_o;
    roundReg_15_1_0[1] <= majority_5151_port_o;
    roundReg_0_2_0[1] <= majority_5152_port_o;
    roundReg_1_2_0[1] <= majority_5153_port_o;
    roundReg_2_2_0[1] <= majority_5154_port_o;
    roundReg_3_2_0[1] <= majority_5155_port_o;
    roundReg_4_2_0[1] <= majority_5156_port_o;
    roundReg_5_2_0[1] <= majority_5157_port_o;
    roundReg_6_2_0[1] <= majority_5158_port_o;
    roundReg_7_2_0[1] <= majority_5159_port_o;
    roundReg_8_2_0[1] <= majority_5160_port_o;
    roundReg_9_2_0[1] <= majority_5161_port_o;
    roundReg_10_2_0[1] <= majority_5162_port_o;
    roundReg_11_2_0[1] <= majority_5163_port_o;
    roundReg_12_2_0[1] <= majority_5164_port_o;
    roundReg_13_2_0[1] <= majority_5165_port_o;
    roundReg_14_2_0[1] <= majority_5166_port_o;
    roundReg_15_2_0[1] <= majority_5167_port_o;
    roundReg_0_3_0[1] <= majority_5168_port_o;
    roundReg_1_3_0[1] <= majority_5169_port_o;
    roundReg_2_3_0[1] <= majority_5170_port_o;
    roundReg_3_3_0[1] <= majority_5171_port_o;
    roundReg_4_3_0[1] <= majority_5172_port_o;
    roundReg_5_3_0[1] <= majority_5173_port_o;
    roundReg_6_3_0[1] <= majority_5174_port_o;
    roundReg_7_3_0[1] <= majority_5175_port_o;
    roundReg_8_3_0[1] <= majority_5176_port_o;
    roundReg_9_3_0[1] <= majority_5177_port_o;
    roundReg_10_3_0[1] <= majority_5178_port_o;
    roundReg_11_3_0[1] <= majority_5179_port_o;
    roundReg_12_3_0[1] <= majority_5180_port_o;
    roundReg_13_3_0[1] <= majority_5181_port_o;
    roundReg_14_3_0[1] <= majority_5182_port_o;
    roundReg_15_3_0[1] <= majority_5183_port_o;
    roundReg_0_0_1[1] <= majority_5184_port_o;
    roundReg_1_0_1[1] <= majority_5185_port_o;
    roundReg_2_0_1[1] <= majority_5186_port_o;
    roundReg_3_0_1[1] <= majority_5187_port_o;
    roundReg_4_0_1[1] <= majority_5188_port_o;
    roundReg_5_0_1[1] <= majority_5189_port_o;
    roundReg_6_0_1[1] <= majority_5190_port_o;
    roundReg_7_0_1[1] <= majority_5191_port_o;
    roundReg_8_0_1[1] <= majority_5192_port_o;
    roundReg_9_0_1[1] <= majority_5193_port_o;
    roundReg_10_0_1[1] <= majority_5194_port_o;
    roundReg_11_0_1[1] <= majority_5195_port_o;
    roundReg_12_0_1[1] <= majority_5196_port_o;
    roundReg_13_0_1[1] <= majority_5197_port_o;
    roundReg_14_0_1[1] <= majority_5198_port_o;
    roundReg_15_0_1[1] <= majority_5199_port_o;
    roundReg_0_1_1[1] <= majority_5200_port_o;
    roundReg_1_1_1[1] <= majority_5201_port_o;
    roundReg_2_1_1[1] <= majority_5202_port_o;
    roundReg_3_1_1[1] <= majority_5203_port_o;
    roundReg_4_1_1[1] <= majority_5204_port_o;
    roundReg_5_1_1[1] <= majority_5205_port_o;
    roundReg_6_1_1[1] <= majority_5206_port_o;
    roundReg_7_1_1[1] <= majority_5207_port_o;
    roundReg_8_1_1[1] <= majority_5208_port_o;
    roundReg_9_1_1[1] <= majority_5209_port_o;
    roundReg_10_1_1[1] <= majority_5210_port_o;
    roundReg_11_1_1[1] <= majority_5211_port_o;
    roundReg_12_1_1[1] <= majority_5212_port_o;
    roundReg_13_1_1[1] <= majority_5213_port_o;
    roundReg_14_1_1[1] <= majority_5214_port_o;
    roundReg_15_1_1[1] <= majority_5215_port_o;
    roundReg_0_2_1[1] <= majority_5216_port_o;
    roundReg_1_2_1[1] <= majority_5217_port_o;
    roundReg_2_2_1[1] <= majority_5218_port_o;
    roundReg_3_2_1[1] <= majority_5219_port_o;
    roundReg_4_2_1[1] <= majority_5220_port_o;
    roundReg_5_2_1[1] <= majority_5221_port_o;
    roundReg_6_2_1[1] <= majority_5222_port_o;
    roundReg_7_2_1[1] <= majority_5223_port_o;
    roundReg_8_2_1[1] <= majority_5224_port_o;
    roundReg_9_2_1[1] <= majority_5225_port_o;
    roundReg_10_2_1[1] <= majority_5226_port_o;
    roundReg_11_2_1[1] <= majority_5227_port_o;
    roundReg_12_2_1[1] <= majority_5228_port_o;
    roundReg_13_2_1[1] <= majority_5229_port_o;
    roundReg_14_2_1[1] <= majority_5230_port_o;
    roundReg_15_2_1[1] <= majority_5231_port_o;
    roundReg_0_3_1[1] <= majority_5232_port_o;
    roundReg_1_3_1[1] <= majority_5233_port_o;
    roundReg_2_3_1[1] <= majority_5234_port_o;
    roundReg_3_3_1[1] <= majority_5235_port_o;
    roundReg_4_3_1[1] <= majority_5236_port_o;
    roundReg_5_3_1[1] <= majority_5237_port_o;
    roundReg_6_3_1[1] <= majority_5238_port_o;
    roundReg_7_3_1[1] <= majority_5239_port_o;
    roundReg_8_3_1[1] <= majority_5240_port_o;
    roundReg_9_3_1[1] <= majority_5241_port_o;
    roundReg_10_3_1[1] <= majority_5242_port_o;
    roundReg_11_3_1[1] <= majority_5243_port_o;
    roundReg_12_3_1[1] <= majority_5244_port_o;
    roundReg_13_3_1[1] <= majority_5245_port_o;
    roundReg_14_3_1[1] <= majority_5246_port_o;
    roundReg_15_3_1[1] <= majority_5247_port_o;
    roundReg_0_0_2[1] <= majority_5248_port_o;
    roundReg_1_0_2[1] <= majority_5249_port_o;
    roundReg_2_0_2[1] <= majority_5250_port_o;
    roundReg_3_0_2[1] <= majority_5251_port_o;
    roundReg_4_0_2[1] <= majority_5252_port_o;
    roundReg_5_0_2[1] <= majority_5253_port_o;
    roundReg_6_0_2[1] <= majority_5254_port_o;
    roundReg_7_0_2[1] <= majority_5255_port_o;
    roundReg_8_0_2[1] <= majority_5256_port_o;
    roundReg_9_0_2[1] <= majority_5257_port_o;
    roundReg_10_0_2[1] <= majority_5258_port_o;
    roundReg_11_0_2[1] <= majority_5259_port_o;
    roundReg_12_0_2[1] <= majority_5260_port_o;
    roundReg_13_0_2[1] <= majority_5261_port_o;
    roundReg_14_0_2[1] <= majority_5262_port_o;
    roundReg_15_0_2[1] <= majority_5263_port_o;
    roundReg_0_1_2[1] <= majority_5264_port_o;
    roundReg_1_1_2[1] <= majority_5265_port_o;
    roundReg_2_1_2[1] <= majority_5266_port_o;
    roundReg_3_1_2[1] <= majority_5267_port_o;
    roundReg_4_1_2[1] <= majority_5268_port_o;
    roundReg_5_1_2[1] <= majority_5269_port_o;
    roundReg_6_1_2[1] <= majority_5270_port_o;
    roundReg_7_1_2[1] <= majority_5271_port_o;
    roundReg_8_1_2[1] <= majority_5272_port_o;
    roundReg_9_1_2[1] <= majority_5273_port_o;
    roundReg_10_1_2[1] <= majority_5274_port_o;
    roundReg_11_1_2[1] <= majority_5275_port_o;
    roundReg_12_1_2[1] <= majority_5276_port_o;
    roundReg_13_1_2[1] <= majority_5277_port_o;
    roundReg_14_1_2[1] <= majority_5278_port_o;
    roundReg_15_1_2[1] <= majority_5279_port_o;
    roundReg_0_2_2[1] <= majority_5280_port_o;
    roundReg_1_2_2[1] <= majority_5281_port_o;
    roundReg_2_2_2[1] <= majority_5282_port_o;
    roundReg_3_2_2[1] <= majority_5283_port_o;
    roundReg_4_2_2[1] <= majority_5284_port_o;
    roundReg_5_2_2[1] <= majority_5285_port_o;
    roundReg_6_2_2[1] <= majority_5286_port_o;
    roundReg_7_2_2[1] <= majority_5287_port_o;
    roundReg_8_2_2[1] <= majority_5288_port_o;
    roundReg_9_2_2[1] <= majority_5289_port_o;
    roundReg_10_2_2[1] <= majority_5290_port_o;
    roundReg_11_2_2[1] <= majority_5291_port_o;
    roundReg_12_2_2[1] <= majority_5292_port_o;
    roundReg_13_2_2[1] <= majority_5293_port_o;
    roundReg_14_2_2[1] <= majority_5294_port_o;
    roundReg_15_2_2[1] <= majority_5295_port_o;
    roundReg_0_3_2[1] <= majority_5296_port_o;
    roundReg_1_3_2[1] <= majority_5297_port_o;
    roundReg_2_3_2[1] <= majority_5298_port_o;
    roundReg_3_3_2[1] <= majority_5299_port_o;
    roundReg_4_3_2[1] <= majority_5300_port_o;
    roundReg_5_3_2[1] <= majority_5301_port_o;
    roundReg_6_3_2[1] <= majority_5302_port_o;
    roundReg_7_3_2[1] <= majority_5303_port_o;
    roundReg_8_3_2[1] <= majority_5304_port_o;
    roundReg_9_3_2[1] <= majority_5305_port_o;
    roundReg_10_3_2[1] <= majority_5306_port_o;
    roundReg_11_3_2[1] <= majority_5307_port_o;
    roundReg_12_3_2[1] <= majority_5308_port_o;
    roundReg_13_3_2[1] <= majority_5309_port_o;
    roundReg_14_3_2[1] <= majority_5310_port_o;
    roundReg_15_3_2[1] <= majority_5311_port_o;
    roundReg_0_0_3[1] <= majority_5312_port_o;
    roundReg_1_0_3[1] <= majority_5313_port_o;
    roundReg_2_0_3[1] <= majority_5314_port_o;
    roundReg_3_0_3[1] <= majority_5315_port_o;
    roundReg_4_0_3[1] <= majority_5316_port_o;
    roundReg_5_0_3[1] <= majority_5317_port_o;
    roundReg_6_0_3[1] <= majority_5318_port_o;
    roundReg_7_0_3[1] <= majority_5319_port_o;
    roundReg_8_0_3[1] <= majority_5320_port_o;
    roundReg_9_0_3[1] <= majority_5321_port_o;
    roundReg_10_0_3[1] <= majority_5322_port_o;
    roundReg_11_0_3[1] <= majority_5323_port_o;
    roundReg_12_0_3[1] <= majority_5324_port_o;
    roundReg_13_0_3[1] <= majority_5325_port_o;
    roundReg_14_0_3[1] <= majority_5326_port_o;
    roundReg_15_0_3[1] <= majority_5327_port_o;
    roundReg_0_1_3[1] <= majority_5328_port_o;
    roundReg_1_1_3[1] <= majority_5329_port_o;
    roundReg_2_1_3[1] <= majority_5330_port_o;
    roundReg_3_1_3[1] <= majority_5331_port_o;
    roundReg_4_1_3[1] <= majority_5332_port_o;
    roundReg_5_1_3[1] <= majority_5333_port_o;
    roundReg_6_1_3[1] <= majority_5334_port_o;
    roundReg_7_1_3[1] <= majority_5335_port_o;
    roundReg_8_1_3[1] <= majority_5336_port_o;
    roundReg_9_1_3[1] <= majority_5337_port_o;
    roundReg_10_1_3[1] <= majority_5338_port_o;
    roundReg_11_1_3[1] <= majority_5339_port_o;
    roundReg_12_1_3[1] <= majority_5340_port_o;
    roundReg_13_1_3[1] <= majority_5341_port_o;
    roundReg_14_1_3[1] <= majority_5342_port_o;
    roundReg_15_1_3[1] <= majority_5343_port_o;
    roundReg_0_2_3[1] <= majority_5344_port_o;
    roundReg_1_2_3[1] <= majority_5345_port_o;
    roundReg_2_2_3[1] <= majority_5346_port_o;
    roundReg_3_2_3[1] <= majority_5347_port_o;
    roundReg_4_2_3[1] <= majority_5348_port_o;
    roundReg_5_2_3[1] <= majority_5349_port_o;
    roundReg_6_2_3[1] <= majority_5350_port_o;
    roundReg_7_2_3[1] <= majority_5351_port_o;
    roundReg_8_2_3[1] <= majority_5352_port_o;
    roundReg_9_2_3[1] <= majority_5353_port_o;
    roundReg_10_2_3[1] <= majority_5354_port_o;
    roundReg_11_2_3[1] <= majority_5355_port_o;
    roundReg_12_2_3[1] <= majority_5356_port_o;
    roundReg_13_2_3[1] <= majority_5357_port_o;
    roundReg_14_2_3[1] <= majority_5358_port_o;
    roundReg_15_2_3[1] <= majority_5359_port_o;
    roundReg_0_3_3[1] <= majority_5360_port_o;
    roundReg_1_3_3[1] <= majority_5361_port_o;
    roundReg_2_3_3[1] <= majority_5362_port_o;
    roundReg_3_3_3[1] <= majority_5363_port_o;
    roundReg_4_3_3[1] <= majority_5364_port_o;
    roundReg_5_3_3[1] <= majority_5365_port_o;
    roundReg_6_3_3[1] <= majority_5366_port_o;
    roundReg_7_3_3[1] <= majority_5367_port_o;
    roundReg_8_3_3[1] <= majority_5368_port_o;
    roundReg_9_3_3[1] <= majority_5369_port_o;
    roundReg_10_3_3[1] <= majority_5370_port_o;
    roundReg_11_3_3[1] <= majority_5371_port_o;
    roundReg_12_3_3[1] <= majority_5372_port_o;
    roundReg_13_3_3[1] <= majority_5373_port_o;
    roundReg_14_3_3[1] <= majority_5374_port_o;
    roundReg_15_3_3[1] <= majority_5375_port_o;
    roundReg_0_0_4[1] <= majority_5376_port_o;
    roundReg_1_0_4[1] <= majority_5377_port_o;
    roundReg_2_0_4[1] <= majority_5378_port_o;
    roundReg_3_0_4[1] <= majority_5379_port_o;
    roundReg_4_0_4[1] <= majority_5380_port_o;
    roundReg_5_0_4[1] <= majority_5381_port_o;
    roundReg_6_0_4[1] <= majority_5382_port_o;
    roundReg_7_0_4[1] <= majority_5383_port_o;
    roundReg_8_0_4[1] <= majority_5384_port_o;
    roundReg_9_0_4[1] <= majority_5385_port_o;
    roundReg_10_0_4[1] <= majority_5386_port_o;
    roundReg_11_0_4[1] <= majority_5387_port_o;
    roundReg_12_0_4[1] <= majority_5388_port_o;
    roundReg_13_0_4[1] <= majority_5389_port_o;
    roundReg_14_0_4[1] <= majority_5390_port_o;
    roundReg_15_0_4[1] <= majority_5391_port_o;
    roundReg_0_1_4[1] <= majority_5392_port_o;
    roundReg_1_1_4[1] <= majority_5393_port_o;
    roundReg_2_1_4[1] <= majority_5394_port_o;
    roundReg_3_1_4[1] <= majority_5395_port_o;
    roundReg_4_1_4[1] <= majority_5396_port_o;
    roundReg_5_1_4[1] <= majority_5397_port_o;
    roundReg_6_1_4[1] <= majority_5398_port_o;
    roundReg_7_1_4[1] <= majority_5399_port_o;
    roundReg_8_1_4[1] <= majority_5400_port_o;
    roundReg_9_1_4[1] <= majority_5401_port_o;
    roundReg_10_1_4[1] <= majority_5402_port_o;
    roundReg_11_1_4[1] <= majority_5403_port_o;
    roundReg_12_1_4[1] <= majority_5404_port_o;
    roundReg_13_1_4[1] <= majority_5405_port_o;
    roundReg_14_1_4[1] <= majority_5406_port_o;
    roundReg_15_1_4[1] <= majority_5407_port_o;
    roundReg_0_2_4[1] <= majority_5408_port_o;
    roundReg_1_2_4[1] <= majority_5409_port_o;
    roundReg_2_2_4[1] <= majority_5410_port_o;
    roundReg_3_2_4[1] <= majority_5411_port_o;
    roundReg_4_2_4[1] <= majority_5412_port_o;
    roundReg_5_2_4[1] <= majority_5413_port_o;
    roundReg_6_2_4[1] <= majority_5414_port_o;
    roundReg_7_2_4[1] <= majority_5415_port_o;
    roundReg_8_2_4[1] <= majority_5416_port_o;
    roundReg_9_2_4[1] <= majority_5417_port_o;
    roundReg_10_2_4[1] <= majority_5418_port_o;
    roundReg_11_2_4[1] <= majority_5419_port_o;
    roundReg_12_2_4[1] <= majority_5420_port_o;
    roundReg_13_2_4[1] <= majority_5421_port_o;
    roundReg_14_2_4[1] <= majority_5422_port_o;
    roundReg_15_2_4[1] <= majority_5423_port_o;
    roundReg_0_3_4[1] <= majority_5424_port_o;
    roundReg_1_3_4[1] <= majority_5425_port_o;
    roundReg_2_3_4[1] <= majority_5426_port_o;
    roundReg_3_3_4[1] <= majority_5427_port_o;
    roundReg_4_3_4[1] <= majority_5428_port_o;
    roundReg_5_3_4[1] <= majority_5429_port_o;
    roundReg_6_3_4[1] <= majority_5430_port_o;
    roundReg_7_3_4[1] <= majority_5431_port_o;
    roundReg_8_3_4[1] <= majority_5432_port_o;
    roundReg_9_3_4[1] <= majority_5433_port_o;
    roundReg_10_3_4[1] <= majority_5434_port_o;
    roundReg_11_3_4[1] <= majority_5435_port_o;
    roundReg_12_3_4[1] <= majority_5436_port_o;
    roundReg_13_3_4[1] <= majority_5437_port_o;
    roundReg_14_3_4[1] <= majority_5438_port_o;
    roundReg_15_3_4[1] <= majority_5439_port_o;
    roundReg_0_0_5[1] <= majority_5440_port_o;
    roundReg_1_0_5[1] <= majority_5441_port_o;
    roundReg_2_0_5[1] <= majority_5442_port_o;
    roundReg_3_0_5[1] <= majority_5443_port_o;
    roundReg_4_0_5[1] <= majority_5444_port_o;
    roundReg_5_0_5[1] <= majority_5445_port_o;
    roundReg_6_0_5[1] <= majority_5446_port_o;
    roundReg_7_0_5[1] <= majority_5447_port_o;
    roundReg_8_0_5[1] <= majority_5448_port_o;
    roundReg_9_0_5[1] <= majority_5449_port_o;
    roundReg_10_0_5[1] <= majority_5450_port_o;
    roundReg_11_0_5[1] <= majority_5451_port_o;
    roundReg_12_0_5[1] <= majority_5452_port_o;
    roundReg_13_0_5[1] <= majority_5453_port_o;
    roundReg_14_0_5[1] <= majority_5454_port_o;
    roundReg_15_0_5[1] <= majority_5455_port_o;
    roundReg_0_1_5[1] <= majority_5456_port_o;
    roundReg_1_1_5[1] <= majority_5457_port_o;
    roundReg_2_1_5[1] <= majority_5458_port_o;
    roundReg_3_1_5[1] <= majority_5459_port_o;
    roundReg_4_1_5[1] <= majority_5460_port_o;
    roundReg_5_1_5[1] <= majority_5461_port_o;
    roundReg_6_1_5[1] <= majority_5462_port_o;
    roundReg_7_1_5[1] <= majority_5463_port_o;
    roundReg_8_1_5[1] <= majority_5464_port_o;
    roundReg_9_1_5[1] <= majority_5465_port_o;
    roundReg_10_1_5[1] <= majority_5466_port_o;
    roundReg_11_1_5[1] <= majority_5467_port_o;
    roundReg_12_1_5[1] <= majority_5468_port_o;
    roundReg_13_1_5[1] <= majority_5469_port_o;
    roundReg_14_1_5[1] <= majority_5470_port_o;
    roundReg_15_1_5[1] <= majority_5471_port_o;
    roundReg_0_2_5[1] <= majority_5472_port_o;
    roundReg_1_2_5[1] <= majority_5473_port_o;
    roundReg_2_2_5[1] <= majority_5474_port_o;
    roundReg_3_2_5[1] <= majority_5475_port_o;
    roundReg_4_2_5[1] <= majority_5476_port_o;
    roundReg_5_2_5[1] <= majority_5477_port_o;
    roundReg_6_2_5[1] <= majority_5478_port_o;
    roundReg_7_2_5[1] <= majority_5479_port_o;
    roundReg_8_2_5[1] <= majority_5480_port_o;
    roundReg_9_2_5[1] <= majority_5481_port_o;
    roundReg_10_2_5[1] <= majority_5482_port_o;
    roundReg_11_2_5[1] <= majority_5483_port_o;
    roundReg_12_2_5[1] <= majority_5484_port_o;
    roundReg_13_2_5[1] <= majority_5485_port_o;
    roundReg_14_2_5[1] <= majority_5486_port_o;
    roundReg_15_2_5[1] <= majority_5487_port_o;
    roundReg_0_3_5[1] <= majority_5488_port_o;
    roundReg_1_3_5[1] <= majority_5489_port_o;
    roundReg_2_3_5[1] <= majority_5490_port_o;
    roundReg_3_3_5[1] <= majority_5491_port_o;
    roundReg_4_3_5[1] <= majority_5492_port_o;
    roundReg_5_3_5[1] <= majority_5493_port_o;
    roundReg_6_3_5[1] <= majority_5494_port_o;
    roundReg_7_3_5[1] <= majority_5495_port_o;
    roundReg_8_3_5[1] <= majority_5496_port_o;
    roundReg_9_3_5[1] <= majority_5497_port_o;
    roundReg_10_3_5[1] <= majority_5498_port_o;
    roundReg_11_3_5[1] <= majority_5499_port_o;
    roundReg_12_3_5[1] <= majority_5500_port_o;
    roundReg_13_3_5[1] <= majority_5501_port_o;
    roundReg_14_3_5[1] <= majority_5502_port_o;
    roundReg_15_3_5[1] <= majority_5503_port_o;
    roundReg_0_0_6[1] <= majority_5504_port_o;
    roundReg_1_0_6[1] <= majority_5505_port_o;
    roundReg_2_0_6[1] <= majority_5506_port_o;
    roundReg_3_0_6[1] <= majority_5507_port_o;
    roundReg_4_0_6[1] <= majority_5508_port_o;
    roundReg_5_0_6[1] <= majority_5509_port_o;
    roundReg_6_0_6[1] <= majority_5510_port_o;
    roundReg_7_0_6[1] <= majority_5511_port_o;
    roundReg_8_0_6[1] <= majority_5512_port_o;
    roundReg_9_0_6[1] <= majority_5513_port_o;
    roundReg_10_0_6[1] <= majority_5514_port_o;
    roundReg_11_0_6[1] <= majority_5515_port_o;
    roundReg_12_0_6[1] <= majority_5516_port_o;
    roundReg_13_0_6[1] <= majority_5517_port_o;
    roundReg_14_0_6[1] <= majority_5518_port_o;
    roundReg_15_0_6[1] <= majority_5519_port_o;
    roundReg_0_1_6[1] <= majority_5520_port_o;
    roundReg_1_1_6[1] <= majority_5521_port_o;
    roundReg_2_1_6[1] <= majority_5522_port_o;
    roundReg_3_1_6[1] <= majority_5523_port_o;
    roundReg_4_1_6[1] <= majority_5524_port_o;
    roundReg_5_1_6[1] <= majority_5525_port_o;
    roundReg_6_1_6[1] <= majority_5526_port_o;
    roundReg_7_1_6[1] <= majority_5527_port_o;
    roundReg_8_1_6[1] <= majority_5528_port_o;
    roundReg_9_1_6[1] <= majority_5529_port_o;
    roundReg_10_1_6[1] <= majority_5530_port_o;
    roundReg_11_1_6[1] <= majority_5531_port_o;
    roundReg_12_1_6[1] <= majority_5532_port_o;
    roundReg_13_1_6[1] <= majority_5533_port_o;
    roundReg_14_1_6[1] <= majority_5534_port_o;
    roundReg_15_1_6[1] <= majority_5535_port_o;
    roundReg_0_2_6[1] <= majority_5536_port_o;
    roundReg_1_2_6[1] <= majority_5537_port_o;
    roundReg_2_2_6[1] <= majority_5538_port_o;
    roundReg_3_2_6[1] <= majority_5539_port_o;
    roundReg_4_2_6[1] <= majority_5540_port_o;
    roundReg_5_2_6[1] <= majority_5541_port_o;
    roundReg_6_2_6[1] <= majority_5542_port_o;
    roundReg_7_2_6[1] <= majority_5543_port_o;
    roundReg_8_2_6[1] <= majority_5544_port_o;
    roundReg_9_2_6[1] <= majority_5545_port_o;
    roundReg_10_2_6[1] <= majority_5546_port_o;
    roundReg_11_2_6[1] <= majority_5547_port_o;
    roundReg_12_2_6[1] <= majority_5548_port_o;
    roundReg_13_2_6[1] <= majority_5549_port_o;
    roundReg_14_2_6[1] <= majority_5550_port_o;
    roundReg_15_2_6[1] <= majority_5551_port_o;
    roundReg_0_3_6[1] <= majority_5552_port_o;
    roundReg_1_3_6[1] <= majority_5553_port_o;
    roundReg_2_3_6[1] <= majority_5554_port_o;
    roundReg_3_3_6[1] <= majority_5555_port_o;
    roundReg_4_3_6[1] <= majority_5556_port_o;
    roundReg_5_3_6[1] <= majority_5557_port_o;
    roundReg_6_3_6[1] <= majority_5558_port_o;
    roundReg_7_3_6[1] <= majority_5559_port_o;
    roundReg_8_3_6[1] <= majority_5560_port_o;
    roundReg_9_3_6[1] <= majority_5561_port_o;
    roundReg_10_3_6[1] <= majority_5562_port_o;
    roundReg_11_3_6[1] <= majority_5563_port_o;
    roundReg_12_3_6[1] <= majority_5564_port_o;
    roundReg_13_3_6[1] <= majority_5565_port_o;
    roundReg_14_3_6[1] <= majority_5566_port_o;
    roundReg_15_3_6[1] <= majority_5567_port_o;
    roundReg_0_0_7[1] <= majority_5568_port_o;
    roundReg_1_0_7[1] <= majority_5569_port_o;
    roundReg_2_0_7[1] <= majority_5570_port_o;
    roundReg_3_0_7[1] <= majority_5571_port_o;
    roundReg_4_0_7[1] <= majority_5572_port_o;
    roundReg_5_0_7[1] <= majority_5573_port_o;
    roundReg_6_0_7[1] <= majority_5574_port_o;
    roundReg_7_0_7[1] <= majority_5575_port_o;
    roundReg_8_0_7[1] <= majority_5576_port_o;
    roundReg_9_0_7[1] <= majority_5577_port_o;
    roundReg_10_0_7[1] <= majority_5578_port_o;
    roundReg_11_0_7[1] <= majority_5579_port_o;
    roundReg_12_0_7[1] <= majority_5580_port_o;
    roundReg_13_0_7[1] <= majority_5581_port_o;
    roundReg_14_0_7[1] <= majority_5582_port_o;
    roundReg_15_0_7[1] <= majority_5583_port_o;
    roundReg_0_1_7[1] <= majority_5584_port_o;
    roundReg_1_1_7[1] <= majority_5585_port_o;
    roundReg_2_1_7[1] <= majority_5586_port_o;
    roundReg_3_1_7[1] <= majority_5587_port_o;
    roundReg_4_1_7[1] <= majority_5588_port_o;
    roundReg_5_1_7[1] <= majority_5589_port_o;
    roundReg_6_1_7[1] <= majority_5590_port_o;
    roundReg_7_1_7[1] <= majority_5591_port_o;
    roundReg_8_1_7[1] <= majority_5592_port_o;
    roundReg_9_1_7[1] <= majority_5593_port_o;
    roundReg_10_1_7[1] <= majority_5594_port_o;
    roundReg_11_1_7[1] <= majority_5595_port_o;
    roundReg_12_1_7[1] <= majority_5596_port_o;
    roundReg_13_1_7[1] <= majority_5597_port_o;
    roundReg_14_1_7[1] <= majority_5598_port_o;
    roundReg_15_1_7[1] <= majority_5599_port_o;
    roundReg_0_2_7[1] <= majority_5600_port_o;
    roundReg_1_2_7[1] <= majority_5601_port_o;
    roundReg_2_2_7[1] <= majority_5602_port_o;
    roundReg_3_2_7[1] <= majority_5603_port_o;
    roundReg_4_2_7[1] <= majority_5604_port_o;
    roundReg_5_2_7[1] <= majority_5605_port_o;
    roundReg_6_2_7[1] <= majority_5606_port_o;
    roundReg_7_2_7[1] <= majority_5607_port_o;
    roundReg_8_2_7[1] <= majority_5608_port_o;
    roundReg_9_2_7[1] <= majority_5609_port_o;
    roundReg_10_2_7[1] <= majority_5610_port_o;
    roundReg_11_2_7[1] <= majority_5611_port_o;
    roundReg_12_2_7[1] <= majority_5612_port_o;
    roundReg_13_2_7[1] <= majority_5613_port_o;
    roundReg_14_2_7[1] <= majority_5614_port_o;
    roundReg_15_2_7[1] <= majority_5615_port_o;
    roundReg_0_3_7[1] <= majority_5616_port_o;
    roundReg_1_3_7[1] <= majority_5617_port_o;
    roundReg_2_3_7[1] <= majority_5618_port_o;
    roundReg_3_3_7[1] <= majority_5619_port_o;
    roundReg_4_3_7[1] <= majority_5620_port_o;
    roundReg_5_3_7[1] <= majority_5621_port_o;
    roundReg_6_3_7[1] <= majority_5622_port_o;
    roundReg_7_3_7[1] <= majority_5623_port_o;
    roundReg_8_3_7[1] <= majority_5624_port_o;
    roundReg_9_3_7[1] <= majority_5625_port_o;
    roundReg_10_3_7[1] <= majority_5626_port_o;
    roundReg_11_3_7[1] <= majority_5627_port_o;
    roundReg_12_3_7[1] <= majority_5628_port_o;
    roundReg_13_3_7[1] <= majority_5629_port_o;
    roundReg_14_3_7[1] <= majority_5630_port_o;
    roundReg_15_3_7[1] <= majority_5631_port_o;
    roundReg_0_0_0[2] <= majority_5632_port_o;
    roundReg_1_0_0[2] <= majority_5633_port_o;
    roundReg_2_0_0[2] <= majority_5634_port_o;
    roundReg_3_0_0[2] <= majority_5635_port_o;
    roundReg_4_0_0[2] <= majority_5636_port_o;
    roundReg_5_0_0[2] <= majority_5637_port_o;
    roundReg_6_0_0[2] <= majority_5638_port_o;
    roundReg_7_0_0[2] <= majority_5639_port_o;
    roundReg_8_0_0[2] <= majority_5640_port_o;
    roundReg_9_0_0[2] <= majority_5641_port_o;
    roundReg_10_0_0[2] <= majority_5642_port_o;
    roundReg_11_0_0[2] <= majority_5643_port_o;
    roundReg_12_0_0[2] <= majority_5644_port_o;
    roundReg_13_0_0[2] <= majority_5645_port_o;
    roundReg_14_0_0[2] <= majority_5646_port_o;
    roundReg_15_0_0[2] <= majority_5647_port_o;
    roundReg_0_1_0[2] <= majority_5648_port_o;
    roundReg_1_1_0[2] <= majority_5649_port_o;
    roundReg_2_1_0[2] <= majority_5650_port_o;
    roundReg_3_1_0[2] <= majority_5651_port_o;
    roundReg_4_1_0[2] <= majority_5652_port_o;
    roundReg_5_1_0[2] <= majority_5653_port_o;
    roundReg_6_1_0[2] <= majority_5654_port_o;
    roundReg_7_1_0[2] <= majority_5655_port_o;
    roundReg_8_1_0[2] <= majority_5656_port_o;
    roundReg_9_1_0[2] <= majority_5657_port_o;
    roundReg_10_1_0[2] <= majority_5658_port_o;
    roundReg_11_1_0[2] <= majority_5659_port_o;
    roundReg_12_1_0[2] <= majority_5660_port_o;
    roundReg_13_1_0[2] <= majority_5661_port_o;
    roundReg_14_1_0[2] <= majority_5662_port_o;
    roundReg_15_1_0[2] <= majority_5663_port_o;
    roundReg_0_2_0[2] <= majority_5664_port_o;
    roundReg_1_2_0[2] <= majority_5665_port_o;
    roundReg_2_2_0[2] <= majority_5666_port_o;
    roundReg_3_2_0[2] <= majority_5667_port_o;
    roundReg_4_2_0[2] <= majority_5668_port_o;
    roundReg_5_2_0[2] <= majority_5669_port_o;
    roundReg_6_2_0[2] <= majority_5670_port_o;
    roundReg_7_2_0[2] <= majority_5671_port_o;
    roundReg_8_2_0[2] <= majority_5672_port_o;
    roundReg_9_2_0[2] <= majority_5673_port_o;
    roundReg_10_2_0[2] <= majority_5674_port_o;
    roundReg_11_2_0[2] <= majority_5675_port_o;
    roundReg_12_2_0[2] <= majority_5676_port_o;
    roundReg_13_2_0[2] <= majority_5677_port_o;
    roundReg_14_2_0[2] <= majority_5678_port_o;
    roundReg_15_2_0[2] <= majority_5679_port_o;
    roundReg_0_3_0[2] <= majority_5680_port_o;
    roundReg_1_3_0[2] <= majority_5681_port_o;
    roundReg_2_3_0[2] <= majority_5682_port_o;
    roundReg_3_3_0[2] <= majority_5683_port_o;
    roundReg_4_3_0[2] <= majority_5684_port_o;
    roundReg_5_3_0[2] <= majority_5685_port_o;
    roundReg_6_3_0[2] <= majority_5686_port_o;
    roundReg_7_3_0[2] <= majority_5687_port_o;
    roundReg_8_3_0[2] <= majority_5688_port_o;
    roundReg_9_3_0[2] <= majority_5689_port_o;
    roundReg_10_3_0[2] <= majority_5690_port_o;
    roundReg_11_3_0[2] <= majority_5691_port_o;
    roundReg_12_3_0[2] <= majority_5692_port_o;
    roundReg_13_3_0[2] <= majority_5693_port_o;
    roundReg_14_3_0[2] <= majority_5694_port_o;
    roundReg_15_3_0[2] <= majority_5695_port_o;
    roundReg_0_0_1[2] <= majority_5696_port_o;
    roundReg_1_0_1[2] <= majority_5697_port_o;
    roundReg_2_0_1[2] <= majority_5698_port_o;
    roundReg_3_0_1[2] <= majority_5699_port_o;
    roundReg_4_0_1[2] <= majority_5700_port_o;
    roundReg_5_0_1[2] <= majority_5701_port_o;
    roundReg_6_0_1[2] <= majority_5702_port_o;
    roundReg_7_0_1[2] <= majority_5703_port_o;
    roundReg_8_0_1[2] <= majority_5704_port_o;
    roundReg_9_0_1[2] <= majority_5705_port_o;
    roundReg_10_0_1[2] <= majority_5706_port_o;
    roundReg_11_0_1[2] <= majority_5707_port_o;
    roundReg_12_0_1[2] <= majority_5708_port_o;
    roundReg_13_0_1[2] <= majority_5709_port_o;
    roundReg_14_0_1[2] <= majority_5710_port_o;
    roundReg_15_0_1[2] <= majority_5711_port_o;
    roundReg_0_1_1[2] <= majority_5712_port_o;
    roundReg_1_1_1[2] <= majority_5713_port_o;
    roundReg_2_1_1[2] <= majority_5714_port_o;
    roundReg_3_1_1[2] <= majority_5715_port_o;
    roundReg_4_1_1[2] <= majority_5716_port_o;
    roundReg_5_1_1[2] <= majority_5717_port_o;
    roundReg_6_1_1[2] <= majority_5718_port_o;
    roundReg_7_1_1[2] <= majority_5719_port_o;
    roundReg_8_1_1[2] <= majority_5720_port_o;
    roundReg_9_1_1[2] <= majority_5721_port_o;
    roundReg_10_1_1[2] <= majority_5722_port_o;
    roundReg_11_1_1[2] <= majority_5723_port_o;
    roundReg_12_1_1[2] <= majority_5724_port_o;
    roundReg_13_1_1[2] <= majority_5725_port_o;
    roundReg_14_1_1[2] <= majority_5726_port_o;
    roundReg_15_1_1[2] <= majority_5727_port_o;
    roundReg_0_2_1[2] <= majority_5728_port_o;
    roundReg_1_2_1[2] <= majority_5729_port_o;
    roundReg_2_2_1[2] <= majority_5730_port_o;
    roundReg_3_2_1[2] <= majority_5731_port_o;
    roundReg_4_2_1[2] <= majority_5732_port_o;
    roundReg_5_2_1[2] <= majority_5733_port_o;
    roundReg_6_2_1[2] <= majority_5734_port_o;
    roundReg_7_2_1[2] <= majority_5735_port_o;
    roundReg_8_2_1[2] <= majority_5736_port_o;
    roundReg_9_2_1[2] <= majority_5737_port_o;
    roundReg_10_2_1[2] <= majority_5738_port_o;
    roundReg_11_2_1[2] <= majority_5739_port_o;
    roundReg_12_2_1[2] <= majority_5740_port_o;
    roundReg_13_2_1[2] <= majority_5741_port_o;
    roundReg_14_2_1[2] <= majority_5742_port_o;
    roundReg_15_2_1[2] <= majority_5743_port_o;
    roundReg_0_3_1[2] <= majority_5744_port_o;
    roundReg_1_3_1[2] <= majority_5745_port_o;
    roundReg_2_3_1[2] <= majority_5746_port_o;
    roundReg_3_3_1[2] <= majority_5747_port_o;
    roundReg_4_3_1[2] <= majority_5748_port_o;
    roundReg_5_3_1[2] <= majority_5749_port_o;
    roundReg_6_3_1[2] <= majority_5750_port_o;
    roundReg_7_3_1[2] <= majority_5751_port_o;
    roundReg_8_3_1[2] <= majority_5752_port_o;
    roundReg_9_3_1[2] <= majority_5753_port_o;
    roundReg_10_3_1[2] <= majority_5754_port_o;
    roundReg_11_3_1[2] <= majority_5755_port_o;
    roundReg_12_3_1[2] <= majority_5756_port_o;
    roundReg_13_3_1[2] <= majority_5757_port_o;
    roundReg_14_3_1[2] <= majority_5758_port_o;
    roundReg_15_3_1[2] <= majority_5759_port_o;
    roundReg_0_0_2[2] <= majority_5760_port_o;
    roundReg_1_0_2[2] <= majority_5761_port_o;
    roundReg_2_0_2[2] <= majority_5762_port_o;
    roundReg_3_0_2[2] <= majority_5763_port_o;
    roundReg_4_0_2[2] <= majority_5764_port_o;
    roundReg_5_0_2[2] <= majority_5765_port_o;
    roundReg_6_0_2[2] <= majority_5766_port_o;
    roundReg_7_0_2[2] <= majority_5767_port_o;
    roundReg_8_0_2[2] <= majority_5768_port_o;
    roundReg_9_0_2[2] <= majority_5769_port_o;
    roundReg_10_0_2[2] <= majority_5770_port_o;
    roundReg_11_0_2[2] <= majority_5771_port_o;
    roundReg_12_0_2[2] <= majority_5772_port_o;
    roundReg_13_0_2[2] <= majority_5773_port_o;
    roundReg_14_0_2[2] <= majority_5774_port_o;
    roundReg_15_0_2[2] <= majority_5775_port_o;
    roundReg_0_1_2[2] <= majority_5776_port_o;
    roundReg_1_1_2[2] <= majority_5777_port_o;
    roundReg_2_1_2[2] <= majority_5778_port_o;
    roundReg_3_1_2[2] <= majority_5779_port_o;
    roundReg_4_1_2[2] <= majority_5780_port_o;
    roundReg_5_1_2[2] <= majority_5781_port_o;
    roundReg_6_1_2[2] <= majority_5782_port_o;
    roundReg_7_1_2[2] <= majority_5783_port_o;
    roundReg_8_1_2[2] <= majority_5784_port_o;
    roundReg_9_1_2[2] <= majority_5785_port_o;
    roundReg_10_1_2[2] <= majority_5786_port_o;
    roundReg_11_1_2[2] <= majority_5787_port_o;
    roundReg_12_1_2[2] <= majority_5788_port_o;
    roundReg_13_1_2[2] <= majority_5789_port_o;
    roundReg_14_1_2[2] <= majority_5790_port_o;
    roundReg_15_1_2[2] <= majority_5791_port_o;
    roundReg_0_2_2[2] <= majority_5792_port_o;
    roundReg_1_2_2[2] <= majority_5793_port_o;
    roundReg_2_2_2[2] <= majority_5794_port_o;
    roundReg_3_2_2[2] <= majority_5795_port_o;
    roundReg_4_2_2[2] <= majority_5796_port_o;
    roundReg_5_2_2[2] <= majority_5797_port_o;
    roundReg_6_2_2[2] <= majority_5798_port_o;
    roundReg_7_2_2[2] <= majority_5799_port_o;
    roundReg_8_2_2[2] <= majority_5800_port_o;
    roundReg_9_2_2[2] <= majority_5801_port_o;
    roundReg_10_2_2[2] <= majority_5802_port_o;
    roundReg_11_2_2[2] <= majority_5803_port_o;
    roundReg_12_2_2[2] <= majority_5804_port_o;
    roundReg_13_2_2[2] <= majority_5805_port_o;
    roundReg_14_2_2[2] <= majority_5806_port_o;
    roundReg_15_2_2[2] <= majority_5807_port_o;
    roundReg_0_3_2[2] <= majority_5808_port_o;
    roundReg_1_3_2[2] <= majority_5809_port_o;
    roundReg_2_3_2[2] <= majority_5810_port_o;
    roundReg_3_3_2[2] <= majority_5811_port_o;
    roundReg_4_3_2[2] <= majority_5812_port_o;
    roundReg_5_3_2[2] <= majority_5813_port_o;
    roundReg_6_3_2[2] <= majority_5814_port_o;
    roundReg_7_3_2[2] <= majority_5815_port_o;
    roundReg_8_3_2[2] <= majority_5816_port_o;
    roundReg_9_3_2[2] <= majority_5817_port_o;
    roundReg_10_3_2[2] <= majority_5818_port_o;
    roundReg_11_3_2[2] <= majority_5819_port_o;
    roundReg_12_3_2[2] <= majority_5820_port_o;
    roundReg_13_3_2[2] <= majority_5821_port_o;
    roundReg_14_3_2[2] <= majority_5822_port_o;
    roundReg_15_3_2[2] <= majority_5823_port_o;
    roundReg_0_0_3[2] <= majority_5824_port_o;
    roundReg_1_0_3[2] <= majority_5825_port_o;
    roundReg_2_0_3[2] <= majority_5826_port_o;
    roundReg_3_0_3[2] <= majority_5827_port_o;
    roundReg_4_0_3[2] <= majority_5828_port_o;
    roundReg_5_0_3[2] <= majority_5829_port_o;
    roundReg_6_0_3[2] <= majority_5830_port_o;
    roundReg_7_0_3[2] <= majority_5831_port_o;
    roundReg_8_0_3[2] <= majority_5832_port_o;
    roundReg_9_0_3[2] <= majority_5833_port_o;
    roundReg_10_0_3[2] <= majority_5834_port_o;
    roundReg_11_0_3[2] <= majority_5835_port_o;
    roundReg_12_0_3[2] <= majority_5836_port_o;
    roundReg_13_0_3[2] <= majority_5837_port_o;
    roundReg_14_0_3[2] <= majority_5838_port_o;
    roundReg_15_0_3[2] <= majority_5839_port_o;
    roundReg_0_1_3[2] <= majority_5840_port_o;
    roundReg_1_1_3[2] <= majority_5841_port_o;
    roundReg_2_1_3[2] <= majority_5842_port_o;
    roundReg_3_1_3[2] <= majority_5843_port_o;
    roundReg_4_1_3[2] <= majority_5844_port_o;
    roundReg_5_1_3[2] <= majority_5845_port_o;
    roundReg_6_1_3[2] <= majority_5846_port_o;
    roundReg_7_1_3[2] <= majority_5847_port_o;
    roundReg_8_1_3[2] <= majority_5848_port_o;
    roundReg_9_1_3[2] <= majority_5849_port_o;
    roundReg_10_1_3[2] <= majority_5850_port_o;
    roundReg_11_1_3[2] <= majority_5851_port_o;
    roundReg_12_1_3[2] <= majority_5852_port_o;
    roundReg_13_1_3[2] <= majority_5853_port_o;
    roundReg_14_1_3[2] <= majority_5854_port_o;
    roundReg_15_1_3[2] <= majority_5855_port_o;
    roundReg_0_2_3[2] <= majority_5856_port_o;
    roundReg_1_2_3[2] <= majority_5857_port_o;
    roundReg_2_2_3[2] <= majority_5858_port_o;
    roundReg_3_2_3[2] <= majority_5859_port_o;
    roundReg_4_2_3[2] <= majority_5860_port_o;
    roundReg_5_2_3[2] <= majority_5861_port_o;
    roundReg_6_2_3[2] <= majority_5862_port_o;
    roundReg_7_2_3[2] <= majority_5863_port_o;
    roundReg_8_2_3[2] <= majority_5864_port_o;
    roundReg_9_2_3[2] <= majority_5865_port_o;
    roundReg_10_2_3[2] <= majority_5866_port_o;
    roundReg_11_2_3[2] <= majority_5867_port_o;
    roundReg_12_2_3[2] <= majority_5868_port_o;
    roundReg_13_2_3[2] <= majority_5869_port_o;
    roundReg_14_2_3[2] <= majority_5870_port_o;
    roundReg_15_2_3[2] <= majority_5871_port_o;
    roundReg_0_3_3[2] <= majority_5872_port_o;
    roundReg_1_3_3[2] <= majority_5873_port_o;
    roundReg_2_3_3[2] <= majority_5874_port_o;
    roundReg_3_3_3[2] <= majority_5875_port_o;
    roundReg_4_3_3[2] <= majority_5876_port_o;
    roundReg_5_3_3[2] <= majority_5877_port_o;
    roundReg_6_3_3[2] <= majority_5878_port_o;
    roundReg_7_3_3[2] <= majority_5879_port_o;
    roundReg_8_3_3[2] <= majority_5880_port_o;
    roundReg_9_3_3[2] <= majority_5881_port_o;
    roundReg_10_3_3[2] <= majority_5882_port_o;
    roundReg_11_3_3[2] <= majority_5883_port_o;
    roundReg_12_3_3[2] <= majority_5884_port_o;
    roundReg_13_3_3[2] <= majority_5885_port_o;
    roundReg_14_3_3[2] <= majority_5886_port_o;
    roundReg_15_3_3[2] <= majority_5887_port_o;
    roundReg_0_0_4[2] <= majority_5888_port_o;
    roundReg_1_0_4[2] <= majority_5889_port_o;
    roundReg_2_0_4[2] <= majority_5890_port_o;
    roundReg_3_0_4[2] <= majority_5891_port_o;
    roundReg_4_0_4[2] <= majority_5892_port_o;
    roundReg_5_0_4[2] <= majority_5893_port_o;
    roundReg_6_0_4[2] <= majority_5894_port_o;
    roundReg_7_0_4[2] <= majority_5895_port_o;
    roundReg_8_0_4[2] <= majority_5896_port_o;
    roundReg_9_0_4[2] <= majority_5897_port_o;
    roundReg_10_0_4[2] <= majority_5898_port_o;
    roundReg_11_0_4[2] <= majority_5899_port_o;
    roundReg_12_0_4[2] <= majority_5900_port_o;
    roundReg_13_0_4[2] <= majority_5901_port_o;
    roundReg_14_0_4[2] <= majority_5902_port_o;
    roundReg_15_0_4[2] <= majority_5903_port_o;
    roundReg_0_1_4[2] <= majority_5904_port_o;
    roundReg_1_1_4[2] <= majority_5905_port_o;
    roundReg_2_1_4[2] <= majority_5906_port_o;
    roundReg_3_1_4[2] <= majority_5907_port_o;
    roundReg_4_1_4[2] <= majority_5908_port_o;
    roundReg_5_1_4[2] <= majority_5909_port_o;
    roundReg_6_1_4[2] <= majority_5910_port_o;
    roundReg_7_1_4[2] <= majority_5911_port_o;
    roundReg_8_1_4[2] <= majority_5912_port_o;
    roundReg_9_1_4[2] <= majority_5913_port_o;
    roundReg_10_1_4[2] <= majority_5914_port_o;
    roundReg_11_1_4[2] <= majority_5915_port_o;
    roundReg_12_1_4[2] <= majority_5916_port_o;
    roundReg_13_1_4[2] <= majority_5917_port_o;
    roundReg_14_1_4[2] <= majority_5918_port_o;
    roundReg_15_1_4[2] <= majority_5919_port_o;
    roundReg_0_2_4[2] <= majority_5920_port_o;
    roundReg_1_2_4[2] <= majority_5921_port_o;
    roundReg_2_2_4[2] <= majority_5922_port_o;
    roundReg_3_2_4[2] <= majority_5923_port_o;
    roundReg_4_2_4[2] <= majority_5924_port_o;
    roundReg_5_2_4[2] <= majority_5925_port_o;
    roundReg_6_2_4[2] <= majority_5926_port_o;
    roundReg_7_2_4[2] <= majority_5927_port_o;
    roundReg_8_2_4[2] <= majority_5928_port_o;
    roundReg_9_2_4[2] <= majority_5929_port_o;
    roundReg_10_2_4[2] <= majority_5930_port_o;
    roundReg_11_2_4[2] <= majority_5931_port_o;
    roundReg_12_2_4[2] <= majority_5932_port_o;
    roundReg_13_2_4[2] <= majority_5933_port_o;
    roundReg_14_2_4[2] <= majority_5934_port_o;
    roundReg_15_2_4[2] <= majority_5935_port_o;
    roundReg_0_3_4[2] <= majority_5936_port_o;
    roundReg_1_3_4[2] <= majority_5937_port_o;
    roundReg_2_3_4[2] <= majority_5938_port_o;
    roundReg_3_3_4[2] <= majority_5939_port_o;
    roundReg_4_3_4[2] <= majority_5940_port_o;
    roundReg_5_3_4[2] <= majority_5941_port_o;
    roundReg_6_3_4[2] <= majority_5942_port_o;
    roundReg_7_3_4[2] <= majority_5943_port_o;
    roundReg_8_3_4[2] <= majority_5944_port_o;
    roundReg_9_3_4[2] <= majority_5945_port_o;
    roundReg_10_3_4[2] <= majority_5946_port_o;
    roundReg_11_3_4[2] <= majority_5947_port_o;
    roundReg_12_3_4[2] <= majority_5948_port_o;
    roundReg_13_3_4[2] <= majority_5949_port_o;
    roundReg_14_3_4[2] <= majority_5950_port_o;
    roundReg_15_3_4[2] <= majority_5951_port_o;
    roundReg_0_0_5[2] <= majority_5952_port_o;
    roundReg_1_0_5[2] <= majority_5953_port_o;
    roundReg_2_0_5[2] <= majority_5954_port_o;
    roundReg_3_0_5[2] <= majority_5955_port_o;
    roundReg_4_0_5[2] <= majority_5956_port_o;
    roundReg_5_0_5[2] <= majority_5957_port_o;
    roundReg_6_0_5[2] <= majority_5958_port_o;
    roundReg_7_0_5[2] <= majority_5959_port_o;
    roundReg_8_0_5[2] <= majority_5960_port_o;
    roundReg_9_0_5[2] <= majority_5961_port_o;
    roundReg_10_0_5[2] <= majority_5962_port_o;
    roundReg_11_0_5[2] <= majority_5963_port_o;
    roundReg_12_0_5[2] <= majority_5964_port_o;
    roundReg_13_0_5[2] <= majority_5965_port_o;
    roundReg_14_0_5[2] <= majority_5966_port_o;
    roundReg_15_0_5[2] <= majority_5967_port_o;
    roundReg_0_1_5[2] <= majority_5968_port_o;
    roundReg_1_1_5[2] <= majority_5969_port_o;
    roundReg_2_1_5[2] <= majority_5970_port_o;
    roundReg_3_1_5[2] <= majority_5971_port_o;
    roundReg_4_1_5[2] <= majority_5972_port_o;
    roundReg_5_1_5[2] <= majority_5973_port_o;
    roundReg_6_1_5[2] <= majority_5974_port_o;
    roundReg_7_1_5[2] <= majority_5975_port_o;
    roundReg_8_1_5[2] <= majority_5976_port_o;
    roundReg_9_1_5[2] <= majority_5977_port_o;
    roundReg_10_1_5[2] <= majority_5978_port_o;
    roundReg_11_1_5[2] <= majority_5979_port_o;
    roundReg_12_1_5[2] <= majority_5980_port_o;
    roundReg_13_1_5[2] <= majority_5981_port_o;
    roundReg_14_1_5[2] <= majority_5982_port_o;
    roundReg_15_1_5[2] <= majority_5983_port_o;
    roundReg_0_2_5[2] <= majority_5984_port_o;
    roundReg_1_2_5[2] <= majority_5985_port_o;
    roundReg_2_2_5[2] <= majority_5986_port_o;
    roundReg_3_2_5[2] <= majority_5987_port_o;
    roundReg_4_2_5[2] <= majority_5988_port_o;
    roundReg_5_2_5[2] <= majority_5989_port_o;
    roundReg_6_2_5[2] <= majority_5990_port_o;
    roundReg_7_2_5[2] <= majority_5991_port_o;
    roundReg_8_2_5[2] <= majority_5992_port_o;
    roundReg_9_2_5[2] <= majority_5993_port_o;
    roundReg_10_2_5[2] <= majority_5994_port_o;
    roundReg_11_2_5[2] <= majority_5995_port_o;
    roundReg_12_2_5[2] <= majority_5996_port_o;
    roundReg_13_2_5[2] <= majority_5997_port_o;
    roundReg_14_2_5[2] <= majority_5998_port_o;
    roundReg_15_2_5[2] <= majority_5999_port_o;
    roundReg_0_3_5[2] <= majority_6000_port_o;
    roundReg_1_3_5[2] <= majority_6001_port_o;
    roundReg_2_3_5[2] <= majority_6002_port_o;
    roundReg_3_3_5[2] <= majority_6003_port_o;
    roundReg_4_3_5[2] <= majority_6004_port_o;
    roundReg_5_3_5[2] <= majority_6005_port_o;
    roundReg_6_3_5[2] <= majority_6006_port_o;
    roundReg_7_3_5[2] <= majority_6007_port_o;
    roundReg_8_3_5[2] <= majority_6008_port_o;
    roundReg_9_3_5[2] <= majority_6009_port_o;
    roundReg_10_3_5[2] <= majority_6010_port_o;
    roundReg_11_3_5[2] <= majority_6011_port_o;
    roundReg_12_3_5[2] <= majority_6012_port_o;
    roundReg_13_3_5[2] <= majority_6013_port_o;
    roundReg_14_3_5[2] <= majority_6014_port_o;
    roundReg_15_3_5[2] <= majority_6015_port_o;
    roundReg_0_0_6[2] <= majority_6016_port_o;
    roundReg_1_0_6[2] <= majority_6017_port_o;
    roundReg_2_0_6[2] <= majority_6018_port_o;
    roundReg_3_0_6[2] <= majority_6019_port_o;
    roundReg_4_0_6[2] <= majority_6020_port_o;
    roundReg_5_0_6[2] <= majority_6021_port_o;
    roundReg_6_0_6[2] <= majority_6022_port_o;
    roundReg_7_0_6[2] <= majority_6023_port_o;
    roundReg_8_0_6[2] <= majority_6024_port_o;
    roundReg_9_0_6[2] <= majority_6025_port_o;
    roundReg_10_0_6[2] <= majority_6026_port_o;
    roundReg_11_0_6[2] <= majority_6027_port_o;
    roundReg_12_0_6[2] <= majority_6028_port_o;
    roundReg_13_0_6[2] <= majority_6029_port_o;
    roundReg_14_0_6[2] <= majority_6030_port_o;
    roundReg_15_0_6[2] <= majority_6031_port_o;
    roundReg_0_1_6[2] <= majority_6032_port_o;
    roundReg_1_1_6[2] <= majority_6033_port_o;
    roundReg_2_1_6[2] <= majority_6034_port_o;
    roundReg_3_1_6[2] <= majority_6035_port_o;
    roundReg_4_1_6[2] <= majority_6036_port_o;
    roundReg_5_1_6[2] <= majority_6037_port_o;
    roundReg_6_1_6[2] <= majority_6038_port_o;
    roundReg_7_1_6[2] <= majority_6039_port_o;
    roundReg_8_1_6[2] <= majority_6040_port_o;
    roundReg_9_1_6[2] <= majority_6041_port_o;
    roundReg_10_1_6[2] <= majority_6042_port_o;
    roundReg_11_1_6[2] <= majority_6043_port_o;
    roundReg_12_1_6[2] <= majority_6044_port_o;
    roundReg_13_1_6[2] <= majority_6045_port_o;
    roundReg_14_1_6[2] <= majority_6046_port_o;
    roundReg_15_1_6[2] <= majority_6047_port_o;
    roundReg_0_2_6[2] <= majority_6048_port_o;
    roundReg_1_2_6[2] <= majority_6049_port_o;
    roundReg_2_2_6[2] <= majority_6050_port_o;
    roundReg_3_2_6[2] <= majority_6051_port_o;
    roundReg_4_2_6[2] <= majority_6052_port_o;
    roundReg_5_2_6[2] <= majority_6053_port_o;
    roundReg_6_2_6[2] <= majority_6054_port_o;
    roundReg_7_2_6[2] <= majority_6055_port_o;
    roundReg_8_2_6[2] <= majority_6056_port_o;
    roundReg_9_2_6[2] <= majority_6057_port_o;
    roundReg_10_2_6[2] <= majority_6058_port_o;
    roundReg_11_2_6[2] <= majority_6059_port_o;
    roundReg_12_2_6[2] <= majority_6060_port_o;
    roundReg_13_2_6[2] <= majority_6061_port_o;
    roundReg_14_2_6[2] <= majority_6062_port_o;
    roundReg_15_2_6[2] <= majority_6063_port_o;
    roundReg_0_3_6[2] <= majority_6064_port_o;
    roundReg_1_3_6[2] <= majority_6065_port_o;
    roundReg_2_3_6[2] <= majority_6066_port_o;
    roundReg_3_3_6[2] <= majority_6067_port_o;
    roundReg_4_3_6[2] <= majority_6068_port_o;
    roundReg_5_3_6[2] <= majority_6069_port_o;
    roundReg_6_3_6[2] <= majority_6070_port_o;
    roundReg_7_3_6[2] <= majority_6071_port_o;
    roundReg_8_3_6[2] <= majority_6072_port_o;
    roundReg_9_3_6[2] <= majority_6073_port_o;
    roundReg_10_3_6[2] <= majority_6074_port_o;
    roundReg_11_3_6[2] <= majority_6075_port_o;
    roundReg_12_3_6[2] <= majority_6076_port_o;
    roundReg_13_3_6[2] <= majority_6077_port_o;
    roundReg_14_3_6[2] <= majority_6078_port_o;
    roundReg_15_3_6[2] <= majority_6079_port_o;
    roundReg_0_0_7[2] <= majority_6080_port_o;
    roundReg_1_0_7[2] <= majority_6081_port_o;
    roundReg_2_0_7[2] <= majority_6082_port_o;
    roundReg_3_0_7[2] <= majority_6083_port_o;
    roundReg_4_0_7[2] <= majority_6084_port_o;
    roundReg_5_0_7[2] <= majority_6085_port_o;
    roundReg_6_0_7[2] <= majority_6086_port_o;
    roundReg_7_0_7[2] <= majority_6087_port_o;
    roundReg_8_0_7[2] <= majority_6088_port_o;
    roundReg_9_0_7[2] <= majority_6089_port_o;
    roundReg_10_0_7[2] <= majority_6090_port_o;
    roundReg_11_0_7[2] <= majority_6091_port_o;
    roundReg_12_0_7[2] <= majority_6092_port_o;
    roundReg_13_0_7[2] <= majority_6093_port_o;
    roundReg_14_0_7[2] <= majority_6094_port_o;
    roundReg_15_0_7[2] <= majority_6095_port_o;
    roundReg_0_1_7[2] <= majority_6096_port_o;
    roundReg_1_1_7[2] <= majority_6097_port_o;
    roundReg_2_1_7[2] <= majority_6098_port_o;
    roundReg_3_1_7[2] <= majority_6099_port_o;
    roundReg_4_1_7[2] <= majority_6100_port_o;
    roundReg_5_1_7[2] <= majority_6101_port_o;
    roundReg_6_1_7[2] <= majority_6102_port_o;
    roundReg_7_1_7[2] <= majority_6103_port_o;
    roundReg_8_1_7[2] <= majority_6104_port_o;
    roundReg_9_1_7[2] <= majority_6105_port_o;
    roundReg_10_1_7[2] <= majority_6106_port_o;
    roundReg_11_1_7[2] <= majority_6107_port_o;
    roundReg_12_1_7[2] <= majority_6108_port_o;
    roundReg_13_1_7[2] <= majority_6109_port_o;
    roundReg_14_1_7[2] <= majority_6110_port_o;
    roundReg_15_1_7[2] <= majority_6111_port_o;
    roundReg_0_2_7[2] <= majority_6112_port_o;
    roundReg_1_2_7[2] <= majority_6113_port_o;
    roundReg_2_2_7[2] <= majority_6114_port_o;
    roundReg_3_2_7[2] <= majority_6115_port_o;
    roundReg_4_2_7[2] <= majority_6116_port_o;
    roundReg_5_2_7[2] <= majority_6117_port_o;
    roundReg_6_2_7[2] <= majority_6118_port_o;
    roundReg_7_2_7[2] <= majority_6119_port_o;
    roundReg_8_2_7[2] <= majority_6120_port_o;
    roundReg_9_2_7[2] <= majority_6121_port_o;
    roundReg_10_2_7[2] <= majority_6122_port_o;
    roundReg_11_2_7[2] <= majority_6123_port_o;
    roundReg_12_2_7[2] <= majority_6124_port_o;
    roundReg_13_2_7[2] <= majority_6125_port_o;
    roundReg_14_2_7[2] <= majority_6126_port_o;
    roundReg_15_2_7[2] <= majority_6127_port_o;
    roundReg_0_3_7[2] <= majority_6128_port_o;
    roundReg_1_3_7[2] <= majority_6129_port_o;
    roundReg_2_3_7[2] <= majority_6130_port_o;
    roundReg_3_3_7[2] <= majority_6131_port_o;
    roundReg_4_3_7[2] <= majority_6132_port_o;
    roundReg_5_3_7[2] <= majority_6133_port_o;
    roundReg_6_3_7[2] <= majority_6134_port_o;
    roundReg_7_3_7[2] <= majority_6135_port_o;
    roundReg_8_3_7[2] <= majority_6136_port_o;
    roundReg_9_3_7[2] <= majority_6137_port_o;
    roundReg_10_3_7[2] <= majority_6138_port_o;
    roundReg_11_3_7[2] <= majority_6139_port_o;
    roundReg_12_3_7[2] <= majority_6140_port_o;
    roundReg_13_3_7[2] <= majority_6141_port_o;
    roundReg_14_3_7[2] <= majority_6142_port_o;
    roundReg_15_3_7[2] <= majority_6143_port_o;
  end


endmodule

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

module Aes_MixColumn (
  input      [2:0]    port_state_in_0_0_0,
  input      [2:0]    port_state_in_0_0_1,
  input      [2:0]    port_state_in_0_0_2,
  input      [2:0]    port_state_in_0_0_3,
  input      [2:0]    port_state_in_0_0_4,
  input      [2:0]    port_state_in_0_0_5,
  input      [2:0]    port_state_in_0_0_6,
  input      [2:0]    port_state_in_0_0_7,
  input      [2:0]    port_state_in_0_1_0,
  input      [2:0]    port_state_in_0_1_1,
  input      [2:0]    port_state_in_0_1_2,
  input      [2:0]    port_state_in_0_1_3,
  input      [2:0]    port_state_in_0_1_4,
  input      [2:0]    port_state_in_0_1_5,
  input      [2:0]    port_state_in_0_1_6,
  input      [2:0]    port_state_in_0_1_7,
  input      [2:0]    port_state_in_0_2_0,
  input      [2:0]    port_state_in_0_2_1,
  input      [2:0]    port_state_in_0_2_2,
  input      [2:0]    port_state_in_0_2_3,
  input      [2:0]    port_state_in_0_2_4,
  input      [2:0]    port_state_in_0_2_5,
  input      [2:0]    port_state_in_0_2_6,
  input      [2:0]    port_state_in_0_2_7,
  input      [2:0]    port_state_in_0_3_0,
  input      [2:0]    port_state_in_0_3_1,
  input      [2:0]    port_state_in_0_3_2,
  input      [2:0]    port_state_in_0_3_3,
  input      [2:0]    port_state_in_0_3_4,
  input      [2:0]    port_state_in_0_3_5,
  input      [2:0]    port_state_in_0_3_6,
  input      [2:0]    port_state_in_0_3_7,
  input      [2:0]    port_state_in_1_0_0,
  input      [2:0]    port_state_in_1_0_1,
  input      [2:0]    port_state_in_1_0_2,
  input      [2:0]    port_state_in_1_0_3,
  input      [2:0]    port_state_in_1_0_4,
  input      [2:0]    port_state_in_1_0_5,
  input      [2:0]    port_state_in_1_0_6,
  input      [2:0]    port_state_in_1_0_7,
  input      [2:0]    port_state_in_1_1_0,
  input      [2:0]    port_state_in_1_1_1,
  input      [2:0]    port_state_in_1_1_2,
  input      [2:0]    port_state_in_1_1_3,
  input      [2:0]    port_state_in_1_1_4,
  input      [2:0]    port_state_in_1_1_5,
  input      [2:0]    port_state_in_1_1_6,
  input      [2:0]    port_state_in_1_1_7,
  input      [2:0]    port_state_in_1_2_0,
  input      [2:0]    port_state_in_1_2_1,
  input      [2:0]    port_state_in_1_2_2,
  input      [2:0]    port_state_in_1_2_3,
  input      [2:0]    port_state_in_1_2_4,
  input      [2:0]    port_state_in_1_2_5,
  input      [2:0]    port_state_in_1_2_6,
  input      [2:0]    port_state_in_1_2_7,
  input      [2:0]    port_state_in_1_3_0,
  input      [2:0]    port_state_in_1_3_1,
  input      [2:0]    port_state_in_1_3_2,
  input      [2:0]    port_state_in_1_3_3,
  input      [2:0]    port_state_in_1_3_4,
  input      [2:0]    port_state_in_1_3_5,
  input      [2:0]    port_state_in_1_3_6,
  input      [2:0]    port_state_in_1_3_7,
  input      [2:0]    port_state_in_2_0_0,
  input      [2:0]    port_state_in_2_0_1,
  input      [2:0]    port_state_in_2_0_2,
  input      [2:0]    port_state_in_2_0_3,
  input      [2:0]    port_state_in_2_0_4,
  input      [2:0]    port_state_in_2_0_5,
  input      [2:0]    port_state_in_2_0_6,
  input      [2:0]    port_state_in_2_0_7,
  input      [2:0]    port_state_in_2_1_0,
  input      [2:0]    port_state_in_2_1_1,
  input      [2:0]    port_state_in_2_1_2,
  input      [2:0]    port_state_in_2_1_3,
  input      [2:0]    port_state_in_2_1_4,
  input      [2:0]    port_state_in_2_1_5,
  input      [2:0]    port_state_in_2_1_6,
  input      [2:0]    port_state_in_2_1_7,
  input      [2:0]    port_state_in_2_2_0,
  input      [2:0]    port_state_in_2_2_1,
  input      [2:0]    port_state_in_2_2_2,
  input      [2:0]    port_state_in_2_2_3,
  input      [2:0]    port_state_in_2_2_4,
  input      [2:0]    port_state_in_2_2_5,
  input      [2:0]    port_state_in_2_2_6,
  input      [2:0]    port_state_in_2_2_7,
  input      [2:0]    port_state_in_2_3_0,
  input      [2:0]    port_state_in_2_3_1,
  input      [2:0]    port_state_in_2_3_2,
  input      [2:0]    port_state_in_2_3_3,
  input      [2:0]    port_state_in_2_3_4,
  input      [2:0]    port_state_in_2_3_5,
  input      [2:0]    port_state_in_2_3_6,
  input      [2:0]    port_state_in_2_3_7,
  input      [2:0]    port_state_in_3_0_0,
  input      [2:0]    port_state_in_3_0_1,
  input      [2:0]    port_state_in_3_0_2,
  input      [2:0]    port_state_in_3_0_3,
  input      [2:0]    port_state_in_3_0_4,
  input      [2:0]    port_state_in_3_0_5,
  input      [2:0]    port_state_in_3_0_6,
  input      [2:0]    port_state_in_3_0_7,
  input      [2:0]    port_state_in_3_1_0,
  input      [2:0]    port_state_in_3_1_1,
  input      [2:0]    port_state_in_3_1_2,
  input      [2:0]    port_state_in_3_1_3,
  input      [2:0]    port_state_in_3_1_4,
  input      [2:0]    port_state_in_3_1_5,
  input      [2:0]    port_state_in_3_1_6,
  input      [2:0]    port_state_in_3_1_7,
  input      [2:0]    port_state_in_3_2_0,
  input      [2:0]    port_state_in_3_2_1,
  input      [2:0]    port_state_in_3_2_2,
  input      [2:0]    port_state_in_3_2_3,
  input      [2:0]    port_state_in_3_2_4,
  input      [2:0]    port_state_in_3_2_5,
  input      [2:0]    port_state_in_3_2_6,
  input      [2:0]    port_state_in_3_2_7,
  input      [2:0]    port_state_in_3_3_0,
  input      [2:0]    port_state_in_3_3_1,
  input      [2:0]    port_state_in_3_3_2,
  input      [2:0]    port_state_in_3_3_3,
  input      [2:0]    port_state_in_3_3_4,
  input      [2:0]    port_state_in_3_3_5,
  input      [2:0]    port_state_in_3_3_6,
  input      [2:0]    port_state_in_3_3_7,
  input      [2:0]    port_state_in_4_0_0,
  input      [2:0]    port_state_in_4_0_1,
  input      [2:0]    port_state_in_4_0_2,
  input      [2:0]    port_state_in_4_0_3,
  input      [2:0]    port_state_in_4_0_4,
  input      [2:0]    port_state_in_4_0_5,
  input      [2:0]    port_state_in_4_0_6,
  input      [2:0]    port_state_in_4_0_7,
  input      [2:0]    port_state_in_4_1_0,
  input      [2:0]    port_state_in_4_1_1,
  input      [2:0]    port_state_in_4_1_2,
  input      [2:0]    port_state_in_4_1_3,
  input      [2:0]    port_state_in_4_1_4,
  input      [2:0]    port_state_in_4_1_5,
  input      [2:0]    port_state_in_4_1_6,
  input      [2:0]    port_state_in_4_1_7,
  input      [2:0]    port_state_in_4_2_0,
  input      [2:0]    port_state_in_4_2_1,
  input      [2:0]    port_state_in_4_2_2,
  input      [2:0]    port_state_in_4_2_3,
  input      [2:0]    port_state_in_4_2_4,
  input      [2:0]    port_state_in_4_2_5,
  input      [2:0]    port_state_in_4_2_6,
  input      [2:0]    port_state_in_4_2_7,
  input      [2:0]    port_state_in_4_3_0,
  input      [2:0]    port_state_in_4_3_1,
  input      [2:0]    port_state_in_4_3_2,
  input      [2:0]    port_state_in_4_3_3,
  input      [2:0]    port_state_in_4_3_4,
  input      [2:0]    port_state_in_4_3_5,
  input      [2:0]    port_state_in_4_3_6,
  input      [2:0]    port_state_in_4_3_7,
  input      [2:0]    port_state_in_5_0_0,
  input      [2:0]    port_state_in_5_0_1,
  input      [2:0]    port_state_in_5_0_2,
  input      [2:0]    port_state_in_5_0_3,
  input      [2:0]    port_state_in_5_0_4,
  input      [2:0]    port_state_in_5_0_5,
  input      [2:0]    port_state_in_5_0_6,
  input      [2:0]    port_state_in_5_0_7,
  input      [2:0]    port_state_in_5_1_0,
  input      [2:0]    port_state_in_5_1_1,
  input      [2:0]    port_state_in_5_1_2,
  input      [2:0]    port_state_in_5_1_3,
  input      [2:0]    port_state_in_5_1_4,
  input      [2:0]    port_state_in_5_1_5,
  input      [2:0]    port_state_in_5_1_6,
  input      [2:0]    port_state_in_5_1_7,
  input      [2:0]    port_state_in_5_2_0,
  input      [2:0]    port_state_in_5_2_1,
  input      [2:0]    port_state_in_5_2_2,
  input      [2:0]    port_state_in_5_2_3,
  input      [2:0]    port_state_in_5_2_4,
  input      [2:0]    port_state_in_5_2_5,
  input      [2:0]    port_state_in_5_2_6,
  input      [2:0]    port_state_in_5_2_7,
  input      [2:0]    port_state_in_5_3_0,
  input      [2:0]    port_state_in_5_3_1,
  input      [2:0]    port_state_in_5_3_2,
  input      [2:0]    port_state_in_5_3_3,
  input      [2:0]    port_state_in_5_3_4,
  input      [2:0]    port_state_in_5_3_5,
  input      [2:0]    port_state_in_5_3_6,
  input      [2:0]    port_state_in_5_3_7,
  input      [2:0]    port_state_in_6_0_0,
  input      [2:0]    port_state_in_6_0_1,
  input      [2:0]    port_state_in_6_0_2,
  input      [2:0]    port_state_in_6_0_3,
  input      [2:0]    port_state_in_6_0_4,
  input      [2:0]    port_state_in_6_0_5,
  input      [2:0]    port_state_in_6_0_6,
  input      [2:0]    port_state_in_6_0_7,
  input      [2:0]    port_state_in_6_1_0,
  input      [2:0]    port_state_in_6_1_1,
  input      [2:0]    port_state_in_6_1_2,
  input      [2:0]    port_state_in_6_1_3,
  input      [2:0]    port_state_in_6_1_4,
  input      [2:0]    port_state_in_6_1_5,
  input      [2:0]    port_state_in_6_1_6,
  input      [2:0]    port_state_in_6_1_7,
  input      [2:0]    port_state_in_6_2_0,
  input      [2:0]    port_state_in_6_2_1,
  input      [2:0]    port_state_in_6_2_2,
  input      [2:0]    port_state_in_6_2_3,
  input      [2:0]    port_state_in_6_2_4,
  input      [2:0]    port_state_in_6_2_5,
  input      [2:0]    port_state_in_6_2_6,
  input      [2:0]    port_state_in_6_2_7,
  input      [2:0]    port_state_in_6_3_0,
  input      [2:0]    port_state_in_6_3_1,
  input      [2:0]    port_state_in_6_3_2,
  input      [2:0]    port_state_in_6_3_3,
  input      [2:0]    port_state_in_6_3_4,
  input      [2:0]    port_state_in_6_3_5,
  input      [2:0]    port_state_in_6_3_6,
  input      [2:0]    port_state_in_6_3_7,
  input      [2:0]    port_state_in_7_0_0,
  input      [2:0]    port_state_in_7_0_1,
  input      [2:0]    port_state_in_7_0_2,
  input      [2:0]    port_state_in_7_0_3,
  input      [2:0]    port_state_in_7_0_4,
  input      [2:0]    port_state_in_7_0_5,
  input      [2:0]    port_state_in_7_0_6,
  input      [2:0]    port_state_in_7_0_7,
  input      [2:0]    port_state_in_7_1_0,
  input      [2:0]    port_state_in_7_1_1,
  input      [2:0]    port_state_in_7_1_2,
  input      [2:0]    port_state_in_7_1_3,
  input      [2:0]    port_state_in_7_1_4,
  input      [2:0]    port_state_in_7_1_5,
  input      [2:0]    port_state_in_7_1_6,
  input      [2:0]    port_state_in_7_1_7,
  input      [2:0]    port_state_in_7_2_0,
  input      [2:0]    port_state_in_7_2_1,
  input      [2:0]    port_state_in_7_2_2,
  input      [2:0]    port_state_in_7_2_3,
  input      [2:0]    port_state_in_7_2_4,
  input      [2:0]    port_state_in_7_2_5,
  input      [2:0]    port_state_in_7_2_6,
  input      [2:0]    port_state_in_7_2_7,
  input      [2:0]    port_state_in_7_3_0,
  input      [2:0]    port_state_in_7_3_1,
  input      [2:0]    port_state_in_7_3_2,
  input      [2:0]    port_state_in_7_3_3,
  input      [2:0]    port_state_in_7_3_4,
  input      [2:0]    port_state_in_7_3_5,
  input      [2:0]    port_state_in_7_3_6,
  input      [2:0]    port_state_in_7_3_7,
  input      [2:0]    port_state_in_8_0_0,
  input      [2:0]    port_state_in_8_0_1,
  input      [2:0]    port_state_in_8_0_2,
  input      [2:0]    port_state_in_8_0_3,
  input      [2:0]    port_state_in_8_0_4,
  input      [2:0]    port_state_in_8_0_5,
  input      [2:0]    port_state_in_8_0_6,
  input      [2:0]    port_state_in_8_0_7,
  input      [2:0]    port_state_in_8_1_0,
  input      [2:0]    port_state_in_8_1_1,
  input      [2:0]    port_state_in_8_1_2,
  input      [2:0]    port_state_in_8_1_3,
  input      [2:0]    port_state_in_8_1_4,
  input      [2:0]    port_state_in_8_1_5,
  input      [2:0]    port_state_in_8_1_6,
  input      [2:0]    port_state_in_8_1_7,
  input      [2:0]    port_state_in_8_2_0,
  input      [2:0]    port_state_in_8_2_1,
  input      [2:0]    port_state_in_8_2_2,
  input      [2:0]    port_state_in_8_2_3,
  input      [2:0]    port_state_in_8_2_4,
  input      [2:0]    port_state_in_8_2_5,
  input      [2:0]    port_state_in_8_2_6,
  input      [2:0]    port_state_in_8_2_7,
  input      [2:0]    port_state_in_8_3_0,
  input      [2:0]    port_state_in_8_3_1,
  input      [2:0]    port_state_in_8_3_2,
  input      [2:0]    port_state_in_8_3_3,
  input      [2:0]    port_state_in_8_3_4,
  input      [2:0]    port_state_in_8_3_5,
  input      [2:0]    port_state_in_8_3_6,
  input      [2:0]    port_state_in_8_3_7,
  input      [2:0]    port_state_in_9_0_0,
  input      [2:0]    port_state_in_9_0_1,
  input      [2:0]    port_state_in_9_0_2,
  input      [2:0]    port_state_in_9_0_3,
  input      [2:0]    port_state_in_9_0_4,
  input      [2:0]    port_state_in_9_0_5,
  input      [2:0]    port_state_in_9_0_6,
  input      [2:0]    port_state_in_9_0_7,
  input      [2:0]    port_state_in_9_1_0,
  input      [2:0]    port_state_in_9_1_1,
  input      [2:0]    port_state_in_9_1_2,
  input      [2:0]    port_state_in_9_1_3,
  input      [2:0]    port_state_in_9_1_4,
  input      [2:0]    port_state_in_9_1_5,
  input      [2:0]    port_state_in_9_1_6,
  input      [2:0]    port_state_in_9_1_7,
  input      [2:0]    port_state_in_9_2_0,
  input      [2:0]    port_state_in_9_2_1,
  input      [2:0]    port_state_in_9_2_2,
  input      [2:0]    port_state_in_9_2_3,
  input      [2:0]    port_state_in_9_2_4,
  input      [2:0]    port_state_in_9_2_5,
  input      [2:0]    port_state_in_9_2_6,
  input      [2:0]    port_state_in_9_2_7,
  input      [2:0]    port_state_in_9_3_0,
  input      [2:0]    port_state_in_9_3_1,
  input      [2:0]    port_state_in_9_3_2,
  input      [2:0]    port_state_in_9_3_3,
  input      [2:0]    port_state_in_9_3_4,
  input      [2:0]    port_state_in_9_3_5,
  input      [2:0]    port_state_in_9_3_6,
  input      [2:0]    port_state_in_9_3_7,
  input      [2:0]    port_state_in_10_0_0,
  input      [2:0]    port_state_in_10_0_1,
  input      [2:0]    port_state_in_10_0_2,
  input      [2:0]    port_state_in_10_0_3,
  input      [2:0]    port_state_in_10_0_4,
  input      [2:0]    port_state_in_10_0_5,
  input      [2:0]    port_state_in_10_0_6,
  input      [2:0]    port_state_in_10_0_7,
  input      [2:0]    port_state_in_10_1_0,
  input      [2:0]    port_state_in_10_1_1,
  input      [2:0]    port_state_in_10_1_2,
  input      [2:0]    port_state_in_10_1_3,
  input      [2:0]    port_state_in_10_1_4,
  input      [2:0]    port_state_in_10_1_5,
  input      [2:0]    port_state_in_10_1_6,
  input      [2:0]    port_state_in_10_1_7,
  input      [2:0]    port_state_in_10_2_0,
  input      [2:0]    port_state_in_10_2_1,
  input      [2:0]    port_state_in_10_2_2,
  input      [2:0]    port_state_in_10_2_3,
  input      [2:0]    port_state_in_10_2_4,
  input      [2:0]    port_state_in_10_2_5,
  input      [2:0]    port_state_in_10_2_6,
  input      [2:0]    port_state_in_10_2_7,
  input      [2:0]    port_state_in_10_3_0,
  input      [2:0]    port_state_in_10_3_1,
  input      [2:0]    port_state_in_10_3_2,
  input      [2:0]    port_state_in_10_3_3,
  input      [2:0]    port_state_in_10_3_4,
  input      [2:0]    port_state_in_10_3_5,
  input      [2:0]    port_state_in_10_3_6,
  input      [2:0]    port_state_in_10_3_7,
  input      [2:0]    port_state_in_11_0_0,
  input      [2:0]    port_state_in_11_0_1,
  input      [2:0]    port_state_in_11_0_2,
  input      [2:0]    port_state_in_11_0_3,
  input      [2:0]    port_state_in_11_0_4,
  input      [2:0]    port_state_in_11_0_5,
  input      [2:0]    port_state_in_11_0_6,
  input      [2:0]    port_state_in_11_0_7,
  input      [2:0]    port_state_in_11_1_0,
  input      [2:0]    port_state_in_11_1_1,
  input      [2:0]    port_state_in_11_1_2,
  input      [2:0]    port_state_in_11_1_3,
  input      [2:0]    port_state_in_11_1_4,
  input      [2:0]    port_state_in_11_1_5,
  input      [2:0]    port_state_in_11_1_6,
  input      [2:0]    port_state_in_11_1_7,
  input      [2:0]    port_state_in_11_2_0,
  input      [2:0]    port_state_in_11_2_1,
  input      [2:0]    port_state_in_11_2_2,
  input      [2:0]    port_state_in_11_2_3,
  input      [2:0]    port_state_in_11_2_4,
  input      [2:0]    port_state_in_11_2_5,
  input      [2:0]    port_state_in_11_2_6,
  input      [2:0]    port_state_in_11_2_7,
  input      [2:0]    port_state_in_11_3_0,
  input      [2:0]    port_state_in_11_3_1,
  input      [2:0]    port_state_in_11_3_2,
  input      [2:0]    port_state_in_11_3_3,
  input      [2:0]    port_state_in_11_3_4,
  input      [2:0]    port_state_in_11_3_5,
  input      [2:0]    port_state_in_11_3_6,
  input      [2:0]    port_state_in_11_3_7,
  input      [2:0]    port_state_in_12_0_0,
  input      [2:0]    port_state_in_12_0_1,
  input      [2:0]    port_state_in_12_0_2,
  input      [2:0]    port_state_in_12_0_3,
  input      [2:0]    port_state_in_12_0_4,
  input      [2:0]    port_state_in_12_0_5,
  input      [2:0]    port_state_in_12_0_6,
  input      [2:0]    port_state_in_12_0_7,
  input      [2:0]    port_state_in_12_1_0,
  input      [2:0]    port_state_in_12_1_1,
  input      [2:0]    port_state_in_12_1_2,
  input      [2:0]    port_state_in_12_1_3,
  input      [2:0]    port_state_in_12_1_4,
  input      [2:0]    port_state_in_12_1_5,
  input      [2:0]    port_state_in_12_1_6,
  input      [2:0]    port_state_in_12_1_7,
  input      [2:0]    port_state_in_12_2_0,
  input      [2:0]    port_state_in_12_2_1,
  input      [2:0]    port_state_in_12_2_2,
  input      [2:0]    port_state_in_12_2_3,
  input      [2:0]    port_state_in_12_2_4,
  input      [2:0]    port_state_in_12_2_5,
  input      [2:0]    port_state_in_12_2_6,
  input      [2:0]    port_state_in_12_2_7,
  input      [2:0]    port_state_in_12_3_0,
  input      [2:0]    port_state_in_12_3_1,
  input      [2:0]    port_state_in_12_3_2,
  input      [2:0]    port_state_in_12_3_3,
  input      [2:0]    port_state_in_12_3_4,
  input      [2:0]    port_state_in_12_3_5,
  input      [2:0]    port_state_in_12_3_6,
  input      [2:0]    port_state_in_12_3_7,
  input      [2:0]    port_state_in_13_0_0,
  input      [2:0]    port_state_in_13_0_1,
  input      [2:0]    port_state_in_13_0_2,
  input      [2:0]    port_state_in_13_0_3,
  input      [2:0]    port_state_in_13_0_4,
  input      [2:0]    port_state_in_13_0_5,
  input      [2:0]    port_state_in_13_0_6,
  input      [2:0]    port_state_in_13_0_7,
  input      [2:0]    port_state_in_13_1_0,
  input      [2:0]    port_state_in_13_1_1,
  input      [2:0]    port_state_in_13_1_2,
  input      [2:0]    port_state_in_13_1_3,
  input      [2:0]    port_state_in_13_1_4,
  input      [2:0]    port_state_in_13_1_5,
  input      [2:0]    port_state_in_13_1_6,
  input      [2:0]    port_state_in_13_1_7,
  input      [2:0]    port_state_in_13_2_0,
  input      [2:0]    port_state_in_13_2_1,
  input      [2:0]    port_state_in_13_2_2,
  input      [2:0]    port_state_in_13_2_3,
  input      [2:0]    port_state_in_13_2_4,
  input      [2:0]    port_state_in_13_2_5,
  input      [2:0]    port_state_in_13_2_6,
  input      [2:0]    port_state_in_13_2_7,
  input      [2:0]    port_state_in_13_3_0,
  input      [2:0]    port_state_in_13_3_1,
  input      [2:0]    port_state_in_13_3_2,
  input      [2:0]    port_state_in_13_3_3,
  input      [2:0]    port_state_in_13_3_4,
  input      [2:0]    port_state_in_13_3_5,
  input      [2:0]    port_state_in_13_3_6,
  input      [2:0]    port_state_in_13_3_7,
  input      [2:0]    port_state_in_14_0_0,
  input      [2:0]    port_state_in_14_0_1,
  input      [2:0]    port_state_in_14_0_2,
  input      [2:0]    port_state_in_14_0_3,
  input      [2:0]    port_state_in_14_0_4,
  input      [2:0]    port_state_in_14_0_5,
  input      [2:0]    port_state_in_14_0_6,
  input      [2:0]    port_state_in_14_0_7,
  input      [2:0]    port_state_in_14_1_0,
  input      [2:0]    port_state_in_14_1_1,
  input      [2:0]    port_state_in_14_1_2,
  input      [2:0]    port_state_in_14_1_3,
  input      [2:0]    port_state_in_14_1_4,
  input      [2:0]    port_state_in_14_1_5,
  input      [2:0]    port_state_in_14_1_6,
  input      [2:0]    port_state_in_14_1_7,
  input      [2:0]    port_state_in_14_2_0,
  input      [2:0]    port_state_in_14_2_1,
  input      [2:0]    port_state_in_14_2_2,
  input      [2:0]    port_state_in_14_2_3,
  input      [2:0]    port_state_in_14_2_4,
  input      [2:0]    port_state_in_14_2_5,
  input      [2:0]    port_state_in_14_2_6,
  input      [2:0]    port_state_in_14_2_7,
  input      [2:0]    port_state_in_14_3_0,
  input      [2:0]    port_state_in_14_3_1,
  input      [2:0]    port_state_in_14_3_2,
  input      [2:0]    port_state_in_14_3_3,
  input      [2:0]    port_state_in_14_3_4,
  input      [2:0]    port_state_in_14_3_5,
  input      [2:0]    port_state_in_14_3_6,
  input      [2:0]    port_state_in_14_3_7,
  input      [2:0]    port_state_in_15_0_0,
  input      [2:0]    port_state_in_15_0_1,
  input      [2:0]    port_state_in_15_0_2,
  input      [2:0]    port_state_in_15_0_3,
  input      [2:0]    port_state_in_15_0_4,
  input      [2:0]    port_state_in_15_0_5,
  input      [2:0]    port_state_in_15_0_6,
  input      [2:0]    port_state_in_15_0_7,
  input      [2:0]    port_state_in_15_1_0,
  input      [2:0]    port_state_in_15_1_1,
  input      [2:0]    port_state_in_15_1_2,
  input      [2:0]    port_state_in_15_1_3,
  input      [2:0]    port_state_in_15_1_4,
  input      [2:0]    port_state_in_15_1_5,
  input      [2:0]    port_state_in_15_1_6,
  input      [2:0]    port_state_in_15_1_7,
  input      [2:0]    port_state_in_15_2_0,
  input      [2:0]    port_state_in_15_2_1,
  input      [2:0]    port_state_in_15_2_2,
  input      [2:0]    port_state_in_15_2_3,
  input      [2:0]    port_state_in_15_2_4,
  input      [2:0]    port_state_in_15_2_5,
  input      [2:0]    port_state_in_15_2_6,
  input      [2:0]    port_state_in_15_2_7,
  input      [2:0]    port_state_in_15_3_0,
  input      [2:0]    port_state_in_15_3_1,
  input      [2:0]    port_state_in_15_3_2,
  input      [2:0]    port_state_in_15_3_3,
  input      [2:0]    port_state_in_15_3_4,
  input      [2:0]    port_state_in_15_3_5,
  input      [2:0]    port_state_in_15_3_6,
  input      [2:0]    port_state_in_15_3_7,
  output     [2:0]    port_state_out_0_0_0,
  output     [2:0]    port_state_out_0_0_1,
  output     [2:0]    port_state_out_0_0_2,
  output     [2:0]    port_state_out_0_0_3,
  output     [2:0]    port_state_out_0_0_4,
  output     [2:0]    port_state_out_0_0_5,
  output     [2:0]    port_state_out_0_0_6,
  output     [2:0]    port_state_out_0_0_7,
  output     [2:0]    port_state_out_0_1_0,
  output     [2:0]    port_state_out_0_1_1,
  output     [2:0]    port_state_out_0_1_2,
  output     [2:0]    port_state_out_0_1_3,
  output     [2:0]    port_state_out_0_1_4,
  output     [2:0]    port_state_out_0_1_5,
  output     [2:0]    port_state_out_0_1_6,
  output     [2:0]    port_state_out_0_1_7,
  output     [2:0]    port_state_out_0_2_0,
  output     [2:0]    port_state_out_0_2_1,
  output     [2:0]    port_state_out_0_2_2,
  output     [2:0]    port_state_out_0_2_3,
  output     [2:0]    port_state_out_0_2_4,
  output     [2:0]    port_state_out_0_2_5,
  output     [2:0]    port_state_out_0_2_6,
  output     [2:0]    port_state_out_0_2_7,
  output     [2:0]    port_state_out_0_3_0,
  output     [2:0]    port_state_out_0_3_1,
  output     [2:0]    port_state_out_0_3_2,
  output     [2:0]    port_state_out_0_3_3,
  output     [2:0]    port_state_out_0_3_4,
  output     [2:0]    port_state_out_0_3_5,
  output     [2:0]    port_state_out_0_3_6,
  output     [2:0]    port_state_out_0_3_7,
  output     [2:0]    port_state_out_1_0_0,
  output     [2:0]    port_state_out_1_0_1,
  output     [2:0]    port_state_out_1_0_2,
  output     [2:0]    port_state_out_1_0_3,
  output     [2:0]    port_state_out_1_0_4,
  output     [2:0]    port_state_out_1_0_5,
  output     [2:0]    port_state_out_1_0_6,
  output     [2:0]    port_state_out_1_0_7,
  output     [2:0]    port_state_out_1_1_0,
  output     [2:0]    port_state_out_1_1_1,
  output     [2:0]    port_state_out_1_1_2,
  output     [2:0]    port_state_out_1_1_3,
  output     [2:0]    port_state_out_1_1_4,
  output     [2:0]    port_state_out_1_1_5,
  output     [2:0]    port_state_out_1_1_6,
  output     [2:0]    port_state_out_1_1_7,
  output     [2:0]    port_state_out_1_2_0,
  output     [2:0]    port_state_out_1_2_1,
  output     [2:0]    port_state_out_1_2_2,
  output     [2:0]    port_state_out_1_2_3,
  output     [2:0]    port_state_out_1_2_4,
  output     [2:0]    port_state_out_1_2_5,
  output     [2:0]    port_state_out_1_2_6,
  output     [2:0]    port_state_out_1_2_7,
  output     [2:0]    port_state_out_1_3_0,
  output     [2:0]    port_state_out_1_3_1,
  output     [2:0]    port_state_out_1_3_2,
  output     [2:0]    port_state_out_1_3_3,
  output     [2:0]    port_state_out_1_3_4,
  output     [2:0]    port_state_out_1_3_5,
  output     [2:0]    port_state_out_1_3_6,
  output     [2:0]    port_state_out_1_3_7,
  output     [2:0]    port_state_out_2_0_0,
  output     [2:0]    port_state_out_2_0_1,
  output     [2:0]    port_state_out_2_0_2,
  output     [2:0]    port_state_out_2_0_3,
  output     [2:0]    port_state_out_2_0_4,
  output     [2:0]    port_state_out_2_0_5,
  output     [2:0]    port_state_out_2_0_6,
  output     [2:0]    port_state_out_2_0_7,
  output     [2:0]    port_state_out_2_1_0,
  output     [2:0]    port_state_out_2_1_1,
  output     [2:0]    port_state_out_2_1_2,
  output     [2:0]    port_state_out_2_1_3,
  output     [2:0]    port_state_out_2_1_4,
  output     [2:0]    port_state_out_2_1_5,
  output     [2:0]    port_state_out_2_1_6,
  output     [2:0]    port_state_out_2_1_7,
  output     [2:0]    port_state_out_2_2_0,
  output     [2:0]    port_state_out_2_2_1,
  output     [2:0]    port_state_out_2_2_2,
  output     [2:0]    port_state_out_2_2_3,
  output     [2:0]    port_state_out_2_2_4,
  output     [2:0]    port_state_out_2_2_5,
  output     [2:0]    port_state_out_2_2_6,
  output     [2:0]    port_state_out_2_2_7,
  output     [2:0]    port_state_out_2_3_0,
  output     [2:0]    port_state_out_2_3_1,
  output     [2:0]    port_state_out_2_3_2,
  output     [2:0]    port_state_out_2_3_3,
  output     [2:0]    port_state_out_2_3_4,
  output     [2:0]    port_state_out_2_3_5,
  output     [2:0]    port_state_out_2_3_6,
  output     [2:0]    port_state_out_2_3_7,
  output     [2:0]    port_state_out_3_0_0,
  output     [2:0]    port_state_out_3_0_1,
  output     [2:0]    port_state_out_3_0_2,
  output     [2:0]    port_state_out_3_0_3,
  output     [2:0]    port_state_out_3_0_4,
  output     [2:0]    port_state_out_3_0_5,
  output     [2:0]    port_state_out_3_0_6,
  output     [2:0]    port_state_out_3_0_7,
  output     [2:0]    port_state_out_3_1_0,
  output     [2:0]    port_state_out_3_1_1,
  output     [2:0]    port_state_out_3_1_2,
  output     [2:0]    port_state_out_3_1_3,
  output     [2:0]    port_state_out_3_1_4,
  output     [2:0]    port_state_out_3_1_5,
  output     [2:0]    port_state_out_3_1_6,
  output     [2:0]    port_state_out_3_1_7,
  output     [2:0]    port_state_out_3_2_0,
  output     [2:0]    port_state_out_3_2_1,
  output     [2:0]    port_state_out_3_2_2,
  output     [2:0]    port_state_out_3_2_3,
  output     [2:0]    port_state_out_3_2_4,
  output     [2:0]    port_state_out_3_2_5,
  output     [2:0]    port_state_out_3_2_6,
  output     [2:0]    port_state_out_3_2_7,
  output     [2:0]    port_state_out_3_3_0,
  output     [2:0]    port_state_out_3_3_1,
  output     [2:0]    port_state_out_3_3_2,
  output     [2:0]    port_state_out_3_3_3,
  output     [2:0]    port_state_out_3_3_4,
  output     [2:0]    port_state_out_3_3_5,
  output     [2:0]    port_state_out_3_3_6,
  output     [2:0]    port_state_out_3_3_7,
  output     [2:0]    port_state_out_4_0_0,
  output     [2:0]    port_state_out_4_0_1,
  output     [2:0]    port_state_out_4_0_2,
  output     [2:0]    port_state_out_4_0_3,
  output     [2:0]    port_state_out_4_0_4,
  output     [2:0]    port_state_out_4_0_5,
  output     [2:0]    port_state_out_4_0_6,
  output     [2:0]    port_state_out_4_0_7,
  output     [2:0]    port_state_out_4_1_0,
  output     [2:0]    port_state_out_4_1_1,
  output     [2:0]    port_state_out_4_1_2,
  output     [2:0]    port_state_out_4_1_3,
  output     [2:0]    port_state_out_4_1_4,
  output     [2:0]    port_state_out_4_1_5,
  output     [2:0]    port_state_out_4_1_6,
  output     [2:0]    port_state_out_4_1_7,
  output     [2:0]    port_state_out_4_2_0,
  output     [2:0]    port_state_out_4_2_1,
  output     [2:0]    port_state_out_4_2_2,
  output     [2:0]    port_state_out_4_2_3,
  output     [2:0]    port_state_out_4_2_4,
  output     [2:0]    port_state_out_4_2_5,
  output     [2:0]    port_state_out_4_2_6,
  output     [2:0]    port_state_out_4_2_7,
  output     [2:0]    port_state_out_4_3_0,
  output     [2:0]    port_state_out_4_3_1,
  output     [2:0]    port_state_out_4_3_2,
  output     [2:0]    port_state_out_4_3_3,
  output     [2:0]    port_state_out_4_3_4,
  output     [2:0]    port_state_out_4_3_5,
  output     [2:0]    port_state_out_4_3_6,
  output     [2:0]    port_state_out_4_3_7,
  output     [2:0]    port_state_out_5_0_0,
  output     [2:0]    port_state_out_5_0_1,
  output     [2:0]    port_state_out_5_0_2,
  output     [2:0]    port_state_out_5_0_3,
  output     [2:0]    port_state_out_5_0_4,
  output     [2:0]    port_state_out_5_0_5,
  output     [2:0]    port_state_out_5_0_6,
  output     [2:0]    port_state_out_5_0_7,
  output     [2:0]    port_state_out_5_1_0,
  output     [2:0]    port_state_out_5_1_1,
  output     [2:0]    port_state_out_5_1_2,
  output     [2:0]    port_state_out_5_1_3,
  output     [2:0]    port_state_out_5_1_4,
  output     [2:0]    port_state_out_5_1_5,
  output     [2:0]    port_state_out_5_1_6,
  output     [2:0]    port_state_out_5_1_7,
  output     [2:0]    port_state_out_5_2_0,
  output     [2:0]    port_state_out_5_2_1,
  output     [2:0]    port_state_out_5_2_2,
  output     [2:0]    port_state_out_5_2_3,
  output     [2:0]    port_state_out_5_2_4,
  output     [2:0]    port_state_out_5_2_5,
  output     [2:0]    port_state_out_5_2_6,
  output     [2:0]    port_state_out_5_2_7,
  output     [2:0]    port_state_out_5_3_0,
  output     [2:0]    port_state_out_5_3_1,
  output     [2:0]    port_state_out_5_3_2,
  output     [2:0]    port_state_out_5_3_3,
  output     [2:0]    port_state_out_5_3_4,
  output     [2:0]    port_state_out_5_3_5,
  output     [2:0]    port_state_out_5_3_6,
  output     [2:0]    port_state_out_5_3_7,
  output     [2:0]    port_state_out_6_0_0,
  output     [2:0]    port_state_out_6_0_1,
  output     [2:0]    port_state_out_6_0_2,
  output     [2:0]    port_state_out_6_0_3,
  output     [2:0]    port_state_out_6_0_4,
  output     [2:0]    port_state_out_6_0_5,
  output     [2:0]    port_state_out_6_0_6,
  output     [2:0]    port_state_out_6_0_7,
  output     [2:0]    port_state_out_6_1_0,
  output     [2:0]    port_state_out_6_1_1,
  output     [2:0]    port_state_out_6_1_2,
  output     [2:0]    port_state_out_6_1_3,
  output     [2:0]    port_state_out_6_1_4,
  output     [2:0]    port_state_out_6_1_5,
  output     [2:0]    port_state_out_6_1_6,
  output     [2:0]    port_state_out_6_1_7,
  output     [2:0]    port_state_out_6_2_0,
  output     [2:0]    port_state_out_6_2_1,
  output     [2:0]    port_state_out_6_2_2,
  output     [2:0]    port_state_out_6_2_3,
  output     [2:0]    port_state_out_6_2_4,
  output     [2:0]    port_state_out_6_2_5,
  output     [2:0]    port_state_out_6_2_6,
  output     [2:0]    port_state_out_6_2_7,
  output     [2:0]    port_state_out_6_3_0,
  output     [2:0]    port_state_out_6_3_1,
  output     [2:0]    port_state_out_6_3_2,
  output     [2:0]    port_state_out_6_3_3,
  output     [2:0]    port_state_out_6_3_4,
  output     [2:0]    port_state_out_6_3_5,
  output     [2:0]    port_state_out_6_3_6,
  output     [2:0]    port_state_out_6_3_7,
  output     [2:0]    port_state_out_7_0_0,
  output     [2:0]    port_state_out_7_0_1,
  output     [2:0]    port_state_out_7_0_2,
  output     [2:0]    port_state_out_7_0_3,
  output     [2:0]    port_state_out_7_0_4,
  output     [2:0]    port_state_out_7_0_5,
  output     [2:0]    port_state_out_7_0_6,
  output     [2:0]    port_state_out_7_0_7,
  output     [2:0]    port_state_out_7_1_0,
  output     [2:0]    port_state_out_7_1_1,
  output     [2:0]    port_state_out_7_1_2,
  output     [2:0]    port_state_out_7_1_3,
  output     [2:0]    port_state_out_7_1_4,
  output     [2:0]    port_state_out_7_1_5,
  output     [2:0]    port_state_out_7_1_6,
  output     [2:0]    port_state_out_7_1_7,
  output     [2:0]    port_state_out_7_2_0,
  output     [2:0]    port_state_out_7_2_1,
  output     [2:0]    port_state_out_7_2_2,
  output     [2:0]    port_state_out_7_2_3,
  output     [2:0]    port_state_out_7_2_4,
  output     [2:0]    port_state_out_7_2_5,
  output     [2:0]    port_state_out_7_2_6,
  output     [2:0]    port_state_out_7_2_7,
  output     [2:0]    port_state_out_7_3_0,
  output     [2:0]    port_state_out_7_3_1,
  output     [2:0]    port_state_out_7_3_2,
  output     [2:0]    port_state_out_7_3_3,
  output     [2:0]    port_state_out_7_3_4,
  output     [2:0]    port_state_out_7_3_5,
  output     [2:0]    port_state_out_7_3_6,
  output     [2:0]    port_state_out_7_3_7,
  output     [2:0]    port_state_out_8_0_0,
  output     [2:0]    port_state_out_8_0_1,
  output     [2:0]    port_state_out_8_0_2,
  output     [2:0]    port_state_out_8_0_3,
  output     [2:0]    port_state_out_8_0_4,
  output     [2:0]    port_state_out_8_0_5,
  output     [2:0]    port_state_out_8_0_6,
  output     [2:0]    port_state_out_8_0_7,
  output     [2:0]    port_state_out_8_1_0,
  output     [2:0]    port_state_out_8_1_1,
  output     [2:0]    port_state_out_8_1_2,
  output     [2:0]    port_state_out_8_1_3,
  output     [2:0]    port_state_out_8_1_4,
  output     [2:0]    port_state_out_8_1_5,
  output     [2:0]    port_state_out_8_1_6,
  output     [2:0]    port_state_out_8_1_7,
  output     [2:0]    port_state_out_8_2_0,
  output     [2:0]    port_state_out_8_2_1,
  output     [2:0]    port_state_out_8_2_2,
  output     [2:0]    port_state_out_8_2_3,
  output     [2:0]    port_state_out_8_2_4,
  output     [2:0]    port_state_out_8_2_5,
  output     [2:0]    port_state_out_8_2_6,
  output     [2:0]    port_state_out_8_2_7,
  output     [2:0]    port_state_out_8_3_0,
  output     [2:0]    port_state_out_8_3_1,
  output     [2:0]    port_state_out_8_3_2,
  output     [2:0]    port_state_out_8_3_3,
  output     [2:0]    port_state_out_8_3_4,
  output     [2:0]    port_state_out_8_3_5,
  output     [2:0]    port_state_out_8_3_6,
  output     [2:0]    port_state_out_8_3_7,
  output     [2:0]    port_state_out_9_0_0,
  output     [2:0]    port_state_out_9_0_1,
  output     [2:0]    port_state_out_9_0_2,
  output     [2:0]    port_state_out_9_0_3,
  output     [2:0]    port_state_out_9_0_4,
  output     [2:0]    port_state_out_9_0_5,
  output     [2:0]    port_state_out_9_0_6,
  output     [2:0]    port_state_out_9_0_7,
  output     [2:0]    port_state_out_9_1_0,
  output     [2:0]    port_state_out_9_1_1,
  output     [2:0]    port_state_out_9_1_2,
  output     [2:0]    port_state_out_9_1_3,
  output     [2:0]    port_state_out_9_1_4,
  output     [2:0]    port_state_out_9_1_5,
  output     [2:0]    port_state_out_9_1_6,
  output     [2:0]    port_state_out_9_1_7,
  output     [2:0]    port_state_out_9_2_0,
  output     [2:0]    port_state_out_9_2_1,
  output     [2:0]    port_state_out_9_2_2,
  output     [2:0]    port_state_out_9_2_3,
  output     [2:0]    port_state_out_9_2_4,
  output     [2:0]    port_state_out_9_2_5,
  output     [2:0]    port_state_out_9_2_6,
  output     [2:0]    port_state_out_9_2_7,
  output     [2:0]    port_state_out_9_3_0,
  output     [2:0]    port_state_out_9_3_1,
  output     [2:0]    port_state_out_9_3_2,
  output     [2:0]    port_state_out_9_3_3,
  output     [2:0]    port_state_out_9_3_4,
  output     [2:0]    port_state_out_9_3_5,
  output     [2:0]    port_state_out_9_3_6,
  output     [2:0]    port_state_out_9_3_7,
  output     [2:0]    port_state_out_10_0_0,
  output     [2:0]    port_state_out_10_0_1,
  output     [2:0]    port_state_out_10_0_2,
  output     [2:0]    port_state_out_10_0_3,
  output     [2:0]    port_state_out_10_0_4,
  output     [2:0]    port_state_out_10_0_5,
  output     [2:0]    port_state_out_10_0_6,
  output     [2:0]    port_state_out_10_0_7,
  output     [2:0]    port_state_out_10_1_0,
  output     [2:0]    port_state_out_10_1_1,
  output     [2:0]    port_state_out_10_1_2,
  output     [2:0]    port_state_out_10_1_3,
  output     [2:0]    port_state_out_10_1_4,
  output     [2:0]    port_state_out_10_1_5,
  output     [2:0]    port_state_out_10_1_6,
  output     [2:0]    port_state_out_10_1_7,
  output     [2:0]    port_state_out_10_2_0,
  output     [2:0]    port_state_out_10_2_1,
  output     [2:0]    port_state_out_10_2_2,
  output     [2:0]    port_state_out_10_2_3,
  output     [2:0]    port_state_out_10_2_4,
  output     [2:0]    port_state_out_10_2_5,
  output     [2:0]    port_state_out_10_2_6,
  output     [2:0]    port_state_out_10_2_7,
  output     [2:0]    port_state_out_10_3_0,
  output     [2:0]    port_state_out_10_3_1,
  output     [2:0]    port_state_out_10_3_2,
  output     [2:0]    port_state_out_10_3_3,
  output     [2:0]    port_state_out_10_3_4,
  output     [2:0]    port_state_out_10_3_5,
  output     [2:0]    port_state_out_10_3_6,
  output     [2:0]    port_state_out_10_3_7,
  output     [2:0]    port_state_out_11_0_0,
  output     [2:0]    port_state_out_11_0_1,
  output     [2:0]    port_state_out_11_0_2,
  output     [2:0]    port_state_out_11_0_3,
  output     [2:0]    port_state_out_11_0_4,
  output     [2:0]    port_state_out_11_0_5,
  output     [2:0]    port_state_out_11_0_6,
  output     [2:0]    port_state_out_11_0_7,
  output     [2:0]    port_state_out_11_1_0,
  output     [2:0]    port_state_out_11_1_1,
  output     [2:0]    port_state_out_11_1_2,
  output     [2:0]    port_state_out_11_1_3,
  output     [2:0]    port_state_out_11_1_4,
  output     [2:0]    port_state_out_11_1_5,
  output     [2:0]    port_state_out_11_1_6,
  output     [2:0]    port_state_out_11_1_7,
  output     [2:0]    port_state_out_11_2_0,
  output     [2:0]    port_state_out_11_2_1,
  output     [2:0]    port_state_out_11_2_2,
  output     [2:0]    port_state_out_11_2_3,
  output     [2:0]    port_state_out_11_2_4,
  output     [2:0]    port_state_out_11_2_5,
  output     [2:0]    port_state_out_11_2_6,
  output     [2:0]    port_state_out_11_2_7,
  output     [2:0]    port_state_out_11_3_0,
  output     [2:0]    port_state_out_11_3_1,
  output     [2:0]    port_state_out_11_3_2,
  output     [2:0]    port_state_out_11_3_3,
  output     [2:0]    port_state_out_11_3_4,
  output     [2:0]    port_state_out_11_3_5,
  output     [2:0]    port_state_out_11_3_6,
  output     [2:0]    port_state_out_11_3_7,
  output     [2:0]    port_state_out_12_0_0,
  output     [2:0]    port_state_out_12_0_1,
  output     [2:0]    port_state_out_12_0_2,
  output     [2:0]    port_state_out_12_0_3,
  output     [2:0]    port_state_out_12_0_4,
  output     [2:0]    port_state_out_12_0_5,
  output     [2:0]    port_state_out_12_0_6,
  output     [2:0]    port_state_out_12_0_7,
  output     [2:0]    port_state_out_12_1_0,
  output     [2:0]    port_state_out_12_1_1,
  output     [2:0]    port_state_out_12_1_2,
  output     [2:0]    port_state_out_12_1_3,
  output     [2:0]    port_state_out_12_1_4,
  output     [2:0]    port_state_out_12_1_5,
  output     [2:0]    port_state_out_12_1_6,
  output     [2:0]    port_state_out_12_1_7,
  output     [2:0]    port_state_out_12_2_0,
  output     [2:0]    port_state_out_12_2_1,
  output     [2:0]    port_state_out_12_2_2,
  output     [2:0]    port_state_out_12_2_3,
  output     [2:0]    port_state_out_12_2_4,
  output     [2:0]    port_state_out_12_2_5,
  output     [2:0]    port_state_out_12_2_6,
  output     [2:0]    port_state_out_12_2_7,
  output     [2:0]    port_state_out_12_3_0,
  output     [2:0]    port_state_out_12_3_1,
  output     [2:0]    port_state_out_12_3_2,
  output     [2:0]    port_state_out_12_3_3,
  output     [2:0]    port_state_out_12_3_4,
  output     [2:0]    port_state_out_12_3_5,
  output     [2:0]    port_state_out_12_3_6,
  output     [2:0]    port_state_out_12_3_7,
  output     [2:0]    port_state_out_13_0_0,
  output     [2:0]    port_state_out_13_0_1,
  output     [2:0]    port_state_out_13_0_2,
  output     [2:0]    port_state_out_13_0_3,
  output     [2:0]    port_state_out_13_0_4,
  output     [2:0]    port_state_out_13_0_5,
  output     [2:0]    port_state_out_13_0_6,
  output     [2:0]    port_state_out_13_0_7,
  output     [2:0]    port_state_out_13_1_0,
  output     [2:0]    port_state_out_13_1_1,
  output     [2:0]    port_state_out_13_1_2,
  output     [2:0]    port_state_out_13_1_3,
  output     [2:0]    port_state_out_13_1_4,
  output     [2:0]    port_state_out_13_1_5,
  output     [2:0]    port_state_out_13_1_6,
  output     [2:0]    port_state_out_13_1_7,
  output     [2:0]    port_state_out_13_2_0,
  output     [2:0]    port_state_out_13_2_1,
  output     [2:0]    port_state_out_13_2_2,
  output     [2:0]    port_state_out_13_2_3,
  output     [2:0]    port_state_out_13_2_4,
  output     [2:0]    port_state_out_13_2_5,
  output     [2:0]    port_state_out_13_2_6,
  output     [2:0]    port_state_out_13_2_7,
  output     [2:0]    port_state_out_13_3_0,
  output     [2:0]    port_state_out_13_3_1,
  output     [2:0]    port_state_out_13_3_2,
  output     [2:0]    port_state_out_13_3_3,
  output     [2:0]    port_state_out_13_3_4,
  output     [2:0]    port_state_out_13_3_5,
  output     [2:0]    port_state_out_13_3_6,
  output     [2:0]    port_state_out_13_3_7,
  output     [2:0]    port_state_out_14_0_0,
  output     [2:0]    port_state_out_14_0_1,
  output     [2:0]    port_state_out_14_0_2,
  output     [2:0]    port_state_out_14_0_3,
  output     [2:0]    port_state_out_14_0_4,
  output     [2:0]    port_state_out_14_0_5,
  output     [2:0]    port_state_out_14_0_6,
  output     [2:0]    port_state_out_14_0_7,
  output     [2:0]    port_state_out_14_1_0,
  output     [2:0]    port_state_out_14_1_1,
  output     [2:0]    port_state_out_14_1_2,
  output     [2:0]    port_state_out_14_1_3,
  output     [2:0]    port_state_out_14_1_4,
  output     [2:0]    port_state_out_14_1_5,
  output     [2:0]    port_state_out_14_1_6,
  output     [2:0]    port_state_out_14_1_7,
  output     [2:0]    port_state_out_14_2_0,
  output     [2:0]    port_state_out_14_2_1,
  output     [2:0]    port_state_out_14_2_2,
  output     [2:0]    port_state_out_14_2_3,
  output     [2:0]    port_state_out_14_2_4,
  output     [2:0]    port_state_out_14_2_5,
  output     [2:0]    port_state_out_14_2_6,
  output     [2:0]    port_state_out_14_2_7,
  output     [2:0]    port_state_out_14_3_0,
  output     [2:0]    port_state_out_14_3_1,
  output     [2:0]    port_state_out_14_3_2,
  output     [2:0]    port_state_out_14_3_3,
  output     [2:0]    port_state_out_14_3_4,
  output     [2:0]    port_state_out_14_3_5,
  output     [2:0]    port_state_out_14_3_6,
  output     [2:0]    port_state_out_14_3_7,
  output     [2:0]    port_state_out_15_0_0,
  output     [2:0]    port_state_out_15_0_1,
  output     [2:0]    port_state_out_15_0_2,
  output     [2:0]    port_state_out_15_0_3,
  output     [2:0]    port_state_out_15_0_4,
  output     [2:0]    port_state_out_15_0_5,
  output     [2:0]    port_state_out_15_0_6,
  output     [2:0]    port_state_out_15_0_7,
  output     [2:0]    port_state_out_15_1_0,
  output     [2:0]    port_state_out_15_1_1,
  output     [2:0]    port_state_out_15_1_2,
  output     [2:0]    port_state_out_15_1_3,
  output     [2:0]    port_state_out_15_1_4,
  output     [2:0]    port_state_out_15_1_5,
  output     [2:0]    port_state_out_15_1_6,
  output     [2:0]    port_state_out_15_1_7,
  output     [2:0]    port_state_out_15_2_0,
  output     [2:0]    port_state_out_15_2_1,
  output     [2:0]    port_state_out_15_2_2,
  output     [2:0]    port_state_out_15_2_3,
  output     [2:0]    port_state_out_15_2_4,
  output     [2:0]    port_state_out_15_2_5,
  output     [2:0]    port_state_out_15_2_6,
  output     [2:0]    port_state_out_15_2_7,
  output     [2:0]    port_state_out_15_3_0,
  output     [2:0]    port_state_out_15_3_1,
  output     [2:0]    port_state_out_15_3_2,
  output     [2:0]    port_state_out_15_3_3,
  output     [2:0]    port_state_out_15_3_4,
  output     [2:0]    port_state_out_15_3_5,
  output     [2:0]    port_state_out_15_3_6,
  output     [2:0]    port_state_out_15_3_7
);

  wire       [2:0]    mul2_64_port_byte_out_0;
  wire       [2:0]    mul2_64_port_byte_out_1;
  wire       [2:0]    mul2_64_port_byte_out_2;
  wire       [2:0]    mul2_64_port_byte_out_3;
  wire       [2:0]    mul2_64_port_byte_out_4;
  wire       [2:0]    mul2_64_port_byte_out_5;
  wire       [2:0]    mul2_64_port_byte_out_6;
  wire       [2:0]    mul2_64_port_byte_out_7;
  wire       [2:0]    mul3_64_port_byte_out_0;
  wire       [2:0]    mul3_64_port_byte_out_1;
  wire       [2:0]    mul3_64_port_byte_out_2;
  wire       [2:0]    mul3_64_port_byte_out_3;
  wire       [2:0]    mul3_64_port_byte_out_4;
  wire       [2:0]    mul3_64_port_byte_out_5;
  wire       [2:0]    mul3_64_port_byte_out_6;
  wire       [2:0]    mul3_64_port_byte_out_7;
  wire       [2:0]    mul2_65_port_byte_out_0;
  wire       [2:0]    mul2_65_port_byte_out_1;
  wire       [2:0]    mul2_65_port_byte_out_2;
  wire       [2:0]    mul2_65_port_byte_out_3;
  wire       [2:0]    mul2_65_port_byte_out_4;
  wire       [2:0]    mul2_65_port_byte_out_5;
  wire       [2:0]    mul2_65_port_byte_out_6;
  wire       [2:0]    mul2_65_port_byte_out_7;
  wire       [2:0]    mul3_65_port_byte_out_0;
  wire       [2:0]    mul3_65_port_byte_out_1;
  wire       [2:0]    mul3_65_port_byte_out_2;
  wire       [2:0]    mul3_65_port_byte_out_3;
  wire       [2:0]    mul3_65_port_byte_out_4;
  wire       [2:0]    mul3_65_port_byte_out_5;
  wire       [2:0]    mul3_65_port_byte_out_6;
  wire       [2:0]    mul3_65_port_byte_out_7;
  wire       [2:0]    mul2_66_port_byte_out_0;
  wire       [2:0]    mul2_66_port_byte_out_1;
  wire       [2:0]    mul2_66_port_byte_out_2;
  wire       [2:0]    mul2_66_port_byte_out_3;
  wire       [2:0]    mul2_66_port_byte_out_4;
  wire       [2:0]    mul2_66_port_byte_out_5;
  wire       [2:0]    mul2_66_port_byte_out_6;
  wire       [2:0]    mul2_66_port_byte_out_7;
  wire       [2:0]    mul3_66_port_byte_out_0;
  wire       [2:0]    mul3_66_port_byte_out_1;
  wire       [2:0]    mul3_66_port_byte_out_2;
  wire       [2:0]    mul3_66_port_byte_out_3;
  wire       [2:0]    mul3_66_port_byte_out_4;
  wire       [2:0]    mul3_66_port_byte_out_5;
  wire       [2:0]    mul3_66_port_byte_out_6;
  wire       [2:0]    mul3_66_port_byte_out_7;
  wire       [2:0]    mul2_67_port_byte_out_0;
  wire       [2:0]    mul2_67_port_byte_out_1;
  wire       [2:0]    mul2_67_port_byte_out_2;
  wire       [2:0]    mul2_67_port_byte_out_3;
  wire       [2:0]    mul2_67_port_byte_out_4;
  wire       [2:0]    mul2_67_port_byte_out_5;
  wire       [2:0]    mul2_67_port_byte_out_6;
  wire       [2:0]    mul2_67_port_byte_out_7;
  wire       [2:0]    mul3_67_port_byte_out_0;
  wire       [2:0]    mul3_67_port_byte_out_1;
  wire       [2:0]    mul3_67_port_byte_out_2;
  wire       [2:0]    mul3_67_port_byte_out_3;
  wire       [2:0]    mul3_67_port_byte_out_4;
  wire       [2:0]    mul3_67_port_byte_out_5;
  wire       [2:0]    mul3_67_port_byte_out_6;
  wire       [2:0]    mul3_67_port_byte_out_7;
  wire       [2:0]    mul2_68_port_byte_out_0;
  wire       [2:0]    mul2_68_port_byte_out_1;
  wire       [2:0]    mul2_68_port_byte_out_2;
  wire       [2:0]    mul2_68_port_byte_out_3;
  wire       [2:0]    mul2_68_port_byte_out_4;
  wire       [2:0]    mul2_68_port_byte_out_5;
  wire       [2:0]    mul2_68_port_byte_out_6;
  wire       [2:0]    mul2_68_port_byte_out_7;
  wire       [2:0]    mul3_68_port_byte_out_0;
  wire       [2:0]    mul3_68_port_byte_out_1;
  wire       [2:0]    mul3_68_port_byte_out_2;
  wire       [2:0]    mul3_68_port_byte_out_3;
  wire       [2:0]    mul3_68_port_byte_out_4;
  wire       [2:0]    mul3_68_port_byte_out_5;
  wire       [2:0]    mul3_68_port_byte_out_6;
  wire       [2:0]    mul3_68_port_byte_out_7;
  wire       [2:0]    mul2_69_port_byte_out_0;
  wire       [2:0]    mul2_69_port_byte_out_1;
  wire       [2:0]    mul2_69_port_byte_out_2;
  wire       [2:0]    mul2_69_port_byte_out_3;
  wire       [2:0]    mul2_69_port_byte_out_4;
  wire       [2:0]    mul2_69_port_byte_out_5;
  wire       [2:0]    mul2_69_port_byte_out_6;
  wire       [2:0]    mul2_69_port_byte_out_7;
  wire       [2:0]    mul3_69_port_byte_out_0;
  wire       [2:0]    mul3_69_port_byte_out_1;
  wire       [2:0]    mul3_69_port_byte_out_2;
  wire       [2:0]    mul3_69_port_byte_out_3;
  wire       [2:0]    mul3_69_port_byte_out_4;
  wire       [2:0]    mul3_69_port_byte_out_5;
  wire       [2:0]    mul3_69_port_byte_out_6;
  wire       [2:0]    mul3_69_port_byte_out_7;
  wire       [2:0]    mul2_70_port_byte_out_0;
  wire       [2:0]    mul2_70_port_byte_out_1;
  wire       [2:0]    mul2_70_port_byte_out_2;
  wire       [2:0]    mul2_70_port_byte_out_3;
  wire       [2:0]    mul2_70_port_byte_out_4;
  wire       [2:0]    mul2_70_port_byte_out_5;
  wire       [2:0]    mul2_70_port_byte_out_6;
  wire       [2:0]    mul2_70_port_byte_out_7;
  wire       [2:0]    mul3_70_port_byte_out_0;
  wire       [2:0]    mul3_70_port_byte_out_1;
  wire       [2:0]    mul3_70_port_byte_out_2;
  wire       [2:0]    mul3_70_port_byte_out_3;
  wire       [2:0]    mul3_70_port_byte_out_4;
  wire       [2:0]    mul3_70_port_byte_out_5;
  wire       [2:0]    mul3_70_port_byte_out_6;
  wire       [2:0]    mul3_70_port_byte_out_7;
  wire       [2:0]    mul2_71_port_byte_out_0;
  wire       [2:0]    mul2_71_port_byte_out_1;
  wire       [2:0]    mul2_71_port_byte_out_2;
  wire       [2:0]    mul2_71_port_byte_out_3;
  wire       [2:0]    mul2_71_port_byte_out_4;
  wire       [2:0]    mul2_71_port_byte_out_5;
  wire       [2:0]    mul2_71_port_byte_out_6;
  wire       [2:0]    mul2_71_port_byte_out_7;
  wire       [2:0]    mul3_71_port_byte_out_0;
  wire       [2:0]    mul3_71_port_byte_out_1;
  wire       [2:0]    mul3_71_port_byte_out_2;
  wire       [2:0]    mul3_71_port_byte_out_3;
  wire       [2:0]    mul3_71_port_byte_out_4;
  wire       [2:0]    mul3_71_port_byte_out_5;
  wire       [2:0]    mul3_71_port_byte_out_6;
  wire       [2:0]    mul3_71_port_byte_out_7;
  wire       [2:0]    mul2_72_port_byte_out_0;
  wire       [2:0]    mul2_72_port_byte_out_1;
  wire       [2:0]    mul2_72_port_byte_out_2;
  wire       [2:0]    mul2_72_port_byte_out_3;
  wire       [2:0]    mul2_72_port_byte_out_4;
  wire       [2:0]    mul2_72_port_byte_out_5;
  wire       [2:0]    mul2_72_port_byte_out_6;
  wire       [2:0]    mul2_72_port_byte_out_7;
  wire       [2:0]    mul3_72_port_byte_out_0;
  wire       [2:0]    mul3_72_port_byte_out_1;
  wire       [2:0]    mul3_72_port_byte_out_2;
  wire       [2:0]    mul3_72_port_byte_out_3;
  wire       [2:0]    mul3_72_port_byte_out_4;
  wire       [2:0]    mul3_72_port_byte_out_5;
  wire       [2:0]    mul3_72_port_byte_out_6;
  wire       [2:0]    mul3_72_port_byte_out_7;
  wire       [2:0]    mul2_73_port_byte_out_0;
  wire       [2:0]    mul2_73_port_byte_out_1;
  wire       [2:0]    mul2_73_port_byte_out_2;
  wire       [2:0]    mul2_73_port_byte_out_3;
  wire       [2:0]    mul2_73_port_byte_out_4;
  wire       [2:0]    mul2_73_port_byte_out_5;
  wire       [2:0]    mul2_73_port_byte_out_6;
  wire       [2:0]    mul2_73_port_byte_out_7;
  wire       [2:0]    mul3_73_port_byte_out_0;
  wire       [2:0]    mul3_73_port_byte_out_1;
  wire       [2:0]    mul3_73_port_byte_out_2;
  wire       [2:0]    mul3_73_port_byte_out_3;
  wire       [2:0]    mul3_73_port_byte_out_4;
  wire       [2:0]    mul3_73_port_byte_out_5;
  wire       [2:0]    mul3_73_port_byte_out_6;
  wire       [2:0]    mul3_73_port_byte_out_7;
  wire       [2:0]    mul2_74_port_byte_out_0;
  wire       [2:0]    mul2_74_port_byte_out_1;
  wire       [2:0]    mul2_74_port_byte_out_2;
  wire       [2:0]    mul2_74_port_byte_out_3;
  wire       [2:0]    mul2_74_port_byte_out_4;
  wire       [2:0]    mul2_74_port_byte_out_5;
  wire       [2:0]    mul2_74_port_byte_out_6;
  wire       [2:0]    mul2_74_port_byte_out_7;
  wire       [2:0]    mul3_74_port_byte_out_0;
  wire       [2:0]    mul3_74_port_byte_out_1;
  wire       [2:0]    mul3_74_port_byte_out_2;
  wire       [2:0]    mul3_74_port_byte_out_3;
  wire       [2:0]    mul3_74_port_byte_out_4;
  wire       [2:0]    mul3_74_port_byte_out_5;
  wire       [2:0]    mul3_74_port_byte_out_6;
  wire       [2:0]    mul3_74_port_byte_out_7;
  wire       [2:0]    mul2_75_port_byte_out_0;
  wire       [2:0]    mul2_75_port_byte_out_1;
  wire       [2:0]    mul2_75_port_byte_out_2;
  wire       [2:0]    mul2_75_port_byte_out_3;
  wire       [2:0]    mul2_75_port_byte_out_4;
  wire       [2:0]    mul2_75_port_byte_out_5;
  wire       [2:0]    mul2_75_port_byte_out_6;
  wire       [2:0]    mul2_75_port_byte_out_7;
  wire       [2:0]    mul3_75_port_byte_out_0;
  wire       [2:0]    mul3_75_port_byte_out_1;
  wire       [2:0]    mul3_75_port_byte_out_2;
  wire       [2:0]    mul3_75_port_byte_out_3;
  wire       [2:0]    mul3_75_port_byte_out_4;
  wire       [2:0]    mul3_75_port_byte_out_5;
  wire       [2:0]    mul3_75_port_byte_out_6;
  wire       [2:0]    mul3_75_port_byte_out_7;
  wire       [2:0]    mul2_76_port_byte_out_0;
  wire       [2:0]    mul2_76_port_byte_out_1;
  wire       [2:0]    mul2_76_port_byte_out_2;
  wire       [2:0]    mul2_76_port_byte_out_3;
  wire       [2:0]    mul2_76_port_byte_out_4;
  wire       [2:0]    mul2_76_port_byte_out_5;
  wire       [2:0]    mul2_76_port_byte_out_6;
  wire       [2:0]    mul2_76_port_byte_out_7;
  wire       [2:0]    mul3_76_port_byte_out_0;
  wire       [2:0]    mul3_76_port_byte_out_1;
  wire       [2:0]    mul3_76_port_byte_out_2;
  wire       [2:0]    mul3_76_port_byte_out_3;
  wire       [2:0]    mul3_76_port_byte_out_4;
  wire       [2:0]    mul3_76_port_byte_out_5;
  wire       [2:0]    mul3_76_port_byte_out_6;
  wire       [2:0]    mul3_76_port_byte_out_7;
  wire       [2:0]    mul2_77_port_byte_out_0;
  wire       [2:0]    mul2_77_port_byte_out_1;
  wire       [2:0]    mul2_77_port_byte_out_2;
  wire       [2:0]    mul2_77_port_byte_out_3;
  wire       [2:0]    mul2_77_port_byte_out_4;
  wire       [2:0]    mul2_77_port_byte_out_5;
  wire       [2:0]    mul2_77_port_byte_out_6;
  wire       [2:0]    mul2_77_port_byte_out_7;
  wire       [2:0]    mul3_77_port_byte_out_0;
  wire       [2:0]    mul3_77_port_byte_out_1;
  wire       [2:0]    mul3_77_port_byte_out_2;
  wire       [2:0]    mul3_77_port_byte_out_3;
  wire       [2:0]    mul3_77_port_byte_out_4;
  wire       [2:0]    mul3_77_port_byte_out_5;
  wire       [2:0]    mul3_77_port_byte_out_6;
  wire       [2:0]    mul3_77_port_byte_out_7;
  wire       [2:0]    mul2_78_port_byte_out_0;
  wire       [2:0]    mul2_78_port_byte_out_1;
  wire       [2:0]    mul2_78_port_byte_out_2;
  wire       [2:0]    mul2_78_port_byte_out_3;
  wire       [2:0]    mul2_78_port_byte_out_4;
  wire       [2:0]    mul2_78_port_byte_out_5;
  wire       [2:0]    mul2_78_port_byte_out_6;
  wire       [2:0]    mul2_78_port_byte_out_7;
  wire       [2:0]    mul3_78_port_byte_out_0;
  wire       [2:0]    mul3_78_port_byte_out_1;
  wire       [2:0]    mul3_78_port_byte_out_2;
  wire       [2:0]    mul3_78_port_byte_out_3;
  wire       [2:0]    mul3_78_port_byte_out_4;
  wire       [2:0]    mul3_78_port_byte_out_5;
  wire       [2:0]    mul3_78_port_byte_out_6;
  wire       [2:0]    mul3_78_port_byte_out_7;
  wire       [2:0]    mul2_79_port_byte_out_0;
  wire       [2:0]    mul2_79_port_byte_out_1;
  wire       [2:0]    mul2_79_port_byte_out_2;
  wire       [2:0]    mul2_79_port_byte_out_3;
  wire       [2:0]    mul2_79_port_byte_out_4;
  wire       [2:0]    mul2_79_port_byte_out_5;
  wire       [2:0]    mul2_79_port_byte_out_6;
  wire       [2:0]    mul2_79_port_byte_out_7;
  wire       [2:0]    mul3_79_port_byte_out_0;
  wire       [2:0]    mul3_79_port_byte_out_1;
  wire       [2:0]    mul3_79_port_byte_out_2;
  wire       [2:0]    mul3_79_port_byte_out_3;
  wire       [2:0]    mul3_79_port_byte_out_4;
  wire       [2:0]    mul3_79_port_byte_out_5;
  wire       [2:0]    mul3_79_port_byte_out_6;
  wire       [2:0]    mul3_79_port_byte_out_7;
  wire       [2:0]    mul2_80_port_byte_out_0;
  wire       [2:0]    mul2_80_port_byte_out_1;
  wire       [2:0]    mul2_80_port_byte_out_2;
  wire       [2:0]    mul2_80_port_byte_out_3;
  wire       [2:0]    mul2_80_port_byte_out_4;
  wire       [2:0]    mul2_80_port_byte_out_5;
  wire       [2:0]    mul2_80_port_byte_out_6;
  wire       [2:0]    mul2_80_port_byte_out_7;
  wire       [2:0]    mul3_80_port_byte_out_0;
  wire       [2:0]    mul3_80_port_byte_out_1;
  wire       [2:0]    mul3_80_port_byte_out_2;
  wire       [2:0]    mul3_80_port_byte_out_3;
  wire       [2:0]    mul3_80_port_byte_out_4;
  wire       [2:0]    mul3_80_port_byte_out_5;
  wire       [2:0]    mul3_80_port_byte_out_6;
  wire       [2:0]    mul3_80_port_byte_out_7;
  wire       [2:0]    mul2_81_port_byte_out_0;
  wire       [2:0]    mul2_81_port_byte_out_1;
  wire       [2:0]    mul2_81_port_byte_out_2;
  wire       [2:0]    mul2_81_port_byte_out_3;
  wire       [2:0]    mul2_81_port_byte_out_4;
  wire       [2:0]    mul2_81_port_byte_out_5;
  wire       [2:0]    mul2_81_port_byte_out_6;
  wire       [2:0]    mul2_81_port_byte_out_7;
  wire       [2:0]    mul3_81_port_byte_out_0;
  wire       [2:0]    mul3_81_port_byte_out_1;
  wire       [2:0]    mul3_81_port_byte_out_2;
  wire       [2:0]    mul3_81_port_byte_out_3;
  wire       [2:0]    mul3_81_port_byte_out_4;
  wire       [2:0]    mul3_81_port_byte_out_5;
  wire       [2:0]    mul3_81_port_byte_out_6;
  wire       [2:0]    mul3_81_port_byte_out_7;
  wire       [2:0]    mul2_82_port_byte_out_0;
  wire       [2:0]    mul2_82_port_byte_out_1;
  wire       [2:0]    mul2_82_port_byte_out_2;
  wire       [2:0]    mul2_82_port_byte_out_3;
  wire       [2:0]    mul2_82_port_byte_out_4;
  wire       [2:0]    mul2_82_port_byte_out_5;
  wire       [2:0]    mul2_82_port_byte_out_6;
  wire       [2:0]    mul2_82_port_byte_out_7;
  wire       [2:0]    mul3_82_port_byte_out_0;
  wire       [2:0]    mul3_82_port_byte_out_1;
  wire       [2:0]    mul3_82_port_byte_out_2;
  wire       [2:0]    mul3_82_port_byte_out_3;
  wire       [2:0]    mul3_82_port_byte_out_4;
  wire       [2:0]    mul3_82_port_byte_out_5;
  wire       [2:0]    mul3_82_port_byte_out_6;
  wire       [2:0]    mul3_82_port_byte_out_7;
  wire       [2:0]    mul2_83_port_byte_out_0;
  wire       [2:0]    mul2_83_port_byte_out_1;
  wire       [2:0]    mul2_83_port_byte_out_2;
  wire       [2:0]    mul2_83_port_byte_out_3;
  wire       [2:0]    mul2_83_port_byte_out_4;
  wire       [2:0]    mul2_83_port_byte_out_5;
  wire       [2:0]    mul2_83_port_byte_out_6;
  wire       [2:0]    mul2_83_port_byte_out_7;
  wire       [2:0]    mul3_83_port_byte_out_0;
  wire       [2:0]    mul3_83_port_byte_out_1;
  wire       [2:0]    mul3_83_port_byte_out_2;
  wire       [2:0]    mul3_83_port_byte_out_3;
  wire       [2:0]    mul3_83_port_byte_out_4;
  wire       [2:0]    mul3_83_port_byte_out_5;
  wire       [2:0]    mul3_83_port_byte_out_6;
  wire       [2:0]    mul3_83_port_byte_out_7;
  wire       [2:0]    mul2_84_port_byte_out_0;
  wire       [2:0]    mul2_84_port_byte_out_1;
  wire       [2:0]    mul2_84_port_byte_out_2;
  wire       [2:0]    mul2_84_port_byte_out_3;
  wire       [2:0]    mul2_84_port_byte_out_4;
  wire       [2:0]    mul2_84_port_byte_out_5;
  wire       [2:0]    mul2_84_port_byte_out_6;
  wire       [2:0]    mul2_84_port_byte_out_7;
  wire       [2:0]    mul3_84_port_byte_out_0;
  wire       [2:0]    mul3_84_port_byte_out_1;
  wire       [2:0]    mul3_84_port_byte_out_2;
  wire       [2:0]    mul3_84_port_byte_out_3;
  wire       [2:0]    mul3_84_port_byte_out_4;
  wire       [2:0]    mul3_84_port_byte_out_5;
  wire       [2:0]    mul3_84_port_byte_out_6;
  wire       [2:0]    mul3_84_port_byte_out_7;
  wire       [2:0]    mul2_85_port_byte_out_0;
  wire       [2:0]    mul2_85_port_byte_out_1;
  wire       [2:0]    mul2_85_port_byte_out_2;
  wire       [2:0]    mul2_85_port_byte_out_3;
  wire       [2:0]    mul2_85_port_byte_out_4;
  wire       [2:0]    mul2_85_port_byte_out_5;
  wire       [2:0]    mul2_85_port_byte_out_6;
  wire       [2:0]    mul2_85_port_byte_out_7;
  wire       [2:0]    mul3_85_port_byte_out_0;
  wire       [2:0]    mul3_85_port_byte_out_1;
  wire       [2:0]    mul3_85_port_byte_out_2;
  wire       [2:0]    mul3_85_port_byte_out_3;
  wire       [2:0]    mul3_85_port_byte_out_4;
  wire       [2:0]    mul3_85_port_byte_out_5;
  wire       [2:0]    mul3_85_port_byte_out_6;
  wire       [2:0]    mul3_85_port_byte_out_7;
  wire       [2:0]    mul2_86_port_byte_out_0;
  wire       [2:0]    mul2_86_port_byte_out_1;
  wire       [2:0]    mul2_86_port_byte_out_2;
  wire       [2:0]    mul2_86_port_byte_out_3;
  wire       [2:0]    mul2_86_port_byte_out_4;
  wire       [2:0]    mul2_86_port_byte_out_5;
  wire       [2:0]    mul2_86_port_byte_out_6;
  wire       [2:0]    mul2_86_port_byte_out_7;
  wire       [2:0]    mul3_86_port_byte_out_0;
  wire       [2:0]    mul3_86_port_byte_out_1;
  wire       [2:0]    mul3_86_port_byte_out_2;
  wire       [2:0]    mul3_86_port_byte_out_3;
  wire       [2:0]    mul3_86_port_byte_out_4;
  wire       [2:0]    mul3_86_port_byte_out_5;
  wire       [2:0]    mul3_86_port_byte_out_6;
  wire       [2:0]    mul3_86_port_byte_out_7;
  wire       [2:0]    mul2_87_port_byte_out_0;
  wire       [2:0]    mul2_87_port_byte_out_1;
  wire       [2:0]    mul2_87_port_byte_out_2;
  wire       [2:0]    mul2_87_port_byte_out_3;
  wire       [2:0]    mul2_87_port_byte_out_4;
  wire       [2:0]    mul2_87_port_byte_out_5;
  wire       [2:0]    mul2_87_port_byte_out_6;
  wire       [2:0]    mul2_87_port_byte_out_7;
  wire       [2:0]    mul3_87_port_byte_out_0;
  wire       [2:0]    mul3_87_port_byte_out_1;
  wire       [2:0]    mul3_87_port_byte_out_2;
  wire       [2:0]    mul3_87_port_byte_out_3;
  wire       [2:0]    mul3_87_port_byte_out_4;
  wire       [2:0]    mul3_87_port_byte_out_5;
  wire       [2:0]    mul3_87_port_byte_out_6;
  wire       [2:0]    mul3_87_port_byte_out_7;
  wire       [2:0]    mul2_88_port_byte_out_0;
  wire       [2:0]    mul2_88_port_byte_out_1;
  wire       [2:0]    mul2_88_port_byte_out_2;
  wire       [2:0]    mul2_88_port_byte_out_3;
  wire       [2:0]    mul2_88_port_byte_out_4;
  wire       [2:0]    mul2_88_port_byte_out_5;
  wire       [2:0]    mul2_88_port_byte_out_6;
  wire       [2:0]    mul2_88_port_byte_out_7;
  wire       [2:0]    mul3_88_port_byte_out_0;
  wire       [2:0]    mul3_88_port_byte_out_1;
  wire       [2:0]    mul3_88_port_byte_out_2;
  wire       [2:0]    mul3_88_port_byte_out_3;
  wire       [2:0]    mul3_88_port_byte_out_4;
  wire       [2:0]    mul3_88_port_byte_out_5;
  wire       [2:0]    mul3_88_port_byte_out_6;
  wire       [2:0]    mul3_88_port_byte_out_7;
  wire       [2:0]    mul2_89_port_byte_out_0;
  wire       [2:0]    mul2_89_port_byte_out_1;
  wire       [2:0]    mul2_89_port_byte_out_2;
  wire       [2:0]    mul2_89_port_byte_out_3;
  wire       [2:0]    mul2_89_port_byte_out_4;
  wire       [2:0]    mul2_89_port_byte_out_5;
  wire       [2:0]    mul2_89_port_byte_out_6;
  wire       [2:0]    mul2_89_port_byte_out_7;
  wire       [2:0]    mul3_89_port_byte_out_0;
  wire       [2:0]    mul3_89_port_byte_out_1;
  wire       [2:0]    mul3_89_port_byte_out_2;
  wire       [2:0]    mul3_89_port_byte_out_3;
  wire       [2:0]    mul3_89_port_byte_out_4;
  wire       [2:0]    mul3_89_port_byte_out_5;
  wire       [2:0]    mul3_89_port_byte_out_6;
  wire       [2:0]    mul3_89_port_byte_out_7;
  wire       [2:0]    mul2_90_port_byte_out_0;
  wire       [2:0]    mul2_90_port_byte_out_1;
  wire       [2:0]    mul2_90_port_byte_out_2;
  wire       [2:0]    mul2_90_port_byte_out_3;
  wire       [2:0]    mul2_90_port_byte_out_4;
  wire       [2:0]    mul2_90_port_byte_out_5;
  wire       [2:0]    mul2_90_port_byte_out_6;
  wire       [2:0]    mul2_90_port_byte_out_7;
  wire       [2:0]    mul3_90_port_byte_out_0;
  wire       [2:0]    mul3_90_port_byte_out_1;
  wire       [2:0]    mul3_90_port_byte_out_2;
  wire       [2:0]    mul3_90_port_byte_out_3;
  wire       [2:0]    mul3_90_port_byte_out_4;
  wire       [2:0]    mul3_90_port_byte_out_5;
  wire       [2:0]    mul3_90_port_byte_out_6;
  wire       [2:0]    mul3_90_port_byte_out_7;
  wire       [2:0]    mul2_91_port_byte_out_0;
  wire       [2:0]    mul2_91_port_byte_out_1;
  wire       [2:0]    mul2_91_port_byte_out_2;
  wire       [2:0]    mul2_91_port_byte_out_3;
  wire       [2:0]    mul2_91_port_byte_out_4;
  wire       [2:0]    mul2_91_port_byte_out_5;
  wire       [2:0]    mul2_91_port_byte_out_6;
  wire       [2:0]    mul2_91_port_byte_out_7;
  wire       [2:0]    mul3_91_port_byte_out_0;
  wire       [2:0]    mul3_91_port_byte_out_1;
  wire       [2:0]    mul3_91_port_byte_out_2;
  wire       [2:0]    mul3_91_port_byte_out_3;
  wire       [2:0]    mul3_91_port_byte_out_4;
  wire       [2:0]    mul3_91_port_byte_out_5;
  wire       [2:0]    mul3_91_port_byte_out_6;
  wire       [2:0]    mul3_91_port_byte_out_7;
  wire       [2:0]    mul2_92_port_byte_out_0;
  wire       [2:0]    mul2_92_port_byte_out_1;
  wire       [2:0]    mul2_92_port_byte_out_2;
  wire       [2:0]    mul2_92_port_byte_out_3;
  wire       [2:0]    mul2_92_port_byte_out_4;
  wire       [2:0]    mul2_92_port_byte_out_5;
  wire       [2:0]    mul2_92_port_byte_out_6;
  wire       [2:0]    mul2_92_port_byte_out_7;
  wire       [2:0]    mul3_92_port_byte_out_0;
  wire       [2:0]    mul3_92_port_byte_out_1;
  wire       [2:0]    mul3_92_port_byte_out_2;
  wire       [2:0]    mul3_92_port_byte_out_3;
  wire       [2:0]    mul3_92_port_byte_out_4;
  wire       [2:0]    mul3_92_port_byte_out_5;
  wire       [2:0]    mul3_92_port_byte_out_6;
  wire       [2:0]    mul3_92_port_byte_out_7;
  wire       [2:0]    mul2_93_port_byte_out_0;
  wire       [2:0]    mul2_93_port_byte_out_1;
  wire       [2:0]    mul2_93_port_byte_out_2;
  wire       [2:0]    mul2_93_port_byte_out_3;
  wire       [2:0]    mul2_93_port_byte_out_4;
  wire       [2:0]    mul2_93_port_byte_out_5;
  wire       [2:0]    mul2_93_port_byte_out_6;
  wire       [2:0]    mul2_93_port_byte_out_7;
  wire       [2:0]    mul3_93_port_byte_out_0;
  wire       [2:0]    mul3_93_port_byte_out_1;
  wire       [2:0]    mul3_93_port_byte_out_2;
  wire       [2:0]    mul3_93_port_byte_out_3;
  wire       [2:0]    mul3_93_port_byte_out_4;
  wire       [2:0]    mul3_93_port_byte_out_5;
  wire       [2:0]    mul3_93_port_byte_out_6;
  wire       [2:0]    mul3_93_port_byte_out_7;
  wire       [2:0]    mul2_94_port_byte_out_0;
  wire       [2:0]    mul2_94_port_byte_out_1;
  wire       [2:0]    mul2_94_port_byte_out_2;
  wire       [2:0]    mul2_94_port_byte_out_3;
  wire       [2:0]    mul2_94_port_byte_out_4;
  wire       [2:0]    mul2_94_port_byte_out_5;
  wire       [2:0]    mul2_94_port_byte_out_6;
  wire       [2:0]    mul2_94_port_byte_out_7;
  wire       [2:0]    mul3_94_port_byte_out_0;
  wire       [2:0]    mul3_94_port_byte_out_1;
  wire       [2:0]    mul3_94_port_byte_out_2;
  wire       [2:0]    mul3_94_port_byte_out_3;
  wire       [2:0]    mul3_94_port_byte_out_4;
  wire       [2:0]    mul3_94_port_byte_out_5;
  wire       [2:0]    mul3_94_port_byte_out_6;
  wire       [2:0]    mul3_94_port_byte_out_7;
  wire       [2:0]    mul2_95_port_byte_out_0;
  wire       [2:0]    mul2_95_port_byte_out_1;
  wire       [2:0]    mul2_95_port_byte_out_2;
  wire       [2:0]    mul2_95_port_byte_out_3;
  wire       [2:0]    mul2_95_port_byte_out_4;
  wire       [2:0]    mul2_95_port_byte_out_5;
  wire       [2:0]    mul2_95_port_byte_out_6;
  wire       [2:0]    mul2_95_port_byte_out_7;
  wire       [2:0]    mul3_95_port_byte_out_0;
  wire       [2:0]    mul3_95_port_byte_out_1;
  wire       [2:0]    mul3_95_port_byte_out_2;
  wire       [2:0]    mul3_95_port_byte_out_3;
  wire       [2:0]    mul3_95_port_byte_out_4;
  wire       [2:0]    mul3_95_port_byte_out_5;
  wire       [2:0]    mul3_95_port_byte_out_6;
  wire       [2:0]    mul3_95_port_byte_out_7;
  wire       [2:0]    mul2_96_port_byte_out_0;
  wire       [2:0]    mul2_96_port_byte_out_1;
  wire       [2:0]    mul2_96_port_byte_out_2;
  wire       [2:0]    mul2_96_port_byte_out_3;
  wire       [2:0]    mul2_96_port_byte_out_4;
  wire       [2:0]    mul2_96_port_byte_out_5;
  wire       [2:0]    mul2_96_port_byte_out_6;
  wire       [2:0]    mul2_96_port_byte_out_7;
  wire       [2:0]    mul3_96_port_byte_out_0;
  wire       [2:0]    mul3_96_port_byte_out_1;
  wire       [2:0]    mul3_96_port_byte_out_2;
  wire       [2:0]    mul3_96_port_byte_out_3;
  wire       [2:0]    mul3_96_port_byte_out_4;
  wire       [2:0]    mul3_96_port_byte_out_5;
  wire       [2:0]    mul3_96_port_byte_out_6;
  wire       [2:0]    mul3_96_port_byte_out_7;
  wire       [2:0]    mul2_97_port_byte_out_0;
  wire       [2:0]    mul2_97_port_byte_out_1;
  wire       [2:0]    mul2_97_port_byte_out_2;
  wire       [2:0]    mul2_97_port_byte_out_3;
  wire       [2:0]    mul2_97_port_byte_out_4;
  wire       [2:0]    mul2_97_port_byte_out_5;
  wire       [2:0]    mul2_97_port_byte_out_6;
  wire       [2:0]    mul2_97_port_byte_out_7;
  wire       [2:0]    mul3_97_port_byte_out_0;
  wire       [2:0]    mul3_97_port_byte_out_1;
  wire       [2:0]    mul3_97_port_byte_out_2;
  wire       [2:0]    mul3_97_port_byte_out_3;
  wire       [2:0]    mul3_97_port_byte_out_4;
  wire       [2:0]    mul3_97_port_byte_out_5;
  wire       [2:0]    mul3_97_port_byte_out_6;
  wire       [2:0]    mul3_97_port_byte_out_7;
  wire       [2:0]    mul2_98_port_byte_out_0;
  wire       [2:0]    mul2_98_port_byte_out_1;
  wire       [2:0]    mul2_98_port_byte_out_2;
  wire       [2:0]    mul2_98_port_byte_out_3;
  wire       [2:0]    mul2_98_port_byte_out_4;
  wire       [2:0]    mul2_98_port_byte_out_5;
  wire       [2:0]    mul2_98_port_byte_out_6;
  wire       [2:0]    mul2_98_port_byte_out_7;
  wire       [2:0]    mul3_98_port_byte_out_0;
  wire       [2:0]    mul3_98_port_byte_out_1;
  wire       [2:0]    mul3_98_port_byte_out_2;
  wire       [2:0]    mul3_98_port_byte_out_3;
  wire       [2:0]    mul3_98_port_byte_out_4;
  wire       [2:0]    mul3_98_port_byte_out_5;
  wire       [2:0]    mul3_98_port_byte_out_6;
  wire       [2:0]    mul3_98_port_byte_out_7;
  wire       [2:0]    mul2_99_port_byte_out_0;
  wire       [2:0]    mul2_99_port_byte_out_1;
  wire       [2:0]    mul2_99_port_byte_out_2;
  wire       [2:0]    mul2_99_port_byte_out_3;
  wire       [2:0]    mul2_99_port_byte_out_4;
  wire       [2:0]    mul2_99_port_byte_out_5;
  wire       [2:0]    mul2_99_port_byte_out_6;
  wire       [2:0]    mul2_99_port_byte_out_7;
  wire       [2:0]    mul3_99_port_byte_out_0;
  wire       [2:0]    mul3_99_port_byte_out_1;
  wire       [2:0]    mul3_99_port_byte_out_2;
  wire       [2:0]    mul3_99_port_byte_out_3;
  wire       [2:0]    mul3_99_port_byte_out_4;
  wire       [2:0]    mul3_99_port_byte_out_5;
  wire       [2:0]    mul3_99_port_byte_out_6;
  wire       [2:0]    mul3_99_port_byte_out_7;
  wire       [2:0]    mul2_100_port_byte_out_0;
  wire       [2:0]    mul2_100_port_byte_out_1;
  wire       [2:0]    mul2_100_port_byte_out_2;
  wire       [2:0]    mul2_100_port_byte_out_3;
  wire       [2:0]    mul2_100_port_byte_out_4;
  wire       [2:0]    mul2_100_port_byte_out_5;
  wire       [2:0]    mul2_100_port_byte_out_6;
  wire       [2:0]    mul2_100_port_byte_out_7;
  wire       [2:0]    mul3_100_port_byte_out_0;
  wire       [2:0]    mul3_100_port_byte_out_1;
  wire       [2:0]    mul3_100_port_byte_out_2;
  wire       [2:0]    mul3_100_port_byte_out_3;
  wire       [2:0]    mul3_100_port_byte_out_4;
  wire       [2:0]    mul3_100_port_byte_out_5;
  wire       [2:0]    mul3_100_port_byte_out_6;
  wire       [2:0]    mul3_100_port_byte_out_7;
  wire       [2:0]    mul2_101_port_byte_out_0;
  wire       [2:0]    mul2_101_port_byte_out_1;
  wire       [2:0]    mul2_101_port_byte_out_2;
  wire       [2:0]    mul2_101_port_byte_out_3;
  wire       [2:0]    mul2_101_port_byte_out_4;
  wire       [2:0]    mul2_101_port_byte_out_5;
  wire       [2:0]    mul2_101_port_byte_out_6;
  wire       [2:0]    mul2_101_port_byte_out_7;
  wire       [2:0]    mul3_101_port_byte_out_0;
  wire       [2:0]    mul3_101_port_byte_out_1;
  wire       [2:0]    mul3_101_port_byte_out_2;
  wire       [2:0]    mul3_101_port_byte_out_3;
  wire       [2:0]    mul3_101_port_byte_out_4;
  wire       [2:0]    mul3_101_port_byte_out_5;
  wire       [2:0]    mul3_101_port_byte_out_6;
  wire       [2:0]    mul3_101_port_byte_out_7;
  wire       [2:0]    mul2_102_port_byte_out_0;
  wire       [2:0]    mul2_102_port_byte_out_1;
  wire       [2:0]    mul2_102_port_byte_out_2;
  wire       [2:0]    mul2_102_port_byte_out_3;
  wire       [2:0]    mul2_102_port_byte_out_4;
  wire       [2:0]    mul2_102_port_byte_out_5;
  wire       [2:0]    mul2_102_port_byte_out_6;
  wire       [2:0]    mul2_102_port_byte_out_7;
  wire       [2:0]    mul3_102_port_byte_out_0;
  wire       [2:0]    mul3_102_port_byte_out_1;
  wire       [2:0]    mul3_102_port_byte_out_2;
  wire       [2:0]    mul3_102_port_byte_out_3;
  wire       [2:0]    mul3_102_port_byte_out_4;
  wire       [2:0]    mul3_102_port_byte_out_5;
  wire       [2:0]    mul3_102_port_byte_out_6;
  wire       [2:0]    mul3_102_port_byte_out_7;
  wire       [2:0]    mul2_103_port_byte_out_0;
  wire       [2:0]    mul2_103_port_byte_out_1;
  wire       [2:0]    mul2_103_port_byte_out_2;
  wire       [2:0]    mul2_103_port_byte_out_3;
  wire       [2:0]    mul2_103_port_byte_out_4;
  wire       [2:0]    mul2_103_port_byte_out_5;
  wire       [2:0]    mul2_103_port_byte_out_6;
  wire       [2:0]    mul2_103_port_byte_out_7;
  wire       [2:0]    mul3_103_port_byte_out_0;
  wire       [2:0]    mul3_103_port_byte_out_1;
  wire       [2:0]    mul3_103_port_byte_out_2;
  wire       [2:0]    mul3_103_port_byte_out_3;
  wire       [2:0]    mul3_103_port_byte_out_4;
  wire       [2:0]    mul3_103_port_byte_out_5;
  wire       [2:0]    mul3_103_port_byte_out_6;
  wire       [2:0]    mul3_103_port_byte_out_7;
  wire       [2:0]    mul2_104_port_byte_out_0;
  wire       [2:0]    mul2_104_port_byte_out_1;
  wire       [2:0]    mul2_104_port_byte_out_2;
  wire       [2:0]    mul2_104_port_byte_out_3;
  wire       [2:0]    mul2_104_port_byte_out_4;
  wire       [2:0]    mul2_104_port_byte_out_5;
  wire       [2:0]    mul2_104_port_byte_out_6;
  wire       [2:0]    mul2_104_port_byte_out_7;
  wire       [2:0]    mul3_104_port_byte_out_0;
  wire       [2:0]    mul3_104_port_byte_out_1;
  wire       [2:0]    mul3_104_port_byte_out_2;
  wire       [2:0]    mul3_104_port_byte_out_3;
  wire       [2:0]    mul3_104_port_byte_out_4;
  wire       [2:0]    mul3_104_port_byte_out_5;
  wire       [2:0]    mul3_104_port_byte_out_6;
  wire       [2:0]    mul3_104_port_byte_out_7;
  wire       [2:0]    mul2_105_port_byte_out_0;
  wire       [2:0]    mul2_105_port_byte_out_1;
  wire       [2:0]    mul2_105_port_byte_out_2;
  wire       [2:0]    mul2_105_port_byte_out_3;
  wire       [2:0]    mul2_105_port_byte_out_4;
  wire       [2:0]    mul2_105_port_byte_out_5;
  wire       [2:0]    mul2_105_port_byte_out_6;
  wire       [2:0]    mul2_105_port_byte_out_7;
  wire       [2:0]    mul3_105_port_byte_out_0;
  wire       [2:0]    mul3_105_port_byte_out_1;
  wire       [2:0]    mul3_105_port_byte_out_2;
  wire       [2:0]    mul3_105_port_byte_out_3;
  wire       [2:0]    mul3_105_port_byte_out_4;
  wire       [2:0]    mul3_105_port_byte_out_5;
  wire       [2:0]    mul3_105_port_byte_out_6;
  wire       [2:0]    mul3_105_port_byte_out_7;
  wire       [2:0]    mul2_106_port_byte_out_0;
  wire       [2:0]    mul2_106_port_byte_out_1;
  wire       [2:0]    mul2_106_port_byte_out_2;
  wire       [2:0]    mul2_106_port_byte_out_3;
  wire       [2:0]    mul2_106_port_byte_out_4;
  wire       [2:0]    mul2_106_port_byte_out_5;
  wire       [2:0]    mul2_106_port_byte_out_6;
  wire       [2:0]    mul2_106_port_byte_out_7;
  wire       [2:0]    mul3_106_port_byte_out_0;
  wire       [2:0]    mul3_106_port_byte_out_1;
  wire       [2:0]    mul3_106_port_byte_out_2;
  wire       [2:0]    mul3_106_port_byte_out_3;
  wire       [2:0]    mul3_106_port_byte_out_4;
  wire       [2:0]    mul3_106_port_byte_out_5;
  wire       [2:0]    mul3_106_port_byte_out_6;
  wire       [2:0]    mul3_106_port_byte_out_7;
  wire       [2:0]    mul2_107_port_byte_out_0;
  wire       [2:0]    mul2_107_port_byte_out_1;
  wire       [2:0]    mul2_107_port_byte_out_2;
  wire       [2:0]    mul2_107_port_byte_out_3;
  wire       [2:0]    mul2_107_port_byte_out_4;
  wire       [2:0]    mul2_107_port_byte_out_5;
  wire       [2:0]    mul2_107_port_byte_out_6;
  wire       [2:0]    mul2_107_port_byte_out_7;
  wire       [2:0]    mul3_107_port_byte_out_0;
  wire       [2:0]    mul3_107_port_byte_out_1;
  wire       [2:0]    mul3_107_port_byte_out_2;
  wire       [2:0]    mul3_107_port_byte_out_3;
  wire       [2:0]    mul3_107_port_byte_out_4;
  wire       [2:0]    mul3_107_port_byte_out_5;
  wire       [2:0]    mul3_107_port_byte_out_6;
  wire       [2:0]    mul3_107_port_byte_out_7;
  wire       [2:0]    mul2_108_port_byte_out_0;
  wire       [2:0]    mul2_108_port_byte_out_1;
  wire       [2:0]    mul2_108_port_byte_out_2;
  wire       [2:0]    mul2_108_port_byte_out_3;
  wire       [2:0]    mul2_108_port_byte_out_4;
  wire       [2:0]    mul2_108_port_byte_out_5;
  wire       [2:0]    mul2_108_port_byte_out_6;
  wire       [2:0]    mul2_108_port_byte_out_7;
  wire       [2:0]    mul3_108_port_byte_out_0;
  wire       [2:0]    mul3_108_port_byte_out_1;
  wire       [2:0]    mul3_108_port_byte_out_2;
  wire       [2:0]    mul3_108_port_byte_out_3;
  wire       [2:0]    mul3_108_port_byte_out_4;
  wire       [2:0]    mul3_108_port_byte_out_5;
  wire       [2:0]    mul3_108_port_byte_out_6;
  wire       [2:0]    mul3_108_port_byte_out_7;
  wire       [2:0]    mul2_109_port_byte_out_0;
  wire       [2:0]    mul2_109_port_byte_out_1;
  wire       [2:0]    mul2_109_port_byte_out_2;
  wire       [2:0]    mul2_109_port_byte_out_3;
  wire       [2:0]    mul2_109_port_byte_out_4;
  wire       [2:0]    mul2_109_port_byte_out_5;
  wire       [2:0]    mul2_109_port_byte_out_6;
  wire       [2:0]    mul2_109_port_byte_out_7;
  wire       [2:0]    mul3_109_port_byte_out_0;
  wire       [2:0]    mul3_109_port_byte_out_1;
  wire       [2:0]    mul3_109_port_byte_out_2;
  wire       [2:0]    mul3_109_port_byte_out_3;
  wire       [2:0]    mul3_109_port_byte_out_4;
  wire       [2:0]    mul3_109_port_byte_out_5;
  wire       [2:0]    mul3_109_port_byte_out_6;
  wire       [2:0]    mul3_109_port_byte_out_7;
  wire       [2:0]    mul2_110_port_byte_out_0;
  wire       [2:0]    mul2_110_port_byte_out_1;
  wire       [2:0]    mul2_110_port_byte_out_2;
  wire       [2:0]    mul2_110_port_byte_out_3;
  wire       [2:0]    mul2_110_port_byte_out_4;
  wire       [2:0]    mul2_110_port_byte_out_5;
  wire       [2:0]    mul2_110_port_byte_out_6;
  wire       [2:0]    mul2_110_port_byte_out_7;
  wire       [2:0]    mul3_110_port_byte_out_0;
  wire       [2:0]    mul3_110_port_byte_out_1;
  wire       [2:0]    mul3_110_port_byte_out_2;
  wire       [2:0]    mul3_110_port_byte_out_3;
  wire       [2:0]    mul3_110_port_byte_out_4;
  wire       [2:0]    mul3_110_port_byte_out_5;
  wire       [2:0]    mul3_110_port_byte_out_6;
  wire       [2:0]    mul3_110_port_byte_out_7;
  wire       [2:0]    mul2_111_port_byte_out_0;
  wire       [2:0]    mul2_111_port_byte_out_1;
  wire       [2:0]    mul2_111_port_byte_out_2;
  wire       [2:0]    mul2_111_port_byte_out_3;
  wire       [2:0]    mul2_111_port_byte_out_4;
  wire       [2:0]    mul2_111_port_byte_out_5;
  wire       [2:0]    mul2_111_port_byte_out_6;
  wire       [2:0]    mul2_111_port_byte_out_7;
  wire       [2:0]    mul3_111_port_byte_out_0;
  wire       [2:0]    mul3_111_port_byte_out_1;
  wire       [2:0]    mul3_111_port_byte_out_2;
  wire       [2:0]    mul3_111_port_byte_out_3;
  wire       [2:0]    mul3_111_port_byte_out_4;
  wire       [2:0]    mul3_111_port_byte_out_5;
  wire       [2:0]    mul3_111_port_byte_out_6;
  wire       [2:0]    mul3_111_port_byte_out_7;
  wire       [2:0]    mul2_112_port_byte_out_0;
  wire       [2:0]    mul2_112_port_byte_out_1;
  wire       [2:0]    mul2_112_port_byte_out_2;
  wire       [2:0]    mul2_112_port_byte_out_3;
  wire       [2:0]    mul2_112_port_byte_out_4;
  wire       [2:0]    mul2_112_port_byte_out_5;
  wire       [2:0]    mul2_112_port_byte_out_6;
  wire       [2:0]    mul2_112_port_byte_out_7;
  wire       [2:0]    mul3_112_port_byte_out_0;
  wire       [2:0]    mul3_112_port_byte_out_1;
  wire       [2:0]    mul3_112_port_byte_out_2;
  wire       [2:0]    mul3_112_port_byte_out_3;
  wire       [2:0]    mul3_112_port_byte_out_4;
  wire       [2:0]    mul3_112_port_byte_out_5;
  wire       [2:0]    mul3_112_port_byte_out_6;
  wire       [2:0]    mul3_112_port_byte_out_7;
  wire       [2:0]    mul2_113_port_byte_out_0;
  wire       [2:0]    mul2_113_port_byte_out_1;
  wire       [2:0]    mul2_113_port_byte_out_2;
  wire       [2:0]    mul2_113_port_byte_out_3;
  wire       [2:0]    mul2_113_port_byte_out_4;
  wire       [2:0]    mul2_113_port_byte_out_5;
  wire       [2:0]    mul2_113_port_byte_out_6;
  wire       [2:0]    mul2_113_port_byte_out_7;
  wire       [2:0]    mul3_113_port_byte_out_0;
  wire       [2:0]    mul3_113_port_byte_out_1;
  wire       [2:0]    mul3_113_port_byte_out_2;
  wire       [2:0]    mul3_113_port_byte_out_3;
  wire       [2:0]    mul3_113_port_byte_out_4;
  wire       [2:0]    mul3_113_port_byte_out_5;
  wire       [2:0]    mul3_113_port_byte_out_6;
  wire       [2:0]    mul3_113_port_byte_out_7;
  wire       [2:0]    mul2_114_port_byte_out_0;
  wire       [2:0]    mul2_114_port_byte_out_1;
  wire       [2:0]    mul2_114_port_byte_out_2;
  wire       [2:0]    mul2_114_port_byte_out_3;
  wire       [2:0]    mul2_114_port_byte_out_4;
  wire       [2:0]    mul2_114_port_byte_out_5;
  wire       [2:0]    mul2_114_port_byte_out_6;
  wire       [2:0]    mul2_114_port_byte_out_7;
  wire       [2:0]    mul3_114_port_byte_out_0;
  wire       [2:0]    mul3_114_port_byte_out_1;
  wire       [2:0]    mul3_114_port_byte_out_2;
  wire       [2:0]    mul3_114_port_byte_out_3;
  wire       [2:0]    mul3_114_port_byte_out_4;
  wire       [2:0]    mul3_114_port_byte_out_5;
  wire       [2:0]    mul3_114_port_byte_out_6;
  wire       [2:0]    mul3_114_port_byte_out_7;
  wire       [2:0]    mul2_115_port_byte_out_0;
  wire       [2:0]    mul2_115_port_byte_out_1;
  wire       [2:0]    mul2_115_port_byte_out_2;
  wire       [2:0]    mul2_115_port_byte_out_3;
  wire       [2:0]    mul2_115_port_byte_out_4;
  wire       [2:0]    mul2_115_port_byte_out_5;
  wire       [2:0]    mul2_115_port_byte_out_6;
  wire       [2:0]    mul2_115_port_byte_out_7;
  wire       [2:0]    mul3_115_port_byte_out_0;
  wire       [2:0]    mul3_115_port_byte_out_1;
  wire       [2:0]    mul3_115_port_byte_out_2;
  wire       [2:0]    mul3_115_port_byte_out_3;
  wire       [2:0]    mul3_115_port_byte_out_4;
  wire       [2:0]    mul3_115_port_byte_out_5;
  wire       [2:0]    mul3_115_port_byte_out_6;
  wire       [2:0]    mul3_115_port_byte_out_7;
  wire       [2:0]    mul2_116_port_byte_out_0;
  wire       [2:0]    mul2_116_port_byte_out_1;
  wire       [2:0]    mul2_116_port_byte_out_2;
  wire       [2:0]    mul2_116_port_byte_out_3;
  wire       [2:0]    mul2_116_port_byte_out_4;
  wire       [2:0]    mul2_116_port_byte_out_5;
  wire       [2:0]    mul2_116_port_byte_out_6;
  wire       [2:0]    mul2_116_port_byte_out_7;
  wire       [2:0]    mul3_116_port_byte_out_0;
  wire       [2:0]    mul3_116_port_byte_out_1;
  wire       [2:0]    mul3_116_port_byte_out_2;
  wire       [2:0]    mul3_116_port_byte_out_3;
  wire       [2:0]    mul3_116_port_byte_out_4;
  wire       [2:0]    mul3_116_port_byte_out_5;
  wire       [2:0]    mul3_116_port_byte_out_6;
  wire       [2:0]    mul3_116_port_byte_out_7;
  wire       [2:0]    mul2_117_port_byte_out_0;
  wire       [2:0]    mul2_117_port_byte_out_1;
  wire       [2:0]    mul2_117_port_byte_out_2;
  wire       [2:0]    mul2_117_port_byte_out_3;
  wire       [2:0]    mul2_117_port_byte_out_4;
  wire       [2:0]    mul2_117_port_byte_out_5;
  wire       [2:0]    mul2_117_port_byte_out_6;
  wire       [2:0]    mul2_117_port_byte_out_7;
  wire       [2:0]    mul3_117_port_byte_out_0;
  wire       [2:0]    mul3_117_port_byte_out_1;
  wire       [2:0]    mul3_117_port_byte_out_2;
  wire       [2:0]    mul3_117_port_byte_out_3;
  wire       [2:0]    mul3_117_port_byte_out_4;
  wire       [2:0]    mul3_117_port_byte_out_5;
  wire       [2:0]    mul3_117_port_byte_out_6;
  wire       [2:0]    mul3_117_port_byte_out_7;
  wire       [2:0]    mul2_118_port_byte_out_0;
  wire       [2:0]    mul2_118_port_byte_out_1;
  wire       [2:0]    mul2_118_port_byte_out_2;
  wire       [2:0]    mul2_118_port_byte_out_3;
  wire       [2:0]    mul2_118_port_byte_out_4;
  wire       [2:0]    mul2_118_port_byte_out_5;
  wire       [2:0]    mul2_118_port_byte_out_6;
  wire       [2:0]    mul2_118_port_byte_out_7;
  wire       [2:0]    mul3_118_port_byte_out_0;
  wire       [2:0]    mul3_118_port_byte_out_1;
  wire       [2:0]    mul3_118_port_byte_out_2;
  wire       [2:0]    mul3_118_port_byte_out_3;
  wire       [2:0]    mul3_118_port_byte_out_4;
  wire       [2:0]    mul3_118_port_byte_out_5;
  wire       [2:0]    mul3_118_port_byte_out_6;
  wire       [2:0]    mul3_118_port_byte_out_7;
  wire       [2:0]    mul2_119_port_byte_out_0;
  wire       [2:0]    mul2_119_port_byte_out_1;
  wire       [2:0]    mul2_119_port_byte_out_2;
  wire       [2:0]    mul2_119_port_byte_out_3;
  wire       [2:0]    mul2_119_port_byte_out_4;
  wire       [2:0]    mul2_119_port_byte_out_5;
  wire       [2:0]    mul2_119_port_byte_out_6;
  wire       [2:0]    mul2_119_port_byte_out_7;
  wire       [2:0]    mul3_119_port_byte_out_0;
  wire       [2:0]    mul3_119_port_byte_out_1;
  wire       [2:0]    mul3_119_port_byte_out_2;
  wire       [2:0]    mul3_119_port_byte_out_3;
  wire       [2:0]    mul3_119_port_byte_out_4;
  wire       [2:0]    mul3_119_port_byte_out_5;
  wire       [2:0]    mul3_119_port_byte_out_6;
  wire       [2:0]    mul3_119_port_byte_out_7;
  wire       [2:0]    mul2_120_port_byte_out_0;
  wire       [2:0]    mul2_120_port_byte_out_1;
  wire       [2:0]    mul2_120_port_byte_out_2;
  wire       [2:0]    mul2_120_port_byte_out_3;
  wire       [2:0]    mul2_120_port_byte_out_4;
  wire       [2:0]    mul2_120_port_byte_out_5;
  wire       [2:0]    mul2_120_port_byte_out_6;
  wire       [2:0]    mul2_120_port_byte_out_7;
  wire       [2:0]    mul3_120_port_byte_out_0;
  wire       [2:0]    mul3_120_port_byte_out_1;
  wire       [2:0]    mul3_120_port_byte_out_2;
  wire       [2:0]    mul3_120_port_byte_out_3;
  wire       [2:0]    mul3_120_port_byte_out_4;
  wire       [2:0]    mul3_120_port_byte_out_5;
  wire       [2:0]    mul3_120_port_byte_out_6;
  wire       [2:0]    mul3_120_port_byte_out_7;
  wire       [2:0]    mul2_121_port_byte_out_0;
  wire       [2:0]    mul2_121_port_byte_out_1;
  wire       [2:0]    mul2_121_port_byte_out_2;
  wire       [2:0]    mul2_121_port_byte_out_3;
  wire       [2:0]    mul2_121_port_byte_out_4;
  wire       [2:0]    mul2_121_port_byte_out_5;
  wire       [2:0]    mul2_121_port_byte_out_6;
  wire       [2:0]    mul2_121_port_byte_out_7;
  wire       [2:0]    mul3_121_port_byte_out_0;
  wire       [2:0]    mul3_121_port_byte_out_1;
  wire       [2:0]    mul3_121_port_byte_out_2;
  wire       [2:0]    mul3_121_port_byte_out_3;
  wire       [2:0]    mul3_121_port_byte_out_4;
  wire       [2:0]    mul3_121_port_byte_out_5;
  wire       [2:0]    mul3_121_port_byte_out_6;
  wire       [2:0]    mul3_121_port_byte_out_7;
  wire       [2:0]    mul2_122_port_byte_out_0;
  wire       [2:0]    mul2_122_port_byte_out_1;
  wire       [2:0]    mul2_122_port_byte_out_2;
  wire       [2:0]    mul2_122_port_byte_out_3;
  wire       [2:0]    mul2_122_port_byte_out_4;
  wire       [2:0]    mul2_122_port_byte_out_5;
  wire       [2:0]    mul2_122_port_byte_out_6;
  wire       [2:0]    mul2_122_port_byte_out_7;
  wire       [2:0]    mul3_122_port_byte_out_0;
  wire       [2:0]    mul3_122_port_byte_out_1;
  wire       [2:0]    mul3_122_port_byte_out_2;
  wire       [2:0]    mul3_122_port_byte_out_3;
  wire       [2:0]    mul3_122_port_byte_out_4;
  wire       [2:0]    mul3_122_port_byte_out_5;
  wire       [2:0]    mul3_122_port_byte_out_6;
  wire       [2:0]    mul3_122_port_byte_out_7;
  wire       [2:0]    mul2_123_port_byte_out_0;
  wire       [2:0]    mul2_123_port_byte_out_1;
  wire       [2:0]    mul2_123_port_byte_out_2;
  wire       [2:0]    mul2_123_port_byte_out_3;
  wire       [2:0]    mul2_123_port_byte_out_4;
  wire       [2:0]    mul2_123_port_byte_out_5;
  wire       [2:0]    mul2_123_port_byte_out_6;
  wire       [2:0]    mul2_123_port_byte_out_7;
  wire       [2:0]    mul3_123_port_byte_out_0;
  wire       [2:0]    mul3_123_port_byte_out_1;
  wire       [2:0]    mul3_123_port_byte_out_2;
  wire       [2:0]    mul3_123_port_byte_out_3;
  wire       [2:0]    mul3_123_port_byte_out_4;
  wire       [2:0]    mul3_123_port_byte_out_5;
  wire       [2:0]    mul3_123_port_byte_out_6;
  wire       [2:0]    mul3_123_port_byte_out_7;
  wire       [2:0]    mul2_124_port_byte_out_0;
  wire       [2:0]    mul2_124_port_byte_out_1;
  wire       [2:0]    mul2_124_port_byte_out_2;
  wire       [2:0]    mul2_124_port_byte_out_3;
  wire       [2:0]    mul2_124_port_byte_out_4;
  wire       [2:0]    mul2_124_port_byte_out_5;
  wire       [2:0]    mul2_124_port_byte_out_6;
  wire       [2:0]    mul2_124_port_byte_out_7;
  wire       [2:0]    mul3_124_port_byte_out_0;
  wire       [2:0]    mul3_124_port_byte_out_1;
  wire       [2:0]    mul3_124_port_byte_out_2;
  wire       [2:0]    mul3_124_port_byte_out_3;
  wire       [2:0]    mul3_124_port_byte_out_4;
  wire       [2:0]    mul3_124_port_byte_out_5;
  wire       [2:0]    mul3_124_port_byte_out_6;
  wire       [2:0]    mul3_124_port_byte_out_7;
  wire       [2:0]    mul2_125_port_byte_out_0;
  wire       [2:0]    mul2_125_port_byte_out_1;
  wire       [2:0]    mul2_125_port_byte_out_2;
  wire       [2:0]    mul2_125_port_byte_out_3;
  wire       [2:0]    mul2_125_port_byte_out_4;
  wire       [2:0]    mul2_125_port_byte_out_5;
  wire       [2:0]    mul2_125_port_byte_out_6;
  wire       [2:0]    mul2_125_port_byte_out_7;
  wire       [2:0]    mul3_125_port_byte_out_0;
  wire       [2:0]    mul3_125_port_byte_out_1;
  wire       [2:0]    mul3_125_port_byte_out_2;
  wire       [2:0]    mul3_125_port_byte_out_3;
  wire       [2:0]    mul3_125_port_byte_out_4;
  wire       [2:0]    mul3_125_port_byte_out_5;
  wire       [2:0]    mul3_125_port_byte_out_6;
  wire       [2:0]    mul3_125_port_byte_out_7;
  wire       [2:0]    mul2_126_port_byte_out_0;
  wire       [2:0]    mul2_126_port_byte_out_1;
  wire       [2:0]    mul2_126_port_byte_out_2;
  wire       [2:0]    mul2_126_port_byte_out_3;
  wire       [2:0]    mul2_126_port_byte_out_4;
  wire       [2:0]    mul2_126_port_byte_out_5;
  wire       [2:0]    mul2_126_port_byte_out_6;
  wire       [2:0]    mul2_126_port_byte_out_7;
  wire       [2:0]    mul3_126_port_byte_out_0;
  wire       [2:0]    mul3_126_port_byte_out_1;
  wire       [2:0]    mul3_126_port_byte_out_2;
  wire       [2:0]    mul3_126_port_byte_out_3;
  wire       [2:0]    mul3_126_port_byte_out_4;
  wire       [2:0]    mul3_126_port_byte_out_5;
  wire       [2:0]    mul3_126_port_byte_out_6;
  wire       [2:0]    mul3_126_port_byte_out_7;
  wire       [2:0]    mul2_127_port_byte_out_0;
  wire       [2:0]    mul2_127_port_byte_out_1;
  wire       [2:0]    mul2_127_port_byte_out_2;
  wire       [2:0]    mul2_127_port_byte_out_3;
  wire       [2:0]    mul2_127_port_byte_out_4;
  wire       [2:0]    mul2_127_port_byte_out_5;
  wire       [2:0]    mul2_127_port_byte_out_6;
  wire       [2:0]    mul2_127_port_byte_out_7;
  wire       [2:0]    mul3_127_port_byte_out_0;
  wire       [2:0]    mul3_127_port_byte_out_1;
  wire       [2:0]    mul3_127_port_byte_out_2;
  wire       [2:0]    mul3_127_port_byte_out_3;
  wire       [2:0]    mul3_127_port_byte_out_4;
  wire       [2:0]    mul3_127_port_byte_out_5;
  wire       [2:0]    mul3_127_port_byte_out_6;
  wire       [2:0]    mul3_127_port_byte_out_7;
  wire       [2:0]    state_out_0_0_0;
  wire       [2:0]    state_out_0_0_1;
  wire       [2:0]    state_out_0_0_2;
  wire       [2:0]    state_out_0_0_3;
  wire       [2:0]    state_out_0_0_4;
  wire       [2:0]    state_out_0_0_5;
  wire       [2:0]    state_out_0_0_6;
  wire       [2:0]    state_out_0_0_7;
  wire       [2:0]    state_out_0_1_0;
  wire       [2:0]    state_out_0_1_1;
  wire       [2:0]    state_out_0_1_2;
  wire       [2:0]    state_out_0_1_3;
  wire       [2:0]    state_out_0_1_4;
  wire       [2:0]    state_out_0_1_5;
  wire       [2:0]    state_out_0_1_6;
  wire       [2:0]    state_out_0_1_7;
  wire       [2:0]    state_out_0_2_0;
  wire       [2:0]    state_out_0_2_1;
  wire       [2:0]    state_out_0_2_2;
  wire       [2:0]    state_out_0_2_3;
  wire       [2:0]    state_out_0_2_4;
  wire       [2:0]    state_out_0_2_5;
  wire       [2:0]    state_out_0_2_6;
  wire       [2:0]    state_out_0_2_7;
  wire       [2:0]    state_out_0_3_0;
  wire       [2:0]    state_out_0_3_1;
  wire       [2:0]    state_out_0_3_2;
  wire       [2:0]    state_out_0_3_3;
  wire       [2:0]    state_out_0_3_4;
  wire       [2:0]    state_out_0_3_5;
  wire       [2:0]    state_out_0_3_6;
  wire       [2:0]    state_out_0_3_7;
  wire       [2:0]    state_out_1_0_0;
  wire       [2:0]    state_out_1_0_1;
  wire       [2:0]    state_out_1_0_2;
  wire       [2:0]    state_out_1_0_3;
  wire       [2:0]    state_out_1_0_4;
  wire       [2:0]    state_out_1_0_5;
  wire       [2:0]    state_out_1_0_6;
  wire       [2:0]    state_out_1_0_7;
  wire       [2:0]    state_out_1_1_0;
  wire       [2:0]    state_out_1_1_1;
  wire       [2:0]    state_out_1_1_2;
  wire       [2:0]    state_out_1_1_3;
  wire       [2:0]    state_out_1_1_4;
  wire       [2:0]    state_out_1_1_5;
  wire       [2:0]    state_out_1_1_6;
  wire       [2:0]    state_out_1_1_7;
  wire       [2:0]    state_out_1_2_0;
  wire       [2:0]    state_out_1_2_1;
  wire       [2:0]    state_out_1_2_2;
  wire       [2:0]    state_out_1_2_3;
  wire       [2:0]    state_out_1_2_4;
  wire       [2:0]    state_out_1_2_5;
  wire       [2:0]    state_out_1_2_6;
  wire       [2:0]    state_out_1_2_7;
  wire       [2:0]    state_out_1_3_0;
  wire       [2:0]    state_out_1_3_1;
  wire       [2:0]    state_out_1_3_2;
  wire       [2:0]    state_out_1_3_3;
  wire       [2:0]    state_out_1_3_4;
  wire       [2:0]    state_out_1_3_5;
  wire       [2:0]    state_out_1_3_6;
  wire       [2:0]    state_out_1_3_7;
  wire       [2:0]    state_out_2_0_0;
  wire       [2:0]    state_out_2_0_1;
  wire       [2:0]    state_out_2_0_2;
  wire       [2:0]    state_out_2_0_3;
  wire       [2:0]    state_out_2_0_4;
  wire       [2:0]    state_out_2_0_5;
  wire       [2:0]    state_out_2_0_6;
  wire       [2:0]    state_out_2_0_7;
  wire       [2:0]    state_out_2_1_0;
  wire       [2:0]    state_out_2_1_1;
  wire       [2:0]    state_out_2_1_2;
  wire       [2:0]    state_out_2_1_3;
  wire       [2:0]    state_out_2_1_4;
  wire       [2:0]    state_out_2_1_5;
  wire       [2:0]    state_out_2_1_6;
  wire       [2:0]    state_out_2_1_7;
  wire       [2:0]    state_out_2_2_0;
  wire       [2:0]    state_out_2_2_1;
  wire       [2:0]    state_out_2_2_2;
  wire       [2:0]    state_out_2_2_3;
  wire       [2:0]    state_out_2_2_4;
  wire       [2:0]    state_out_2_2_5;
  wire       [2:0]    state_out_2_2_6;
  wire       [2:0]    state_out_2_2_7;
  wire       [2:0]    state_out_2_3_0;
  wire       [2:0]    state_out_2_3_1;
  wire       [2:0]    state_out_2_3_2;
  wire       [2:0]    state_out_2_3_3;
  wire       [2:0]    state_out_2_3_4;
  wire       [2:0]    state_out_2_3_5;
  wire       [2:0]    state_out_2_3_6;
  wire       [2:0]    state_out_2_3_7;
  wire       [2:0]    state_out_3_0_0;
  wire       [2:0]    state_out_3_0_1;
  wire       [2:0]    state_out_3_0_2;
  wire       [2:0]    state_out_3_0_3;
  wire       [2:0]    state_out_3_0_4;
  wire       [2:0]    state_out_3_0_5;
  wire       [2:0]    state_out_3_0_6;
  wire       [2:0]    state_out_3_0_7;
  wire       [2:0]    state_out_3_1_0;
  wire       [2:0]    state_out_3_1_1;
  wire       [2:0]    state_out_3_1_2;
  wire       [2:0]    state_out_3_1_3;
  wire       [2:0]    state_out_3_1_4;
  wire       [2:0]    state_out_3_1_5;
  wire       [2:0]    state_out_3_1_6;
  wire       [2:0]    state_out_3_1_7;
  wire       [2:0]    state_out_3_2_0;
  wire       [2:0]    state_out_3_2_1;
  wire       [2:0]    state_out_3_2_2;
  wire       [2:0]    state_out_3_2_3;
  wire       [2:0]    state_out_3_2_4;
  wire       [2:0]    state_out_3_2_5;
  wire       [2:0]    state_out_3_2_6;
  wire       [2:0]    state_out_3_2_7;
  wire       [2:0]    state_out_3_3_0;
  wire       [2:0]    state_out_3_3_1;
  wire       [2:0]    state_out_3_3_2;
  wire       [2:0]    state_out_3_3_3;
  wire       [2:0]    state_out_3_3_4;
  wire       [2:0]    state_out_3_3_5;
  wire       [2:0]    state_out_3_3_6;
  wire       [2:0]    state_out_3_3_7;
  wire       [2:0]    state_out_4_0_0;
  wire       [2:0]    state_out_4_0_1;
  wire       [2:0]    state_out_4_0_2;
  wire       [2:0]    state_out_4_0_3;
  wire       [2:0]    state_out_4_0_4;
  wire       [2:0]    state_out_4_0_5;
  wire       [2:0]    state_out_4_0_6;
  wire       [2:0]    state_out_4_0_7;
  wire       [2:0]    state_out_4_1_0;
  wire       [2:0]    state_out_4_1_1;
  wire       [2:0]    state_out_4_1_2;
  wire       [2:0]    state_out_4_1_3;
  wire       [2:0]    state_out_4_1_4;
  wire       [2:0]    state_out_4_1_5;
  wire       [2:0]    state_out_4_1_6;
  wire       [2:0]    state_out_4_1_7;
  wire       [2:0]    state_out_4_2_0;
  wire       [2:0]    state_out_4_2_1;
  wire       [2:0]    state_out_4_2_2;
  wire       [2:0]    state_out_4_2_3;
  wire       [2:0]    state_out_4_2_4;
  wire       [2:0]    state_out_4_2_5;
  wire       [2:0]    state_out_4_2_6;
  wire       [2:0]    state_out_4_2_7;
  wire       [2:0]    state_out_4_3_0;
  wire       [2:0]    state_out_4_3_1;
  wire       [2:0]    state_out_4_3_2;
  wire       [2:0]    state_out_4_3_3;
  wire       [2:0]    state_out_4_3_4;
  wire       [2:0]    state_out_4_3_5;
  wire       [2:0]    state_out_4_3_6;
  wire       [2:0]    state_out_4_3_7;
  wire       [2:0]    state_out_5_0_0;
  wire       [2:0]    state_out_5_0_1;
  wire       [2:0]    state_out_5_0_2;
  wire       [2:0]    state_out_5_0_3;
  wire       [2:0]    state_out_5_0_4;
  wire       [2:0]    state_out_5_0_5;
  wire       [2:0]    state_out_5_0_6;
  wire       [2:0]    state_out_5_0_7;
  wire       [2:0]    state_out_5_1_0;
  wire       [2:0]    state_out_5_1_1;
  wire       [2:0]    state_out_5_1_2;
  wire       [2:0]    state_out_5_1_3;
  wire       [2:0]    state_out_5_1_4;
  wire       [2:0]    state_out_5_1_5;
  wire       [2:0]    state_out_5_1_6;
  wire       [2:0]    state_out_5_1_7;
  wire       [2:0]    state_out_5_2_0;
  wire       [2:0]    state_out_5_2_1;
  wire       [2:0]    state_out_5_2_2;
  wire       [2:0]    state_out_5_2_3;
  wire       [2:0]    state_out_5_2_4;
  wire       [2:0]    state_out_5_2_5;
  wire       [2:0]    state_out_5_2_6;
  wire       [2:0]    state_out_5_2_7;
  wire       [2:0]    state_out_5_3_0;
  wire       [2:0]    state_out_5_3_1;
  wire       [2:0]    state_out_5_3_2;
  wire       [2:0]    state_out_5_3_3;
  wire       [2:0]    state_out_5_3_4;
  wire       [2:0]    state_out_5_3_5;
  wire       [2:0]    state_out_5_3_6;
  wire       [2:0]    state_out_5_3_7;
  wire       [2:0]    state_out_6_0_0;
  wire       [2:0]    state_out_6_0_1;
  wire       [2:0]    state_out_6_0_2;
  wire       [2:0]    state_out_6_0_3;
  wire       [2:0]    state_out_6_0_4;
  wire       [2:0]    state_out_6_0_5;
  wire       [2:0]    state_out_6_0_6;
  wire       [2:0]    state_out_6_0_7;
  wire       [2:0]    state_out_6_1_0;
  wire       [2:0]    state_out_6_1_1;
  wire       [2:0]    state_out_6_1_2;
  wire       [2:0]    state_out_6_1_3;
  wire       [2:0]    state_out_6_1_4;
  wire       [2:0]    state_out_6_1_5;
  wire       [2:0]    state_out_6_1_6;
  wire       [2:0]    state_out_6_1_7;
  wire       [2:0]    state_out_6_2_0;
  wire       [2:0]    state_out_6_2_1;
  wire       [2:0]    state_out_6_2_2;
  wire       [2:0]    state_out_6_2_3;
  wire       [2:0]    state_out_6_2_4;
  wire       [2:0]    state_out_6_2_5;
  wire       [2:0]    state_out_6_2_6;
  wire       [2:0]    state_out_6_2_7;
  wire       [2:0]    state_out_6_3_0;
  wire       [2:0]    state_out_6_3_1;
  wire       [2:0]    state_out_6_3_2;
  wire       [2:0]    state_out_6_3_3;
  wire       [2:0]    state_out_6_3_4;
  wire       [2:0]    state_out_6_3_5;
  wire       [2:0]    state_out_6_3_6;
  wire       [2:0]    state_out_6_3_7;
  wire       [2:0]    state_out_7_0_0;
  wire       [2:0]    state_out_7_0_1;
  wire       [2:0]    state_out_7_0_2;
  wire       [2:0]    state_out_7_0_3;
  wire       [2:0]    state_out_7_0_4;
  wire       [2:0]    state_out_7_0_5;
  wire       [2:0]    state_out_7_0_6;
  wire       [2:0]    state_out_7_0_7;
  wire       [2:0]    state_out_7_1_0;
  wire       [2:0]    state_out_7_1_1;
  wire       [2:0]    state_out_7_1_2;
  wire       [2:0]    state_out_7_1_3;
  wire       [2:0]    state_out_7_1_4;
  wire       [2:0]    state_out_7_1_5;
  wire       [2:0]    state_out_7_1_6;
  wire       [2:0]    state_out_7_1_7;
  wire       [2:0]    state_out_7_2_0;
  wire       [2:0]    state_out_7_2_1;
  wire       [2:0]    state_out_7_2_2;
  wire       [2:0]    state_out_7_2_3;
  wire       [2:0]    state_out_7_2_4;
  wire       [2:0]    state_out_7_2_5;
  wire       [2:0]    state_out_7_2_6;
  wire       [2:0]    state_out_7_2_7;
  wire       [2:0]    state_out_7_3_0;
  wire       [2:0]    state_out_7_3_1;
  wire       [2:0]    state_out_7_3_2;
  wire       [2:0]    state_out_7_3_3;
  wire       [2:0]    state_out_7_3_4;
  wire       [2:0]    state_out_7_3_5;
  wire       [2:0]    state_out_7_3_6;
  wire       [2:0]    state_out_7_3_7;
  wire       [2:0]    state_out_8_0_0;
  wire       [2:0]    state_out_8_0_1;
  wire       [2:0]    state_out_8_0_2;
  wire       [2:0]    state_out_8_0_3;
  wire       [2:0]    state_out_8_0_4;
  wire       [2:0]    state_out_8_0_5;
  wire       [2:0]    state_out_8_0_6;
  wire       [2:0]    state_out_8_0_7;
  wire       [2:0]    state_out_8_1_0;
  wire       [2:0]    state_out_8_1_1;
  wire       [2:0]    state_out_8_1_2;
  wire       [2:0]    state_out_8_1_3;
  wire       [2:0]    state_out_8_1_4;
  wire       [2:0]    state_out_8_1_5;
  wire       [2:0]    state_out_8_1_6;
  wire       [2:0]    state_out_8_1_7;
  wire       [2:0]    state_out_8_2_0;
  wire       [2:0]    state_out_8_2_1;
  wire       [2:0]    state_out_8_2_2;
  wire       [2:0]    state_out_8_2_3;
  wire       [2:0]    state_out_8_2_4;
  wire       [2:0]    state_out_8_2_5;
  wire       [2:0]    state_out_8_2_6;
  wire       [2:0]    state_out_8_2_7;
  wire       [2:0]    state_out_8_3_0;
  wire       [2:0]    state_out_8_3_1;
  wire       [2:0]    state_out_8_3_2;
  wire       [2:0]    state_out_8_3_3;
  wire       [2:0]    state_out_8_3_4;
  wire       [2:0]    state_out_8_3_5;
  wire       [2:0]    state_out_8_3_6;
  wire       [2:0]    state_out_8_3_7;
  wire       [2:0]    state_out_9_0_0;
  wire       [2:0]    state_out_9_0_1;
  wire       [2:0]    state_out_9_0_2;
  wire       [2:0]    state_out_9_0_3;
  wire       [2:0]    state_out_9_0_4;
  wire       [2:0]    state_out_9_0_5;
  wire       [2:0]    state_out_9_0_6;
  wire       [2:0]    state_out_9_0_7;
  wire       [2:0]    state_out_9_1_0;
  wire       [2:0]    state_out_9_1_1;
  wire       [2:0]    state_out_9_1_2;
  wire       [2:0]    state_out_9_1_3;
  wire       [2:0]    state_out_9_1_4;
  wire       [2:0]    state_out_9_1_5;
  wire       [2:0]    state_out_9_1_6;
  wire       [2:0]    state_out_9_1_7;
  wire       [2:0]    state_out_9_2_0;
  wire       [2:0]    state_out_9_2_1;
  wire       [2:0]    state_out_9_2_2;
  wire       [2:0]    state_out_9_2_3;
  wire       [2:0]    state_out_9_2_4;
  wire       [2:0]    state_out_9_2_5;
  wire       [2:0]    state_out_9_2_6;
  wire       [2:0]    state_out_9_2_7;
  wire       [2:0]    state_out_9_3_0;
  wire       [2:0]    state_out_9_3_1;
  wire       [2:0]    state_out_9_3_2;
  wire       [2:0]    state_out_9_3_3;
  wire       [2:0]    state_out_9_3_4;
  wire       [2:0]    state_out_9_3_5;
  wire       [2:0]    state_out_9_3_6;
  wire       [2:0]    state_out_9_3_7;
  wire       [2:0]    state_out_10_0_0;
  wire       [2:0]    state_out_10_0_1;
  wire       [2:0]    state_out_10_0_2;
  wire       [2:0]    state_out_10_0_3;
  wire       [2:0]    state_out_10_0_4;
  wire       [2:0]    state_out_10_0_5;
  wire       [2:0]    state_out_10_0_6;
  wire       [2:0]    state_out_10_0_7;
  wire       [2:0]    state_out_10_1_0;
  wire       [2:0]    state_out_10_1_1;
  wire       [2:0]    state_out_10_1_2;
  wire       [2:0]    state_out_10_1_3;
  wire       [2:0]    state_out_10_1_4;
  wire       [2:0]    state_out_10_1_5;
  wire       [2:0]    state_out_10_1_6;
  wire       [2:0]    state_out_10_1_7;
  wire       [2:0]    state_out_10_2_0;
  wire       [2:0]    state_out_10_2_1;
  wire       [2:0]    state_out_10_2_2;
  wire       [2:0]    state_out_10_2_3;
  wire       [2:0]    state_out_10_2_4;
  wire       [2:0]    state_out_10_2_5;
  wire       [2:0]    state_out_10_2_6;
  wire       [2:0]    state_out_10_2_7;
  wire       [2:0]    state_out_10_3_0;
  wire       [2:0]    state_out_10_3_1;
  wire       [2:0]    state_out_10_3_2;
  wire       [2:0]    state_out_10_3_3;
  wire       [2:0]    state_out_10_3_4;
  wire       [2:0]    state_out_10_3_5;
  wire       [2:0]    state_out_10_3_6;
  wire       [2:0]    state_out_10_3_7;
  wire       [2:0]    state_out_11_0_0;
  wire       [2:0]    state_out_11_0_1;
  wire       [2:0]    state_out_11_0_2;
  wire       [2:0]    state_out_11_0_3;
  wire       [2:0]    state_out_11_0_4;
  wire       [2:0]    state_out_11_0_5;
  wire       [2:0]    state_out_11_0_6;
  wire       [2:0]    state_out_11_0_7;
  wire       [2:0]    state_out_11_1_0;
  wire       [2:0]    state_out_11_1_1;
  wire       [2:0]    state_out_11_1_2;
  wire       [2:0]    state_out_11_1_3;
  wire       [2:0]    state_out_11_1_4;
  wire       [2:0]    state_out_11_1_5;
  wire       [2:0]    state_out_11_1_6;
  wire       [2:0]    state_out_11_1_7;
  wire       [2:0]    state_out_11_2_0;
  wire       [2:0]    state_out_11_2_1;
  wire       [2:0]    state_out_11_2_2;
  wire       [2:0]    state_out_11_2_3;
  wire       [2:0]    state_out_11_2_4;
  wire       [2:0]    state_out_11_2_5;
  wire       [2:0]    state_out_11_2_6;
  wire       [2:0]    state_out_11_2_7;
  wire       [2:0]    state_out_11_3_0;
  wire       [2:0]    state_out_11_3_1;
  wire       [2:0]    state_out_11_3_2;
  wire       [2:0]    state_out_11_3_3;
  wire       [2:0]    state_out_11_3_4;
  wire       [2:0]    state_out_11_3_5;
  wire       [2:0]    state_out_11_3_6;
  wire       [2:0]    state_out_11_3_7;
  wire       [2:0]    state_out_12_0_0;
  wire       [2:0]    state_out_12_0_1;
  wire       [2:0]    state_out_12_0_2;
  wire       [2:0]    state_out_12_0_3;
  wire       [2:0]    state_out_12_0_4;
  wire       [2:0]    state_out_12_0_5;
  wire       [2:0]    state_out_12_0_6;
  wire       [2:0]    state_out_12_0_7;
  wire       [2:0]    state_out_12_1_0;
  wire       [2:0]    state_out_12_1_1;
  wire       [2:0]    state_out_12_1_2;
  wire       [2:0]    state_out_12_1_3;
  wire       [2:0]    state_out_12_1_4;
  wire       [2:0]    state_out_12_1_5;
  wire       [2:0]    state_out_12_1_6;
  wire       [2:0]    state_out_12_1_7;
  wire       [2:0]    state_out_12_2_0;
  wire       [2:0]    state_out_12_2_1;
  wire       [2:0]    state_out_12_2_2;
  wire       [2:0]    state_out_12_2_3;
  wire       [2:0]    state_out_12_2_4;
  wire       [2:0]    state_out_12_2_5;
  wire       [2:0]    state_out_12_2_6;
  wire       [2:0]    state_out_12_2_7;
  wire       [2:0]    state_out_12_3_0;
  wire       [2:0]    state_out_12_3_1;
  wire       [2:0]    state_out_12_3_2;
  wire       [2:0]    state_out_12_3_3;
  wire       [2:0]    state_out_12_3_4;
  wire       [2:0]    state_out_12_3_5;
  wire       [2:0]    state_out_12_3_6;
  wire       [2:0]    state_out_12_3_7;
  wire       [2:0]    state_out_13_0_0;
  wire       [2:0]    state_out_13_0_1;
  wire       [2:0]    state_out_13_0_2;
  wire       [2:0]    state_out_13_0_3;
  wire       [2:0]    state_out_13_0_4;
  wire       [2:0]    state_out_13_0_5;
  wire       [2:0]    state_out_13_0_6;
  wire       [2:0]    state_out_13_0_7;
  wire       [2:0]    state_out_13_1_0;
  wire       [2:0]    state_out_13_1_1;
  wire       [2:0]    state_out_13_1_2;
  wire       [2:0]    state_out_13_1_3;
  wire       [2:0]    state_out_13_1_4;
  wire       [2:0]    state_out_13_1_5;
  wire       [2:0]    state_out_13_1_6;
  wire       [2:0]    state_out_13_1_7;
  wire       [2:0]    state_out_13_2_0;
  wire       [2:0]    state_out_13_2_1;
  wire       [2:0]    state_out_13_2_2;
  wire       [2:0]    state_out_13_2_3;
  wire       [2:0]    state_out_13_2_4;
  wire       [2:0]    state_out_13_2_5;
  wire       [2:0]    state_out_13_2_6;
  wire       [2:0]    state_out_13_2_7;
  wire       [2:0]    state_out_13_3_0;
  wire       [2:0]    state_out_13_3_1;
  wire       [2:0]    state_out_13_3_2;
  wire       [2:0]    state_out_13_3_3;
  wire       [2:0]    state_out_13_3_4;
  wire       [2:0]    state_out_13_3_5;
  wire       [2:0]    state_out_13_3_6;
  wire       [2:0]    state_out_13_3_7;
  wire       [2:0]    state_out_14_0_0;
  wire       [2:0]    state_out_14_0_1;
  wire       [2:0]    state_out_14_0_2;
  wire       [2:0]    state_out_14_0_3;
  wire       [2:0]    state_out_14_0_4;
  wire       [2:0]    state_out_14_0_5;
  wire       [2:0]    state_out_14_0_6;
  wire       [2:0]    state_out_14_0_7;
  wire       [2:0]    state_out_14_1_0;
  wire       [2:0]    state_out_14_1_1;
  wire       [2:0]    state_out_14_1_2;
  wire       [2:0]    state_out_14_1_3;
  wire       [2:0]    state_out_14_1_4;
  wire       [2:0]    state_out_14_1_5;
  wire       [2:0]    state_out_14_1_6;
  wire       [2:0]    state_out_14_1_7;
  wire       [2:0]    state_out_14_2_0;
  wire       [2:0]    state_out_14_2_1;
  wire       [2:0]    state_out_14_2_2;
  wire       [2:0]    state_out_14_2_3;
  wire       [2:0]    state_out_14_2_4;
  wire       [2:0]    state_out_14_2_5;
  wire       [2:0]    state_out_14_2_6;
  wire       [2:0]    state_out_14_2_7;
  wire       [2:0]    state_out_14_3_0;
  wire       [2:0]    state_out_14_3_1;
  wire       [2:0]    state_out_14_3_2;
  wire       [2:0]    state_out_14_3_3;
  wire       [2:0]    state_out_14_3_4;
  wire       [2:0]    state_out_14_3_5;
  wire       [2:0]    state_out_14_3_6;
  wire       [2:0]    state_out_14_3_7;
  wire       [2:0]    state_out_15_0_0;
  wire       [2:0]    state_out_15_0_1;
  wire       [2:0]    state_out_15_0_2;
  wire       [2:0]    state_out_15_0_3;
  wire       [2:0]    state_out_15_0_4;
  wire       [2:0]    state_out_15_0_5;
  wire       [2:0]    state_out_15_0_6;
  wire       [2:0]    state_out_15_0_7;
  wire       [2:0]    state_out_15_1_0;
  wire       [2:0]    state_out_15_1_1;
  wire       [2:0]    state_out_15_1_2;
  wire       [2:0]    state_out_15_1_3;
  wire       [2:0]    state_out_15_1_4;
  wire       [2:0]    state_out_15_1_5;
  wire       [2:0]    state_out_15_1_6;
  wire       [2:0]    state_out_15_1_7;
  wire       [2:0]    state_out_15_2_0;
  wire       [2:0]    state_out_15_2_1;
  wire       [2:0]    state_out_15_2_2;
  wire       [2:0]    state_out_15_2_3;
  wire       [2:0]    state_out_15_2_4;
  wire       [2:0]    state_out_15_2_5;
  wire       [2:0]    state_out_15_2_6;
  wire       [2:0]    state_out_15_2_7;
  wire       [2:0]    state_out_15_3_0;
  wire       [2:0]    state_out_15_3_1;
  wire       [2:0]    state_out_15_3_2;
  wire       [2:0]    state_out_15_3_3;
  wire       [2:0]    state_out_15_3_4;
  wire       [2:0]    state_out_15_3_5;
  wire       [2:0]    state_out_15_3_6;
  wire       [2:0]    state_out_15_3_7;

  Mul2 mul2_64 (
    .port_byte_in_0  (port_state_in_0_0_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_0_0_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_0_0_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_0_0_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_0_0_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_0_0_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_0_0_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_0_0_7[2:0]    ), //i
    .port_byte_out_0 (mul2_64_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul2_64_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul2_64_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul2_64_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul2_64_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul2_64_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul2_64_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul2_64_port_byte_out_7[2:0])  //o
  );
  Mul3 mul3_64 (
    .port_byte_in_0  (port_state_in_1_0_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_1_0_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_1_0_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_1_0_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_1_0_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_1_0_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_1_0_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_1_0_7[2:0]    ), //i
    .port_byte_out_0 (mul3_64_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul3_64_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul3_64_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul3_64_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul3_64_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul3_64_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul3_64_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul3_64_port_byte_out_7[2:0])  //o
  );
  Mul2 mul2_65 (
    .port_byte_in_0  (port_state_in_1_0_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_1_0_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_1_0_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_1_0_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_1_0_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_1_0_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_1_0_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_1_0_7[2:0]    ), //i
    .port_byte_out_0 (mul2_65_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul2_65_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul2_65_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul2_65_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul2_65_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul2_65_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul2_65_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul2_65_port_byte_out_7[2:0])  //o
  );
  Mul3 mul3_65 (
    .port_byte_in_0  (port_state_in_2_0_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_2_0_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_2_0_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_2_0_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_2_0_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_2_0_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_2_0_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_2_0_7[2:0]    ), //i
    .port_byte_out_0 (mul3_65_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul3_65_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul3_65_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul3_65_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul3_65_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul3_65_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul3_65_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul3_65_port_byte_out_7[2:0])  //o
  );
  Mul2 mul2_66 (
    .port_byte_in_0  (port_state_in_2_0_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_2_0_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_2_0_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_2_0_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_2_0_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_2_0_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_2_0_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_2_0_7[2:0]    ), //i
    .port_byte_out_0 (mul2_66_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul2_66_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul2_66_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul2_66_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul2_66_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul2_66_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul2_66_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul2_66_port_byte_out_7[2:0])  //o
  );
  Mul3 mul3_66 (
    .port_byte_in_0  (port_state_in_3_0_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_3_0_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_3_0_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_3_0_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_3_0_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_3_0_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_3_0_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_3_0_7[2:0]    ), //i
    .port_byte_out_0 (mul3_66_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul3_66_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul3_66_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul3_66_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul3_66_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul3_66_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul3_66_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul3_66_port_byte_out_7[2:0])  //o
  );
  Mul2 mul2_67 (
    .port_byte_in_0  (port_state_in_3_0_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_3_0_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_3_0_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_3_0_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_3_0_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_3_0_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_3_0_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_3_0_7[2:0]    ), //i
    .port_byte_out_0 (mul2_67_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul2_67_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul2_67_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul2_67_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul2_67_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul2_67_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul2_67_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul2_67_port_byte_out_7[2:0])  //o
  );
  Mul3 mul3_67 (
    .port_byte_in_0  (port_state_in_0_0_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_0_0_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_0_0_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_0_0_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_0_0_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_0_0_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_0_0_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_0_0_7[2:0]    ), //i
    .port_byte_out_0 (mul3_67_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul3_67_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul3_67_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul3_67_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul3_67_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul3_67_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul3_67_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul3_67_port_byte_out_7[2:0])  //o
  );
  Mul2 mul2_68 (
    .port_byte_in_0  (port_state_in_0_1_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_0_1_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_0_1_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_0_1_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_0_1_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_0_1_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_0_1_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_0_1_7[2:0]    ), //i
    .port_byte_out_0 (mul2_68_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul2_68_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul2_68_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul2_68_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul2_68_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul2_68_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul2_68_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul2_68_port_byte_out_7[2:0])  //o
  );
  Mul3 mul3_68 (
    .port_byte_in_0  (port_state_in_1_1_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_1_1_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_1_1_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_1_1_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_1_1_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_1_1_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_1_1_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_1_1_7[2:0]    ), //i
    .port_byte_out_0 (mul3_68_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul3_68_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul3_68_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul3_68_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul3_68_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul3_68_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul3_68_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul3_68_port_byte_out_7[2:0])  //o
  );
  Mul2 mul2_69 (
    .port_byte_in_0  (port_state_in_1_1_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_1_1_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_1_1_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_1_1_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_1_1_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_1_1_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_1_1_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_1_1_7[2:0]    ), //i
    .port_byte_out_0 (mul2_69_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul2_69_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul2_69_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul2_69_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul2_69_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul2_69_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul2_69_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul2_69_port_byte_out_7[2:0])  //o
  );
  Mul3 mul3_69 (
    .port_byte_in_0  (port_state_in_2_1_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_2_1_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_2_1_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_2_1_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_2_1_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_2_1_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_2_1_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_2_1_7[2:0]    ), //i
    .port_byte_out_0 (mul3_69_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul3_69_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul3_69_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul3_69_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul3_69_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul3_69_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul3_69_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul3_69_port_byte_out_7[2:0])  //o
  );
  Mul2 mul2_70 (
    .port_byte_in_0  (port_state_in_2_1_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_2_1_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_2_1_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_2_1_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_2_1_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_2_1_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_2_1_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_2_1_7[2:0]    ), //i
    .port_byte_out_0 (mul2_70_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul2_70_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul2_70_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul2_70_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul2_70_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul2_70_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul2_70_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul2_70_port_byte_out_7[2:0])  //o
  );
  Mul3 mul3_70 (
    .port_byte_in_0  (port_state_in_3_1_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_3_1_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_3_1_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_3_1_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_3_1_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_3_1_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_3_1_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_3_1_7[2:0]    ), //i
    .port_byte_out_0 (mul3_70_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul3_70_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul3_70_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul3_70_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul3_70_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul3_70_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul3_70_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul3_70_port_byte_out_7[2:0])  //o
  );
  Mul2 mul2_71 (
    .port_byte_in_0  (port_state_in_3_1_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_3_1_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_3_1_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_3_1_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_3_1_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_3_1_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_3_1_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_3_1_7[2:0]    ), //i
    .port_byte_out_0 (mul2_71_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul2_71_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul2_71_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul2_71_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul2_71_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul2_71_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul2_71_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul2_71_port_byte_out_7[2:0])  //o
  );
  Mul3 mul3_71 (
    .port_byte_in_0  (port_state_in_0_1_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_0_1_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_0_1_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_0_1_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_0_1_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_0_1_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_0_1_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_0_1_7[2:0]    ), //i
    .port_byte_out_0 (mul3_71_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul3_71_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul3_71_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul3_71_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul3_71_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul3_71_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul3_71_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul3_71_port_byte_out_7[2:0])  //o
  );
  Mul2 mul2_72 (
    .port_byte_in_0  (port_state_in_0_2_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_0_2_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_0_2_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_0_2_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_0_2_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_0_2_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_0_2_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_0_2_7[2:0]    ), //i
    .port_byte_out_0 (mul2_72_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul2_72_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul2_72_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul2_72_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul2_72_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul2_72_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul2_72_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul2_72_port_byte_out_7[2:0])  //o
  );
  Mul3 mul3_72 (
    .port_byte_in_0  (port_state_in_1_2_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_1_2_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_1_2_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_1_2_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_1_2_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_1_2_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_1_2_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_1_2_7[2:0]    ), //i
    .port_byte_out_0 (mul3_72_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul3_72_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul3_72_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul3_72_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul3_72_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul3_72_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul3_72_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul3_72_port_byte_out_7[2:0])  //o
  );
  Mul2 mul2_73 (
    .port_byte_in_0  (port_state_in_1_2_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_1_2_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_1_2_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_1_2_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_1_2_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_1_2_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_1_2_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_1_2_7[2:0]    ), //i
    .port_byte_out_0 (mul2_73_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul2_73_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul2_73_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul2_73_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul2_73_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul2_73_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul2_73_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul2_73_port_byte_out_7[2:0])  //o
  );
  Mul3 mul3_73 (
    .port_byte_in_0  (port_state_in_2_2_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_2_2_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_2_2_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_2_2_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_2_2_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_2_2_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_2_2_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_2_2_7[2:0]    ), //i
    .port_byte_out_0 (mul3_73_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul3_73_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul3_73_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul3_73_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul3_73_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul3_73_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul3_73_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul3_73_port_byte_out_7[2:0])  //o
  );
  Mul2 mul2_74 (
    .port_byte_in_0  (port_state_in_2_2_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_2_2_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_2_2_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_2_2_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_2_2_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_2_2_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_2_2_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_2_2_7[2:0]    ), //i
    .port_byte_out_0 (mul2_74_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul2_74_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul2_74_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul2_74_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul2_74_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul2_74_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul2_74_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul2_74_port_byte_out_7[2:0])  //o
  );
  Mul3 mul3_74 (
    .port_byte_in_0  (port_state_in_3_2_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_3_2_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_3_2_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_3_2_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_3_2_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_3_2_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_3_2_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_3_2_7[2:0]    ), //i
    .port_byte_out_0 (mul3_74_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul3_74_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul3_74_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul3_74_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul3_74_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul3_74_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul3_74_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul3_74_port_byte_out_7[2:0])  //o
  );
  Mul2 mul2_75 (
    .port_byte_in_0  (port_state_in_3_2_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_3_2_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_3_2_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_3_2_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_3_2_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_3_2_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_3_2_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_3_2_7[2:0]    ), //i
    .port_byte_out_0 (mul2_75_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul2_75_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul2_75_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul2_75_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul2_75_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul2_75_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul2_75_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul2_75_port_byte_out_7[2:0])  //o
  );
  Mul3 mul3_75 (
    .port_byte_in_0  (port_state_in_0_2_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_0_2_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_0_2_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_0_2_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_0_2_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_0_2_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_0_2_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_0_2_7[2:0]    ), //i
    .port_byte_out_0 (mul3_75_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul3_75_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul3_75_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul3_75_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul3_75_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul3_75_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul3_75_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul3_75_port_byte_out_7[2:0])  //o
  );
  Mul2 mul2_76 (
    .port_byte_in_0  (port_state_in_0_3_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_0_3_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_0_3_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_0_3_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_0_3_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_0_3_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_0_3_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_0_3_7[2:0]    ), //i
    .port_byte_out_0 (mul2_76_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul2_76_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul2_76_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul2_76_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul2_76_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul2_76_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul2_76_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul2_76_port_byte_out_7[2:0])  //o
  );
  Mul3 mul3_76 (
    .port_byte_in_0  (port_state_in_1_3_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_1_3_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_1_3_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_1_3_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_1_3_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_1_3_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_1_3_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_1_3_7[2:0]    ), //i
    .port_byte_out_0 (mul3_76_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul3_76_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul3_76_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul3_76_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul3_76_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul3_76_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul3_76_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul3_76_port_byte_out_7[2:0])  //o
  );
  Mul2 mul2_77 (
    .port_byte_in_0  (port_state_in_1_3_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_1_3_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_1_3_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_1_3_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_1_3_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_1_3_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_1_3_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_1_3_7[2:0]    ), //i
    .port_byte_out_0 (mul2_77_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul2_77_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul2_77_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul2_77_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul2_77_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul2_77_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul2_77_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul2_77_port_byte_out_7[2:0])  //o
  );
  Mul3 mul3_77 (
    .port_byte_in_0  (port_state_in_2_3_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_2_3_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_2_3_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_2_3_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_2_3_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_2_3_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_2_3_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_2_3_7[2:0]    ), //i
    .port_byte_out_0 (mul3_77_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul3_77_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul3_77_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul3_77_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul3_77_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul3_77_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul3_77_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul3_77_port_byte_out_7[2:0])  //o
  );
  Mul2 mul2_78 (
    .port_byte_in_0  (port_state_in_2_3_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_2_3_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_2_3_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_2_3_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_2_3_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_2_3_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_2_3_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_2_3_7[2:0]    ), //i
    .port_byte_out_0 (mul2_78_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul2_78_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul2_78_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul2_78_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul2_78_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul2_78_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul2_78_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul2_78_port_byte_out_7[2:0])  //o
  );
  Mul3 mul3_78 (
    .port_byte_in_0  (port_state_in_3_3_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_3_3_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_3_3_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_3_3_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_3_3_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_3_3_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_3_3_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_3_3_7[2:0]    ), //i
    .port_byte_out_0 (mul3_78_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul3_78_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul3_78_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul3_78_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul3_78_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul3_78_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul3_78_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul3_78_port_byte_out_7[2:0])  //o
  );
  Mul2 mul2_79 (
    .port_byte_in_0  (port_state_in_3_3_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_3_3_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_3_3_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_3_3_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_3_3_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_3_3_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_3_3_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_3_3_7[2:0]    ), //i
    .port_byte_out_0 (mul2_79_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul2_79_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul2_79_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul2_79_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul2_79_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul2_79_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul2_79_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul2_79_port_byte_out_7[2:0])  //o
  );
  Mul3 mul3_79 (
    .port_byte_in_0  (port_state_in_0_3_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_0_3_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_0_3_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_0_3_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_0_3_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_0_3_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_0_3_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_0_3_7[2:0]    ), //i
    .port_byte_out_0 (mul3_79_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul3_79_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul3_79_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul3_79_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul3_79_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul3_79_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul3_79_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul3_79_port_byte_out_7[2:0])  //o
  );
  Mul2 mul2_80 (
    .port_byte_in_0  (port_state_in_4_0_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_4_0_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_4_0_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_4_0_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_4_0_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_4_0_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_4_0_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_4_0_7[2:0]    ), //i
    .port_byte_out_0 (mul2_80_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul2_80_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul2_80_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul2_80_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul2_80_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul2_80_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul2_80_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul2_80_port_byte_out_7[2:0])  //o
  );
  Mul3 mul3_80 (
    .port_byte_in_0  (port_state_in_5_0_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_5_0_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_5_0_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_5_0_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_5_0_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_5_0_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_5_0_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_5_0_7[2:0]    ), //i
    .port_byte_out_0 (mul3_80_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul3_80_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul3_80_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul3_80_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul3_80_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul3_80_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul3_80_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul3_80_port_byte_out_7[2:0])  //o
  );
  Mul2 mul2_81 (
    .port_byte_in_0  (port_state_in_5_0_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_5_0_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_5_0_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_5_0_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_5_0_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_5_0_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_5_0_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_5_0_7[2:0]    ), //i
    .port_byte_out_0 (mul2_81_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul2_81_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul2_81_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul2_81_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul2_81_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul2_81_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul2_81_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul2_81_port_byte_out_7[2:0])  //o
  );
  Mul3 mul3_81 (
    .port_byte_in_0  (port_state_in_6_0_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_6_0_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_6_0_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_6_0_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_6_0_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_6_0_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_6_0_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_6_0_7[2:0]    ), //i
    .port_byte_out_0 (mul3_81_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul3_81_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul3_81_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul3_81_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul3_81_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul3_81_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul3_81_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul3_81_port_byte_out_7[2:0])  //o
  );
  Mul2 mul2_82 (
    .port_byte_in_0  (port_state_in_6_0_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_6_0_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_6_0_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_6_0_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_6_0_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_6_0_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_6_0_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_6_0_7[2:0]    ), //i
    .port_byte_out_0 (mul2_82_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul2_82_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul2_82_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul2_82_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul2_82_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul2_82_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul2_82_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul2_82_port_byte_out_7[2:0])  //o
  );
  Mul3 mul3_82 (
    .port_byte_in_0  (port_state_in_7_0_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_7_0_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_7_0_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_7_0_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_7_0_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_7_0_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_7_0_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_7_0_7[2:0]    ), //i
    .port_byte_out_0 (mul3_82_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul3_82_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul3_82_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul3_82_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul3_82_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul3_82_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul3_82_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul3_82_port_byte_out_7[2:0])  //o
  );
  Mul2 mul2_83 (
    .port_byte_in_0  (port_state_in_7_0_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_7_0_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_7_0_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_7_0_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_7_0_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_7_0_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_7_0_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_7_0_7[2:0]    ), //i
    .port_byte_out_0 (mul2_83_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul2_83_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul2_83_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul2_83_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul2_83_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul2_83_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul2_83_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul2_83_port_byte_out_7[2:0])  //o
  );
  Mul3 mul3_83 (
    .port_byte_in_0  (port_state_in_4_0_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_4_0_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_4_0_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_4_0_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_4_0_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_4_0_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_4_0_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_4_0_7[2:0]    ), //i
    .port_byte_out_0 (mul3_83_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul3_83_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul3_83_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul3_83_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul3_83_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul3_83_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul3_83_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul3_83_port_byte_out_7[2:0])  //o
  );
  Mul2 mul2_84 (
    .port_byte_in_0  (port_state_in_4_1_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_4_1_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_4_1_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_4_1_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_4_1_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_4_1_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_4_1_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_4_1_7[2:0]    ), //i
    .port_byte_out_0 (mul2_84_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul2_84_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul2_84_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul2_84_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul2_84_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul2_84_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul2_84_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul2_84_port_byte_out_7[2:0])  //o
  );
  Mul3 mul3_84 (
    .port_byte_in_0  (port_state_in_5_1_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_5_1_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_5_1_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_5_1_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_5_1_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_5_1_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_5_1_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_5_1_7[2:0]    ), //i
    .port_byte_out_0 (mul3_84_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul3_84_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul3_84_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul3_84_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul3_84_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul3_84_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul3_84_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul3_84_port_byte_out_7[2:0])  //o
  );
  Mul2 mul2_85 (
    .port_byte_in_0  (port_state_in_5_1_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_5_1_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_5_1_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_5_1_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_5_1_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_5_1_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_5_1_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_5_1_7[2:0]    ), //i
    .port_byte_out_0 (mul2_85_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul2_85_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul2_85_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul2_85_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul2_85_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul2_85_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul2_85_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul2_85_port_byte_out_7[2:0])  //o
  );
  Mul3 mul3_85 (
    .port_byte_in_0  (port_state_in_6_1_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_6_1_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_6_1_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_6_1_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_6_1_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_6_1_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_6_1_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_6_1_7[2:0]    ), //i
    .port_byte_out_0 (mul3_85_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul3_85_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul3_85_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul3_85_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul3_85_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul3_85_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul3_85_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul3_85_port_byte_out_7[2:0])  //o
  );
  Mul2 mul2_86 (
    .port_byte_in_0  (port_state_in_6_1_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_6_1_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_6_1_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_6_1_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_6_1_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_6_1_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_6_1_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_6_1_7[2:0]    ), //i
    .port_byte_out_0 (mul2_86_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul2_86_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul2_86_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul2_86_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul2_86_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul2_86_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul2_86_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul2_86_port_byte_out_7[2:0])  //o
  );
  Mul3 mul3_86 (
    .port_byte_in_0  (port_state_in_7_1_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_7_1_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_7_1_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_7_1_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_7_1_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_7_1_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_7_1_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_7_1_7[2:0]    ), //i
    .port_byte_out_0 (mul3_86_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul3_86_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul3_86_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul3_86_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul3_86_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul3_86_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul3_86_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul3_86_port_byte_out_7[2:0])  //o
  );
  Mul2 mul2_87 (
    .port_byte_in_0  (port_state_in_7_1_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_7_1_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_7_1_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_7_1_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_7_1_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_7_1_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_7_1_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_7_1_7[2:0]    ), //i
    .port_byte_out_0 (mul2_87_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul2_87_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul2_87_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul2_87_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul2_87_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul2_87_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul2_87_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul2_87_port_byte_out_7[2:0])  //o
  );
  Mul3 mul3_87 (
    .port_byte_in_0  (port_state_in_4_1_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_4_1_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_4_1_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_4_1_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_4_1_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_4_1_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_4_1_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_4_1_7[2:0]    ), //i
    .port_byte_out_0 (mul3_87_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul3_87_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul3_87_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul3_87_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul3_87_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul3_87_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul3_87_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul3_87_port_byte_out_7[2:0])  //o
  );
  Mul2 mul2_88 (
    .port_byte_in_0  (port_state_in_4_2_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_4_2_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_4_2_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_4_2_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_4_2_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_4_2_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_4_2_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_4_2_7[2:0]    ), //i
    .port_byte_out_0 (mul2_88_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul2_88_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul2_88_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul2_88_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul2_88_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul2_88_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul2_88_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul2_88_port_byte_out_7[2:0])  //o
  );
  Mul3 mul3_88 (
    .port_byte_in_0  (port_state_in_5_2_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_5_2_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_5_2_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_5_2_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_5_2_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_5_2_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_5_2_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_5_2_7[2:0]    ), //i
    .port_byte_out_0 (mul3_88_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul3_88_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul3_88_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul3_88_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul3_88_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul3_88_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul3_88_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul3_88_port_byte_out_7[2:0])  //o
  );
  Mul2 mul2_89 (
    .port_byte_in_0  (port_state_in_5_2_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_5_2_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_5_2_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_5_2_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_5_2_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_5_2_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_5_2_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_5_2_7[2:0]    ), //i
    .port_byte_out_0 (mul2_89_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul2_89_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul2_89_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul2_89_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul2_89_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul2_89_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul2_89_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul2_89_port_byte_out_7[2:0])  //o
  );
  Mul3 mul3_89 (
    .port_byte_in_0  (port_state_in_6_2_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_6_2_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_6_2_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_6_2_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_6_2_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_6_2_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_6_2_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_6_2_7[2:0]    ), //i
    .port_byte_out_0 (mul3_89_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul3_89_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul3_89_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul3_89_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul3_89_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul3_89_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul3_89_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul3_89_port_byte_out_7[2:0])  //o
  );
  Mul2 mul2_90 (
    .port_byte_in_0  (port_state_in_6_2_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_6_2_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_6_2_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_6_2_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_6_2_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_6_2_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_6_2_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_6_2_7[2:0]    ), //i
    .port_byte_out_0 (mul2_90_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul2_90_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul2_90_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul2_90_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul2_90_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul2_90_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul2_90_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul2_90_port_byte_out_7[2:0])  //o
  );
  Mul3 mul3_90 (
    .port_byte_in_0  (port_state_in_7_2_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_7_2_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_7_2_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_7_2_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_7_2_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_7_2_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_7_2_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_7_2_7[2:0]    ), //i
    .port_byte_out_0 (mul3_90_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul3_90_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul3_90_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul3_90_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul3_90_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul3_90_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul3_90_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul3_90_port_byte_out_7[2:0])  //o
  );
  Mul2 mul2_91 (
    .port_byte_in_0  (port_state_in_7_2_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_7_2_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_7_2_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_7_2_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_7_2_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_7_2_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_7_2_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_7_2_7[2:0]    ), //i
    .port_byte_out_0 (mul2_91_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul2_91_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul2_91_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul2_91_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul2_91_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul2_91_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul2_91_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul2_91_port_byte_out_7[2:0])  //o
  );
  Mul3 mul3_91 (
    .port_byte_in_0  (port_state_in_4_2_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_4_2_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_4_2_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_4_2_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_4_2_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_4_2_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_4_2_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_4_2_7[2:0]    ), //i
    .port_byte_out_0 (mul3_91_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul3_91_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul3_91_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul3_91_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul3_91_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul3_91_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul3_91_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul3_91_port_byte_out_7[2:0])  //o
  );
  Mul2 mul2_92 (
    .port_byte_in_0  (port_state_in_4_3_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_4_3_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_4_3_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_4_3_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_4_3_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_4_3_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_4_3_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_4_3_7[2:0]    ), //i
    .port_byte_out_0 (mul2_92_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul2_92_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul2_92_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul2_92_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul2_92_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul2_92_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul2_92_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul2_92_port_byte_out_7[2:0])  //o
  );
  Mul3 mul3_92 (
    .port_byte_in_0  (port_state_in_5_3_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_5_3_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_5_3_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_5_3_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_5_3_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_5_3_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_5_3_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_5_3_7[2:0]    ), //i
    .port_byte_out_0 (mul3_92_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul3_92_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul3_92_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul3_92_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul3_92_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul3_92_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul3_92_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul3_92_port_byte_out_7[2:0])  //o
  );
  Mul2 mul2_93 (
    .port_byte_in_0  (port_state_in_5_3_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_5_3_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_5_3_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_5_3_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_5_3_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_5_3_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_5_3_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_5_3_7[2:0]    ), //i
    .port_byte_out_0 (mul2_93_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul2_93_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul2_93_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul2_93_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul2_93_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul2_93_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul2_93_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul2_93_port_byte_out_7[2:0])  //o
  );
  Mul3 mul3_93 (
    .port_byte_in_0  (port_state_in_6_3_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_6_3_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_6_3_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_6_3_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_6_3_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_6_3_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_6_3_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_6_3_7[2:0]    ), //i
    .port_byte_out_0 (mul3_93_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul3_93_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul3_93_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul3_93_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul3_93_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul3_93_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul3_93_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul3_93_port_byte_out_7[2:0])  //o
  );
  Mul2 mul2_94 (
    .port_byte_in_0  (port_state_in_6_3_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_6_3_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_6_3_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_6_3_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_6_3_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_6_3_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_6_3_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_6_3_7[2:0]    ), //i
    .port_byte_out_0 (mul2_94_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul2_94_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul2_94_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul2_94_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul2_94_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul2_94_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul2_94_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul2_94_port_byte_out_7[2:0])  //o
  );
  Mul3 mul3_94 (
    .port_byte_in_0  (port_state_in_7_3_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_7_3_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_7_3_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_7_3_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_7_3_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_7_3_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_7_3_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_7_3_7[2:0]    ), //i
    .port_byte_out_0 (mul3_94_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul3_94_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul3_94_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul3_94_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul3_94_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul3_94_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul3_94_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul3_94_port_byte_out_7[2:0])  //o
  );
  Mul2 mul2_95 (
    .port_byte_in_0  (port_state_in_7_3_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_7_3_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_7_3_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_7_3_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_7_3_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_7_3_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_7_3_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_7_3_7[2:0]    ), //i
    .port_byte_out_0 (mul2_95_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul2_95_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul2_95_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul2_95_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul2_95_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul2_95_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul2_95_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul2_95_port_byte_out_7[2:0])  //o
  );
  Mul3 mul3_95 (
    .port_byte_in_0  (port_state_in_4_3_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_4_3_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_4_3_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_4_3_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_4_3_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_4_3_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_4_3_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_4_3_7[2:0]    ), //i
    .port_byte_out_0 (mul3_95_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul3_95_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul3_95_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul3_95_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul3_95_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul3_95_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul3_95_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul3_95_port_byte_out_7[2:0])  //o
  );
  Mul2 mul2_96 (
    .port_byte_in_0  (port_state_in_8_0_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_8_0_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_8_0_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_8_0_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_8_0_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_8_0_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_8_0_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_8_0_7[2:0]    ), //i
    .port_byte_out_0 (mul2_96_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul2_96_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul2_96_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul2_96_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul2_96_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul2_96_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul2_96_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul2_96_port_byte_out_7[2:0])  //o
  );
  Mul3 mul3_96 (
    .port_byte_in_0  (port_state_in_9_0_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_9_0_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_9_0_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_9_0_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_9_0_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_9_0_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_9_0_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_9_0_7[2:0]    ), //i
    .port_byte_out_0 (mul3_96_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul3_96_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul3_96_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul3_96_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul3_96_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul3_96_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul3_96_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul3_96_port_byte_out_7[2:0])  //o
  );
  Mul2 mul2_97 (
    .port_byte_in_0  (port_state_in_9_0_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_9_0_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_9_0_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_9_0_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_9_0_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_9_0_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_9_0_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_9_0_7[2:0]    ), //i
    .port_byte_out_0 (mul2_97_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul2_97_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul2_97_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul2_97_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul2_97_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul2_97_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul2_97_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul2_97_port_byte_out_7[2:0])  //o
  );
  Mul3 mul3_97 (
    .port_byte_in_0  (port_state_in_10_0_0[2:0]   ), //i
    .port_byte_in_1  (port_state_in_10_0_1[2:0]   ), //i
    .port_byte_in_2  (port_state_in_10_0_2[2:0]   ), //i
    .port_byte_in_3  (port_state_in_10_0_3[2:0]   ), //i
    .port_byte_in_4  (port_state_in_10_0_4[2:0]   ), //i
    .port_byte_in_5  (port_state_in_10_0_5[2:0]   ), //i
    .port_byte_in_6  (port_state_in_10_0_6[2:0]   ), //i
    .port_byte_in_7  (port_state_in_10_0_7[2:0]   ), //i
    .port_byte_out_0 (mul3_97_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul3_97_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul3_97_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul3_97_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul3_97_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul3_97_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul3_97_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul3_97_port_byte_out_7[2:0])  //o
  );
  Mul2 mul2_98 (
    .port_byte_in_0  (port_state_in_10_0_0[2:0]   ), //i
    .port_byte_in_1  (port_state_in_10_0_1[2:0]   ), //i
    .port_byte_in_2  (port_state_in_10_0_2[2:0]   ), //i
    .port_byte_in_3  (port_state_in_10_0_3[2:0]   ), //i
    .port_byte_in_4  (port_state_in_10_0_4[2:0]   ), //i
    .port_byte_in_5  (port_state_in_10_0_5[2:0]   ), //i
    .port_byte_in_6  (port_state_in_10_0_6[2:0]   ), //i
    .port_byte_in_7  (port_state_in_10_0_7[2:0]   ), //i
    .port_byte_out_0 (mul2_98_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul2_98_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul2_98_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul2_98_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul2_98_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul2_98_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul2_98_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul2_98_port_byte_out_7[2:0])  //o
  );
  Mul3 mul3_98 (
    .port_byte_in_0  (port_state_in_11_0_0[2:0]   ), //i
    .port_byte_in_1  (port_state_in_11_0_1[2:0]   ), //i
    .port_byte_in_2  (port_state_in_11_0_2[2:0]   ), //i
    .port_byte_in_3  (port_state_in_11_0_3[2:0]   ), //i
    .port_byte_in_4  (port_state_in_11_0_4[2:0]   ), //i
    .port_byte_in_5  (port_state_in_11_0_5[2:0]   ), //i
    .port_byte_in_6  (port_state_in_11_0_6[2:0]   ), //i
    .port_byte_in_7  (port_state_in_11_0_7[2:0]   ), //i
    .port_byte_out_0 (mul3_98_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul3_98_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul3_98_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul3_98_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul3_98_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul3_98_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul3_98_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul3_98_port_byte_out_7[2:0])  //o
  );
  Mul2 mul2_99 (
    .port_byte_in_0  (port_state_in_11_0_0[2:0]   ), //i
    .port_byte_in_1  (port_state_in_11_0_1[2:0]   ), //i
    .port_byte_in_2  (port_state_in_11_0_2[2:0]   ), //i
    .port_byte_in_3  (port_state_in_11_0_3[2:0]   ), //i
    .port_byte_in_4  (port_state_in_11_0_4[2:0]   ), //i
    .port_byte_in_5  (port_state_in_11_0_5[2:0]   ), //i
    .port_byte_in_6  (port_state_in_11_0_6[2:0]   ), //i
    .port_byte_in_7  (port_state_in_11_0_7[2:0]   ), //i
    .port_byte_out_0 (mul2_99_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul2_99_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul2_99_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul2_99_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul2_99_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul2_99_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul2_99_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul2_99_port_byte_out_7[2:0])  //o
  );
  Mul3 mul3_99 (
    .port_byte_in_0  (port_state_in_8_0_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_8_0_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_8_0_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_8_0_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_8_0_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_8_0_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_8_0_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_8_0_7[2:0]    ), //i
    .port_byte_out_0 (mul3_99_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul3_99_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul3_99_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul3_99_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul3_99_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul3_99_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul3_99_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul3_99_port_byte_out_7[2:0])  //o
  );
  Mul2 mul2_100 (
    .port_byte_in_0  (port_state_in_8_1_0[2:0]     ), //i
    .port_byte_in_1  (port_state_in_8_1_1[2:0]     ), //i
    .port_byte_in_2  (port_state_in_8_1_2[2:0]     ), //i
    .port_byte_in_3  (port_state_in_8_1_3[2:0]     ), //i
    .port_byte_in_4  (port_state_in_8_1_4[2:0]     ), //i
    .port_byte_in_5  (port_state_in_8_1_5[2:0]     ), //i
    .port_byte_in_6  (port_state_in_8_1_6[2:0]     ), //i
    .port_byte_in_7  (port_state_in_8_1_7[2:0]     ), //i
    .port_byte_out_0 (mul2_100_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul2_100_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul2_100_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul2_100_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul2_100_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul2_100_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul2_100_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul2_100_port_byte_out_7[2:0])  //o
  );
  Mul3 mul3_100 (
    .port_byte_in_0  (port_state_in_9_1_0[2:0]     ), //i
    .port_byte_in_1  (port_state_in_9_1_1[2:0]     ), //i
    .port_byte_in_2  (port_state_in_9_1_2[2:0]     ), //i
    .port_byte_in_3  (port_state_in_9_1_3[2:0]     ), //i
    .port_byte_in_4  (port_state_in_9_1_4[2:0]     ), //i
    .port_byte_in_5  (port_state_in_9_1_5[2:0]     ), //i
    .port_byte_in_6  (port_state_in_9_1_6[2:0]     ), //i
    .port_byte_in_7  (port_state_in_9_1_7[2:0]     ), //i
    .port_byte_out_0 (mul3_100_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul3_100_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul3_100_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul3_100_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul3_100_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul3_100_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul3_100_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul3_100_port_byte_out_7[2:0])  //o
  );
  Mul2 mul2_101 (
    .port_byte_in_0  (port_state_in_9_1_0[2:0]     ), //i
    .port_byte_in_1  (port_state_in_9_1_1[2:0]     ), //i
    .port_byte_in_2  (port_state_in_9_1_2[2:0]     ), //i
    .port_byte_in_3  (port_state_in_9_1_3[2:0]     ), //i
    .port_byte_in_4  (port_state_in_9_1_4[2:0]     ), //i
    .port_byte_in_5  (port_state_in_9_1_5[2:0]     ), //i
    .port_byte_in_6  (port_state_in_9_1_6[2:0]     ), //i
    .port_byte_in_7  (port_state_in_9_1_7[2:0]     ), //i
    .port_byte_out_0 (mul2_101_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul2_101_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul2_101_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul2_101_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul2_101_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul2_101_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul2_101_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul2_101_port_byte_out_7[2:0])  //o
  );
  Mul3 mul3_101 (
    .port_byte_in_0  (port_state_in_10_1_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_10_1_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_10_1_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_10_1_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_10_1_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_10_1_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_10_1_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_10_1_7[2:0]    ), //i
    .port_byte_out_0 (mul3_101_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul3_101_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul3_101_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul3_101_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul3_101_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul3_101_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul3_101_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul3_101_port_byte_out_7[2:0])  //o
  );
  Mul2 mul2_102 (
    .port_byte_in_0  (port_state_in_10_1_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_10_1_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_10_1_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_10_1_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_10_1_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_10_1_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_10_1_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_10_1_7[2:0]    ), //i
    .port_byte_out_0 (mul2_102_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul2_102_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul2_102_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul2_102_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul2_102_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul2_102_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul2_102_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul2_102_port_byte_out_7[2:0])  //o
  );
  Mul3 mul3_102 (
    .port_byte_in_0  (port_state_in_11_1_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_11_1_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_11_1_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_11_1_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_11_1_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_11_1_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_11_1_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_11_1_7[2:0]    ), //i
    .port_byte_out_0 (mul3_102_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul3_102_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul3_102_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul3_102_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul3_102_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul3_102_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul3_102_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul3_102_port_byte_out_7[2:0])  //o
  );
  Mul2 mul2_103 (
    .port_byte_in_0  (port_state_in_11_1_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_11_1_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_11_1_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_11_1_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_11_1_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_11_1_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_11_1_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_11_1_7[2:0]    ), //i
    .port_byte_out_0 (mul2_103_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul2_103_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul2_103_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul2_103_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul2_103_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul2_103_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul2_103_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul2_103_port_byte_out_7[2:0])  //o
  );
  Mul3 mul3_103 (
    .port_byte_in_0  (port_state_in_8_1_0[2:0]     ), //i
    .port_byte_in_1  (port_state_in_8_1_1[2:0]     ), //i
    .port_byte_in_2  (port_state_in_8_1_2[2:0]     ), //i
    .port_byte_in_3  (port_state_in_8_1_3[2:0]     ), //i
    .port_byte_in_4  (port_state_in_8_1_4[2:0]     ), //i
    .port_byte_in_5  (port_state_in_8_1_5[2:0]     ), //i
    .port_byte_in_6  (port_state_in_8_1_6[2:0]     ), //i
    .port_byte_in_7  (port_state_in_8_1_7[2:0]     ), //i
    .port_byte_out_0 (mul3_103_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul3_103_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul3_103_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul3_103_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul3_103_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul3_103_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul3_103_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul3_103_port_byte_out_7[2:0])  //o
  );
  Mul2 mul2_104 (
    .port_byte_in_0  (port_state_in_8_2_0[2:0]     ), //i
    .port_byte_in_1  (port_state_in_8_2_1[2:0]     ), //i
    .port_byte_in_2  (port_state_in_8_2_2[2:0]     ), //i
    .port_byte_in_3  (port_state_in_8_2_3[2:0]     ), //i
    .port_byte_in_4  (port_state_in_8_2_4[2:0]     ), //i
    .port_byte_in_5  (port_state_in_8_2_5[2:0]     ), //i
    .port_byte_in_6  (port_state_in_8_2_6[2:0]     ), //i
    .port_byte_in_7  (port_state_in_8_2_7[2:0]     ), //i
    .port_byte_out_0 (mul2_104_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul2_104_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul2_104_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul2_104_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul2_104_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul2_104_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul2_104_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul2_104_port_byte_out_7[2:0])  //o
  );
  Mul3 mul3_104 (
    .port_byte_in_0  (port_state_in_9_2_0[2:0]     ), //i
    .port_byte_in_1  (port_state_in_9_2_1[2:0]     ), //i
    .port_byte_in_2  (port_state_in_9_2_2[2:0]     ), //i
    .port_byte_in_3  (port_state_in_9_2_3[2:0]     ), //i
    .port_byte_in_4  (port_state_in_9_2_4[2:0]     ), //i
    .port_byte_in_5  (port_state_in_9_2_5[2:0]     ), //i
    .port_byte_in_6  (port_state_in_9_2_6[2:0]     ), //i
    .port_byte_in_7  (port_state_in_9_2_7[2:0]     ), //i
    .port_byte_out_0 (mul3_104_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul3_104_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul3_104_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul3_104_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul3_104_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul3_104_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul3_104_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul3_104_port_byte_out_7[2:0])  //o
  );
  Mul2 mul2_105 (
    .port_byte_in_0  (port_state_in_9_2_0[2:0]     ), //i
    .port_byte_in_1  (port_state_in_9_2_1[2:0]     ), //i
    .port_byte_in_2  (port_state_in_9_2_2[2:0]     ), //i
    .port_byte_in_3  (port_state_in_9_2_3[2:0]     ), //i
    .port_byte_in_4  (port_state_in_9_2_4[2:0]     ), //i
    .port_byte_in_5  (port_state_in_9_2_5[2:0]     ), //i
    .port_byte_in_6  (port_state_in_9_2_6[2:0]     ), //i
    .port_byte_in_7  (port_state_in_9_2_7[2:0]     ), //i
    .port_byte_out_0 (mul2_105_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul2_105_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul2_105_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul2_105_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul2_105_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul2_105_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul2_105_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul2_105_port_byte_out_7[2:0])  //o
  );
  Mul3 mul3_105 (
    .port_byte_in_0  (port_state_in_10_2_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_10_2_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_10_2_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_10_2_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_10_2_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_10_2_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_10_2_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_10_2_7[2:0]    ), //i
    .port_byte_out_0 (mul3_105_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul3_105_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul3_105_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul3_105_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul3_105_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul3_105_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul3_105_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul3_105_port_byte_out_7[2:0])  //o
  );
  Mul2 mul2_106 (
    .port_byte_in_0  (port_state_in_10_2_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_10_2_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_10_2_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_10_2_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_10_2_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_10_2_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_10_2_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_10_2_7[2:0]    ), //i
    .port_byte_out_0 (mul2_106_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul2_106_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul2_106_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul2_106_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul2_106_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul2_106_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul2_106_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul2_106_port_byte_out_7[2:0])  //o
  );
  Mul3 mul3_106 (
    .port_byte_in_0  (port_state_in_11_2_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_11_2_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_11_2_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_11_2_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_11_2_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_11_2_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_11_2_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_11_2_7[2:0]    ), //i
    .port_byte_out_0 (mul3_106_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul3_106_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul3_106_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul3_106_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul3_106_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul3_106_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul3_106_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul3_106_port_byte_out_7[2:0])  //o
  );
  Mul2 mul2_107 (
    .port_byte_in_0  (port_state_in_11_2_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_11_2_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_11_2_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_11_2_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_11_2_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_11_2_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_11_2_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_11_2_7[2:0]    ), //i
    .port_byte_out_0 (mul2_107_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul2_107_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul2_107_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul2_107_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul2_107_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul2_107_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul2_107_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul2_107_port_byte_out_7[2:0])  //o
  );
  Mul3 mul3_107 (
    .port_byte_in_0  (port_state_in_8_2_0[2:0]     ), //i
    .port_byte_in_1  (port_state_in_8_2_1[2:0]     ), //i
    .port_byte_in_2  (port_state_in_8_2_2[2:0]     ), //i
    .port_byte_in_3  (port_state_in_8_2_3[2:0]     ), //i
    .port_byte_in_4  (port_state_in_8_2_4[2:0]     ), //i
    .port_byte_in_5  (port_state_in_8_2_5[2:0]     ), //i
    .port_byte_in_6  (port_state_in_8_2_6[2:0]     ), //i
    .port_byte_in_7  (port_state_in_8_2_7[2:0]     ), //i
    .port_byte_out_0 (mul3_107_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul3_107_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul3_107_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul3_107_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul3_107_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul3_107_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul3_107_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul3_107_port_byte_out_7[2:0])  //o
  );
  Mul2 mul2_108 (
    .port_byte_in_0  (port_state_in_8_3_0[2:0]     ), //i
    .port_byte_in_1  (port_state_in_8_3_1[2:0]     ), //i
    .port_byte_in_2  (port_state_in_8_3_2[2:0]     ), //i
    .port_byte_in_3  (port_state_in_8_3_3[2:0]     ), //i
    .port_byte_in_4  (port_state_in_8_3_4[2:0]     ), //i
    .port_byte_in_5  (port_state_in_8_3_5[2:0]     ), //i
    .port_byte_in_6  (port_state_in_8_3_6[2:0]     ), //i
    .port_byte_in_7  (port_state_in_8_3_7[2:0]     ), //i
    .port_byte_out_0 (mul2_108_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul2_108_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul2_108_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul2_108_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul2_108_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul2_108_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul2_108_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul2_108_port_byte_out_7[2:0])  //o
  );
  Mul3 mul3_108 (
    .port_byte_in_0  (port_state_in_9_3_0[2:0]     ), //i
    .port_byte_in_1  (port_state_in_9_3_1[2:0]     ), //i
    .port_byte_in_2  (port_state_in_9_3_2[2:0]     ), //i
    .port_byte_in_3  (port_state_in_9_3_3[2:0]     ), //i
    .port_byte_in_4  (port_state_in_9_3_4[2:0]     ), //i
    .port_byte_in_5  (port_state_in_9_3_5[2:0]     ), //i
    .port_byte_in_6  (port_state_in_9_3_6[2:0]     ), //i
    .port_byte_in_7  (port_state_in_9_3_7[2:0]     ), //i
    .port_byte_out_0 (mul3_108_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul3_108_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul3_108_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul3_108_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul3_108_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul3_108_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul3_108_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul3_108_port_byte_out_7[2:0])  //o
  );
  Mul2 mul2_109 (
    .port_byte_in_0  (port_state_in_9_3_0[2:0]     ), //i
    .port_byte_in_1  (port_state_in_9_3_1[2:0]     ), //i
    .port_byte_in_2  (port_state_in_9_3_2[2:0]     ), //i
    .port_byte_in_3  (port_state_in_9_3_3[2:0]     ), //i
    .port_byte_in_4  (port_state_in_9_3_4[2:0]     ), //i
    .port_byte_in_5  (port_state_in_9_3_5[2:0]     ), //i
    .port_byte_in_6  (port_state_in_9_3_6[2:0]     ), //i
    .port_byte_in_7  (port_state_in_9_3_7[2:0]     ), //i
    .port_byte_out_0 (mul2_109_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul2_109_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul2_109_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul2_109_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul2_109_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul2_109_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul2_109_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul2_109_port_byte_out_7[2:0])  //o
  );
  Mul3 mul3_109 (
    .port_byte_in_0  (port_state_in_10_3_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_10_3_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_10_3_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_10_3_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_10_3_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_10_3_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_10_3_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_10_3_7[2:0]    ), //i
    .port_byte_out_0 (mul3_109_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul3_109_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul3_109_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul3_109_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul3_109_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul3_109_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul3_109_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul3_109_port_byte_out_7[2:0])  //o
  );
  Mul2 mul2_110 (
    .port_byte_in_0  (port_state_in_10_3_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_10_3_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_10_3_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_10_3_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_10_3_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_10_3_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_10_3_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_10_3_7[2:0]    ), //i
    .port_byte_out_0 (mul2_110_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul2_110_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul2_110_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul2_110_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul2_110_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul2_110_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul2_110_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul2_110_port_byte_out_7[2:0])  //o
  );
  Mul3 mul3_110 (
    .port_byte_in_0  (port_state_in_11_3_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_11_3_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_11_3_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_11_3_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_11_3_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_11_3_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_11_3_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_11_3_7[2:0]    ), //i
    .port_byte_out_0 (mul3_110_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul3_110_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul3_110_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul3_110_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul3_110_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul3_110_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul3_110_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul3_110_port_byte_out_7[2:0])  //o
  );
  Mul2 mul2_111 (
    .port_byte_in_0  (port_state_in_11_3_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_11_3_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_11_3_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_11_3_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_11_3_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_11_3_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_11_3_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_11_3_7[2:0]    ), //i
    .port_byte_out_0 (mul2_111_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul2_111_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul2_111_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul2_111_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul2_111_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul2_111_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul2_111_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul2_111_port_byte_out_7[2:0])  //o
  );
  Mul3 mul3_111 (
    .port_byte_in_0  (port_state_in_8_3_0[2:0]     ), //i
    .port_byte_in_1  (port_state_in_8_3_1[2:0]     ), //i
    .port_byte_in_2  (port_state_in_8_3_2[2:0]     ), //i
    .port_byte_in_3  (port_state_in_8_3_3[2:0]     ), //i
    .port_byte_in_4  (port_state_in_8_3_4[2:0]     ), //i
    .port_byte_in_5  (port_state_in_8_3_5[2:0]     ), //i
    .port_byte_in_6  (port_state_in_8_3_6[2:0]     ), //i
    .port_byte_in_7  (port_state_in_8_3_7[2:0]     ), //i
    .port_byte_out_0 (mul3_111_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul3_111_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul3_111_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul3_111_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul3_111_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul3_111_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul3_111_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul3_111_port_byte_out_7[2:0])  //o
  );
  Mul2 mul2_112 (
    .port_byte_in_0  (port_state_in_12_0_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_12_0_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_12_0_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_12_0_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_12_0_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_12_0_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_12_0_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_12_0_7[2:0]    ), //i
    .port_byte_out_0 (mul2_112_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul2_112_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul2_112_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul2_112_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul2_112_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul2_112_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul2_112_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul2_112_port_byte_out_7[2:0])  //o
  );
  Mul3 mul3_112 (
    .port_byte_in_0  (port_state_in_13_0_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_13_0_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_13_0_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_13_0_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_13_0_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_13_0_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_13_0_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_13_0_7[2:0]    ), //i
    .port_byte_out_0 (mul3_112_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul3_112_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul3_112_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul3_112_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul3_112_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul3_112_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul3_112_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul3_112_port_byte_out_7[2:0])  //o
  );
  Mul2 mul2_113 (
    .port_byte_in_0  (port_state_in_13_0_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_13_0_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_13_0_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_13_0_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_13_0_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_13_0_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_13_0_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_13_0_7[2:0]    ), //i
    .port_byte_out_0 (mul2_113_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul2_113_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul2_113_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul2_113_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul2_113_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul2_113_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul2_113_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul2_113_port_byte_out_7[2:0])  //o
  );
  Mul3 mul3_113 (
    .port_byte_in_0  (port_state_in_14_0_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_14_0_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_14_0_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_14_0_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_14_0_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_14_0_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_14_0_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_14_0_7[2:0]    ), //i
    .port_byte_out_0 (mul3_113_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul3_113_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul3_113_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul3_113_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul3_113_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul3_113_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul3_113_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul3_113_port_byte_out_7[2:0])  //o
  );
  Mul2 mul2_114 (
    .port_byte_in_0  (port_state_in_14_0_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_14_0_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_14_0_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_14_0_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_14_0_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_14_0_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_14_0_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_14_0_7[2:0]    ), //i
    .port_byte_out_0 (mul2_114_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul2_114_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul2_114_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul2_114_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul2_114_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul2_114_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul2_114_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul2_114_port_byte_out_7[2:0])  //o
  );
  Mul3 mul3_114 (
    .port_byte_in_0  (port_state_in_15_0_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_15_0_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_15_0_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_15_0_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_15_0_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_15_0_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_15_0_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_15_0_7[2:0]    ), //i
    .port_byte_out_0 (mul3_114_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul3_114_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul3_114_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul3_114_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul3_114_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul3_114_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul3_114_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul3_114_port_byte_out_7[2:0])  //o
  );
  Mul2 mul2_115 (
    .port_byte_in_0  (port_state_in_15_0_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_15_0_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_15_0_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_15_0_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_15_0_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_15_0_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_15_0_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_15_0_7[2:0]    ), //i
    .port_byte_out_0 (mul2_115_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul2_115_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul2_115_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul2_115_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul2_115_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul2_115_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul2_115_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul2_115_port_byte_out_7[2:0])  //o
  );
  Mul3 mul3_115 (
    .port_byte_in_0  (port_state_in_12_0_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_12_0_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_12_0_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_12_0_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_12_0_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_12_0_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_12_0_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_12_0_7[2:0]    ), //i
    .port_byte_out_0 (mul3_115_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul3_115_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul3_115_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul3_115_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul3_115_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul3_115_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul3_115_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul3_115_port_byte_out_7[2:0])  //o
  );
  Mul2 mul2_116 (
    .port_byte_in_0  (port_state_in_12_1_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_12_1_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_12_1_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_12_1_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_12_1_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_12_1_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_12_1_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_12_1_7[2:0]    ), //i
    .port_byte_out_0 (mul2_116_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul2_116_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul2_116_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul2_116_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul2_116_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul2_116_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul2_116_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul2_116_port_byte_out_7[2:0])  //o
  );
  Mul3 mul3_116 (
    .port_byte_in_0  (port_state_in_13_1_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_13_1_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_13_1_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_13_1_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_13_1_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_13_1_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_13_1_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_13_1_7[2:0]    ), //i
    .port_byte_out_0 (mul3_116_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul3_116_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul3_116_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul3_116_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul3_116_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul3_116_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul3_116_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul3_116_port_byte_out_7[2:0])  //o
  );
  Mul2 mul2_117 (
    .port_byte_in_0  (port_state_in_13_1_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_13_1_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_13_1_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_13_1_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_13_1_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_13_1_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_13_1_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_13_1_7[2:0]    ), //i
    .port_byte_out_0 (mul2_117_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul2_117_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul2_117_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul2_117_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul2_117_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul2_117_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul2_117_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul2_117_port_byte_out_7[2:0])  //o
  );
  Mul3 mul3_117 (
    .port_byte_in_0  (port_state_in_14_1_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_14_1_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_14_1_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_14_1_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_14_1_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_14_1_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_14_1_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_14_1_7[2:0]    ), //i
    .port_byte_out_0 (mul3_117_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul3_117_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul3_117_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul3_117_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul3_117_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul3_117_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul3_117_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul3_117_port_byte_out_7[2:0])  //o
  );
  Mul2 mul2_118 (
    .port_byte_in_0  (port_state_in_14_1_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_14_1_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_14_1_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_14_1_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_14_1_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_14_1_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_14_1_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_14_1_7[2:0]    ), //i
    .port_byte_out_0 (mul2_118_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul2_118_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul2_118_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul2_118_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul2_118_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul2_118_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul2_118_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul2_118_port_byte_out_7[2:0])  //o
  );
  Mul3 mul3_118 (
    .port_byte_in_0  (port_state_in_15_1_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_15_1_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_15_1_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_15_1_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_15_1_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_15_1_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_15_1_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_15_1_7[2:0]    ), //i
    .port_byte_out_0 (mul3_118_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul3_118_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul3_118_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul3_118_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul3_118_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul3_118_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul3_118_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul3_118_port_byte_out_7[2:0])  //o
  );
  Mul2 mul2_119 (
    .port_byte_in_0  (port_state_in_15_1_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_15_1_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_15_1_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_15_1_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_15_1_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_15_1_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_15_1_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_15_1_7[2:0]    ), //i
    .port_byte_out_0 (mul2_119_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul2_119_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul2_119_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul2_119_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul2_119_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul2_119_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul2_119_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul2_119_port_byte_out_7[2:0])  //o
  );
  Mul3 mul3_119 (
    .port_byte_in_0  (port_state_in_12_1_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_12_1_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_12_1_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_12_1_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_12_1_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_12_1_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_12_1_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_12_1_7[2:0]    ), //i
    .port_byte_out_0 (mul3_119_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul3_119_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul3_119_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul3_119_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul3_119_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul3_119_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul3_119_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul3_119_port_byte_out_7[2:0])  //o
  );
  Mul2 mul2_120 (
    .port_byte_in_0  (port_state_in_12_2_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_12_2_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_12_2_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_12_2_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_12_2_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_12_2_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_12_2_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_12_2_7[2:0]    ), //i
    .port_byte_out_0 (mul2_120_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul2_120_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul2_120_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul2_120_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul2_120_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul2_120_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul2_120_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul2_120_port_byte_out_7[2:0])  //o
  );
  Mul3 mul3_120 (
    .port_byte_in_0  (port_state_in_13_2_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_13_2_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_13_2_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_13_2_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_13_2_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_13_2_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_13_2_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_13_2_7[2:0]    ), //i
    .port_byte_out_0 (mul3_120_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul3_120_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul3_120_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul3_120_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul3_120_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul3_120_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul3_120_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul3_120_port_byte_out_7[2:0])  //o
  );
  Mul2 mul2_121 (
    .port_byte_in_0  (port_state_in_13_2_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_13_2_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_13_2_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_13_2_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_13_2_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_13_2_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_13_2_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_13_2_7[2:0]    ), //i
    .port_byte_out_0 (mul2_121_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul2_121_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul2_121_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul2_121_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul2_121_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul2_121_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul2_121_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul2_121_port_byte_out_7[2:0])  //o
  );
  Mul3 mul3_121 (
    .port_byte_in_0  (port_state_in_14_2_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_14_2_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_14_2_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_14_2_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_14_2_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_14_2_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_14_2_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_14_2_7[2:0]    ), //i
    .port_byte_out_0 (mul3_121_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul3_121_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul3_121_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul3_121_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul3_121_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul3_121_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul3_121_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul3_121_port_byte_out_7[2:0])  //o
  );
  Mul2 mul2_122 (
    .port_byte_in_0  (port_state_in_14_2_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_14_2_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_14_2_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_14_2_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_14_2_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_14_2_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_14_2_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_14_2_7[2:0]    ), //i
    .port_byte_out_0 (mul2_122_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul2_122_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul2_122_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul2_122_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul2_122_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul2_122_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul2_122_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul2_122_port_byte_out_7[2:0])  //o
  );
  Mul3 mul3_122 (
    .port_byte_in_0  (port_state_in_15_2_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_15_2_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_15_2_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_15_2_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_15_2_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_15_2_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_15_2_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_15_2_7[2:0]    ), //i
    .port_byte_out_0 (mul3_122_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul3_122_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul3_122_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul3_122_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul3_122_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul3_122_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul3_122_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul3_122_port_byte_out_7[2:0])  //o
  );
  Mul2 mul2_123 (
    .port_byte_in_0  (port_state_in_15_2_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_15_2_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_15_2_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_15_2_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_15_2_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_15_2_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_15_2_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_15_2_7[2:0]    ), //i
    .port_byte_out_0 (mul2_123_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul2_123_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul2_123_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul2_123_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul2_123_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul2_123_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul2_123_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul2_123_port_byte_out_7[2:0])  //o
  );
  Mul3 mul3_123 (
    .port_byte_in_0  (port_state_in_12_2_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_12_2_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_12_2_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_12_2_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_12_2_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_12_2_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_12_2_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_12_2_7[2:0]    ), //i
    .port_byte_out_0 (mul3_123_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul3_123_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul3_123_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul3_123_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul3_123_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul3_123_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul3_123_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul3_123_port_byte_out_7[2:0])  //o
  );
  Mul2 mul2_124 (
    .port_byte_in_0  (port_state_in_12_3_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_12_3_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_12_3_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_12_3_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_12_3_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_12_3_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_12_3_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_12_3_7[2:0]    ), //i
    .port_byte_out_0 (mul2_124_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul2_124_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul2_124_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul2_124_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul2_124_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul2_124_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul2_124_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul2_124_port_byte_out_7[2:0])  //o
  );
  Mul3 mul3_124 (
    .port_byte_in_0  (port_state_in_13_3_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_13_3_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_13_3_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_13_3_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_13_3_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_13_3_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_13_3_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_13_3_7[2:0]    ), //i
    .port_byte_out_0 (mul3_124_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul3_124_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul3_124_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul3_124_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul3_124_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul3_124_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul3_124_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul3_124_port_byte_out_7[2:0])  //o
  );
  Mul2 mul2_125 (
    .port_byte_in_0  (port_state_in_13_3_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_13_3_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_13_3_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_13_3_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_13_3_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_13_3_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_13_3_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_13_3_7[2:0]    ), //i
    .port_byte_out_0 (mul2_125_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul2_125_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul2_125_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul2_125_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul2_125_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul2_125_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul2_125_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul2_125_port_byte_out_7[2:0])  //o
  );
  Mul3 mul3_125 (
    .port_byte_in_0  (port_state_in_14_3_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_14_3_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_14_3_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_14_3_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_14_3_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_14_3_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_14_3_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_14_3_7[2:0]    ), //i
    .port_byte_out_0 (mul3_125_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul3_125_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul3_125_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul3_125_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul3_125_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul3_125_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul3_125_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul3_125_port_byte_out_7[2:0])  //o
  );
  Mul2 mul2_126 (
    .port_byte_in_0  (port_state_in_14_3_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_14_3_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_14_3_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_14_3_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_14_3_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_14_3_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_14_3_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_14_3_7[2:0]    ), //i
    .port_byte_out_0 (mul2_126_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul2_126_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul2_126_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul2_126_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul2_126_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul2_126_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul2_126_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul2_126_port_byte_out_7[2:0])  //o
  );
  Mul3 mul3_126 (
    .port_byte_in_0  (port_state_in_15_3_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_15_3_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_15_3_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_15_3_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_15_3_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_15_3_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_15_3_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_15_3_7[2:0]    ), //i
    .port_byte_out_0 (mul3_126_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul3_126_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul3_126_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul3_126_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul3_126_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul3_126_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul3_126_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul3_126_port_byte_out_7[2:0])  //o
  );
  Mul2 mul2_127 (
    .port_byte_in_0  (port_state_in_15_3_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_15_3_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_15_3_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_15_3_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_15_3_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_15_3_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_15_3_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_15_3_7[2:0]    ), //i
    .port_byte_out_0 (mul2_127_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul2_127_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul2_127_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul2_127_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul2_127_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul2_127_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul2_127_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul2_127_port_byte_out_7[2:0])  //o
  );
  Mul3 mul3_127 (
    .port_byte_in_0  (port_state_in_12_3_0[2:0]    ), //i
    .port_byte_in_1  (port_state_in_12_3_1[2:0]    ), //i
    .port_byte_in_2  (port_state_in_12_3_2[2:0]    ), //i
    .port_byte_in_3  (port_state_in_12_3_3[2:0]    ), //i
    .port_byte_in_4  (port_state_in_12_3_4[2:0]    ), //i
    .port_byte_in_5  (port_state_in_12_3_5[2:0]    ), //i
    .port_byte_in_6  (port_state_in_12_3_6[2:0]    ), //i
    .port_byte_in_7  (port_state_in_12_3_7[2:0]    ), //i
    .port_byte_out_0 (mul3_127_port_byte_out_0[2:0]), //o
    .port_byte_out_1 (mul3_127_port_byte_out_1[2:0]), //o
    .port_byte_out_2 (mul3_127_port_byte_out_2[2:0]), //o
    .port_byte_out_3 (mul3_127_port_byte_out_3[2:0]), //o
    .port_byte_out_4 (mul3_127_port_byte_out_4[2:0]), //o
    .port_byte_out_5 (mul3_127_port_byte_out_5[2:0]), //o
    .port_byte_out_6 (mul3_127_port_byte_out_6[2:0]), //o
    .port_byte_out_7 (mul3_127_port_byte_out_7[2:0])  //o
  );
  assign state_out_0_0_0 = (((mul2_64_port_byte_out_0 ^ mul3_64_port_byte_out_0) ^ port_state_in_2_0_0) ^ port_state_in_3_0_0);
  assign state_out_1_0_0 = (((mul2_65_port_byte_out_0 ^ mul3_65_port_byte_out_0) ^ port_state_in_0_0_0) ^ port_state_in_3_0_0);
  assign state_out_2_0_0 = (((mul2_66_port_byte_out_0 ^ mul3_66_port_byte_out_0) ^ port_state_in_0_0_0) ^ port_state_in_1_0_0);
  assign state_out_3_0_0 = (((mul2_67_port_byte_out_0 ^ mul3_67_port_byte_out_0) ^ port_state_in_1_0_0) ^ port_state_in_2_0_0);
  assign state_out_0_0_1 = (((mul2_64_port_byte_out_1 ^ mul3_64_port_byte_out_1) ^ port_state_in_2_0_1) ^ port_state_in_3_0_1);
  assign state_out_1_0_1 = (((mul2_65_port_byte_out_1 ^ mul3_65_port_byte_out_1) ^ port_state_in_0_0_1) ^ port_state_in_3_0_1);
  assign state_out_2_0_1 = (((mul2_66_port_byte_out_1 ^ mul3_66_port_byte_out_1) ^ port_state_in_0_0_1) ^ port_state_in_1_0_1);
  assign state_out_3_0_1 = (((mul2_67_port_byte_out_1 ^ mul3_67_port_byte_out_1) ^ port_state_in_1_0_1) ^ port_state_in_2_0_1);
  assign state_out_0_0_2 = (((mul2_64_port_byte_out_2 ^ mul3_64_port_byte_out_2) ^ port_state_in_2_0_2) ^ port_state_in_3_0_2);
  assign state_out_1_0_2 = (((mul2_65_port_byte_out_2 ^ mul3_65_port_byte_out_2) ^ port_state_in_0_0_2) ^ port_state_in_3_0_2);
  assign state_out_2_0_2 = (((mul2_66_port_byte_out_2 ^ mul3_66_port_byte_out_2) ^ port_state_in_0_0_2) ^ port_state_in_1_0_2);
  assign state_out_3_0_2 = (((mul2_67_port_byte_out_2 ^ mul3_67_port_byte_out_2) ^ port_state_in_1_0_2) ^ port_state_in_2_0_2);
  assign state_out_0_0_3 = (((mul2_64_port_byte_out_3 ^ mul3_64_port_byte_out_3) ^ port_state_in_2_0_3) ^ port_state_in_3_0_3);
  assign state_out_1_0_3 = (((mul2_65_port_byte_out_3 ^ mul3_65_port_byte_out_3) ^ port_state_in_0_0_3) ^ port_state_in_3_0_3);
  assign state_out_2_0_3 = (((mul2_66_port_byte_out_3 ^ mul3_66_port_byte_out_3) ^ port_state_in_0_0_3) ^ port_state_in_1_0_3);
  assign state_out_3_0_3 = (((mul2_67_port_byte_out_3 ^ mul3_67_port_byte_out_3) ^ port_state_in_1_0_3) ^ port_state_in_2_0_3);
  assign state_out_0_0_4 = (((mul2_64_port_byte_out_4 ^ mul3_64_port_byte_out_4) ^ port_state_in_2_0_4) ^ port_state_in_3_0_4);
  assign state_out_1_0_4 = (((mul2_65_port_byte_out_4 ^ mul3_65_port_byte_out_4) ^ port_state_in_0_0_4) ^ port_state_in_3_0_4);
  assign state_out_2_0_4 = (((mul2_66_port_byte_out_4 ^ mul3_66_port_byte_out_4) ^ port_state_in_0_0_4) ^ port_state_in_1_0_4);
  assign state_out_3_0_4 = (((mul2_67_port_byte_out_4 ^ mul3_67_port_byte_out_4) ^ port_state_in_1_0_4) ^ port_state_in_2_0_4);
  assign state_out_0_0_5 = (((mul2_64_port_byte_out_5 ^ mul3_64_port_byte_out_5) ^ port_state_in_2_0_5) ^ port_state_in_3_0_5);
  assign state_out_1_0_5 = (((mul2_65_port_byte_out_5 ^ mul3_65_port_byte_out_5) ^ port_state_in_0_0_5) ^ port_state_in_3_0_5);
  assign state_out_2_0_5 = (((mul2_66_port_byte_out_5 ^ mul3_66_port_byte_out_5) ^ port_state_in_0_0_5) ^ port_state_in_1_0_5);
  assign state_out_3_0_5 = (((mul2_67_port_byte_out_5 ^ mul3_67_port_byte_out_5) ^ port_state_in_1_0_5) ^ port_state_in_2_0_5);
  assign state_out_0_0_6 = (((mul2_64_port_byte_out_6 ^ mul3_64_port_byte_out_6) ^ port_state_in_2_0_6) ^ port_state_in_3_0_6);
  assign state_out_1_0_6 = (((mul2_65_port_byte_out_6 ^ mul3_65_port_byte_out_6) ^ port_state_in_0_0_6) ^ port_state_in_3_0_6);
  assign state_out_2_0_6 = (((mul2_66_port_byte_out_6 ^ mul3_66_port_byte_out_6) ^ port_state_in_0_0_6) ^ port_state_in_1_0_6);
  assign state_out_3_0_6 = (((mul2_67_port_byte_out_6 ^ mul3_67_port_byte_out_6) ^ port_state_in_1_0_6) ^ port_state_in_2_0_6);
  assign state_out_0_0_7 = (((mul2_64_port_byte_out_7 ^ mul3_64_port_byte_out_7) ^ port_state_in_2_0_7) ^ port_state_in_3_0_7);
  assign state_out_1_0_7 = (((mul2_65_port_byte_out_7 ^ mul3_65_port_byte_out_7) ^ port_state_in_0_0_7) ^ port_state_in_3_0_7);
  assign state_out_2_0_7 = (((mul2_66_port_byte_out_7 ^ mul3_66_port_byte_out_7) ^ port_state_in_0_0_7) ^ port_state_in_1_0_7);
  assign state_out_3_0_7 = (((mul2_67_port_byte_out_7 ^ mul3_67_port_byte_out_7) ^ port_state_in_1_0_7) ^ port_state_in_2_0_7);
  assign state_out_0_1_0 = (((mul2_68_port_byte_out_0 ^ mul3_68_port_byte_out_0) ^ port_state_in_2_1_0) ^ port_state_in_3_1_0);
  assign state_out_1_1_0 = (((mul2_69_port_byte_out_0 ^ mul3_69_port_byte_out_0) ^ port_state_in_0_1_0) ^ port_state_in_3_1_0);
  assign state_out_2_1_0 = (((mul2_70_port_byte_out_0 ^ mul3_70_port_byte_out_0) ^ port_state_in_0_1_0) ^ port_state_in_1_1_0);
  assign state_out_3_1_0 = (((mul2_71_port_byte_out_0 ^ mul3_71_port_byte_out_0) ^ port_state_in_1_1_0) ^ port_state_in_2_1_0);
  assign state_out_0_1_1 = (((mul2_68_port_byte_out_1 ^ mul3_68_port_byte_out_1) ^ port_state_in_2_1_1) ^ port_state_in_3_1_1);
  assign state_out_1_1_1 = (((mul2_69_port_byte_out_1 ^ mul3_69_port_byte_out_1) ^ port_state_in_0_1_1) ^ port_state_in_3_1_1);
  assign state_out_2_1_1 = (((mul2_70_port_byte_out_1 ^ mul3_70_port_byte_out_1) ^ port_state_in_0_1_1) ^ port_state_in_1_1_1);
  assign state_out_3_1_1 = (((mul2_71_port_byte_out_1 ^ mul3_71_port_byte_out_1) ^ port_state_in_1_1_1) ^ port_state_in_2_1_1);
  assign state_out_0_1_2 = (((mul2_68_port_byte_out_2 ^ mul3_68_port_byte_out_2) ^ port_state_in_2_1_2) ^ port_state_in_3_1_2);
  assign state_out_1_1_2 = (((mul2_69_port_byte_out_2 ^ mul3_69_port_byte_out_2) ^ port_state_in_0_1_2) ^ port_state_in_3_1_2);
  assign state_out_2_1_2 = (((mul2_70_port_byte_out_2 ^ mul3_70_port_byte_out_2) ^ port_state_in_0_1_2) ^ port_state_in_1_1_2);
  assign state_out_3_1_2 = (((mul2_71_port_byte_out_2 ^ mul3_71_port_byte_out_2) ^ port_state_in_1_1_2) ^ port_state_in_2_1_2);
  assign state_out_0_1_3 = (((mul2_68_port_byte_out_3 ^ mul3_68_port_byte_out_3) ^ port_state_in_2_1_3) ^ port_state_in_3_1_3);
  assign state_out_1_1_3 = (((mul2_69_port_byte_out_3 ^ mul3_69_port_byte_out_3) ^ port_state_in_0_1_3) ^ port_state_in_3_1_3);
  assign state_out_2_1_3 = (((mul2_70_port_byte_out_3 ^ mul3_70_port_byte_out_3) ^ port_state_in_0_1_3) ^ port_state_in_1_1_3);
  assign state_out_3_1_3 = (((mul2_71_port_byte_out_3 ^ mul3_71_port_byte_out_3) ^ port_state_in_1_1_3) ^ port_state_in_2_1_3);
  assign state_out_0_1_4 = (((mul2_68_port_byte_out_4 ^ mul3_68_port_byte_out_4) ^ port_state_in_2_1_4) ^ port_state_in_3_1_4);
  assign state_out_1_1_4 = (((mul2_69_port_byte_out_4 ^ mul3_69_port_byte_out_4) ^ port_state_in_0_1_4) ^ port_state_in_3_1_4);
  assign state_out_2_1_4 = (((mul2_70_port_byte_out_4 ^ mul3_70_port_byte_out_4) ^ port_state_in_0_1_4) ^ port_state_in_1_1_4);
  assign state_out_3_1_4 = (((mul2_71_port_byte_out_4 ^ mul3_71_port_byte_out_4) ^ port_state_in_1_1_4) ^ port_state_in_2_1_4);
  assign state_out_0_1_5 = (((mul2_68_port_byte_out_5 ^ mul3_68_port_byte_out_5) ^ port_state_in_2_1_5) ^ port_state_in_3_1_5);
  assign state_out_1_1_5 = (((mul2_69_port_byte_out_5 ^ mul3_69_port_byte_out_5) ^ port_state_in_0_1_5) ^ port_state_in_3_1_5);
  assign state_out_2_1_5 = (((mul2_70_port_byte_out_5 ^ mul3_70_port_byte_out_5) ^ port_state_in_0_1_5) ^ port_state_in_1_1_5);
  assign state_out_3_1_5 = (((mul2_71_port_byte_out_5 ^ mul3_71_port_byte_out_5) ^ port_state_in_1_1_5) ^ port_state_in_2_1_5);
  assign state_out_0_1_6 = (((mul2_68_port_byte_out_6 ^ mul3_68_port_byte_out_6) ^ port_state_in_2_1_6) ^ port_state_in_3_1_6);
  assign state_out_1_1_6 = (((mul2_69_port_byte_out_6 ^ mul3_69_port_byte_out_6) ^ port_state_in_0_1_6) ^ port_state_in_3_1_6);
  assign state_out_2_1_6 = (((mul2_70_port_byte_out_6 ^ mul3_70_port_byte_out_6) ^ port_state_in_0_1_6) ^ port_state_in_1_1_6);
  assign state_out_3_1_6 = (((mul2_71_port_byte_out_6 ^ mul3_71_port_byte_out_6) ^ port_state_in_1_1_6) ^ port_state_in_2_1_6);
  assign state_out_0_1_7 = (((mul2_68_port_byte_out_7 ^ mul3_68_port_byte_out_7) ^ port_state_in_2_1_7) ^ port_state_in_3_1_7);
  assign state_out_1_1_7 = (((mul2_69_port_byte_out_7 ^ mul3_69_port_byte_out_7) ^ port_state_in_0_1_7) ^ port_state_in_3_1_7);
  assign state_out_2_1_7 = (((mul2_70_port_byte_out_7 ^ mul3_70_port_byte_out_7) ^ port_state_in_0_1_7) ^ port_state_in_1_1_7);
  assign state_out_3_1_7 = (((mul2_71_port_byte_out_7 ^ mul3_71_port_byte_out_7) ^ port_state_in_1_1_7) ^ port_state_in_2_1_7);
  assign state_out_0_2_0 = (((mul2_72_port_byte_out_0 ^ mul3_72_port_byte_out_0) ^ port_state_in_2_2_0) ^ port_state_in_3_2_0);
  assign state_out_1_2_0 = (((mul2_73_port_byte_out_0 ^ mul3_73_port_byte_out_0) ^ port_state_in_0_2_0) ^ port_state_in_3_2_0);
  assign state_out_2_2_0 = (((mul2_74_port_byte_out_0 ^ mul3_74_port_byte_out_0) ^ port_state_in_0_2_0) ^ port_state_in_1_2_0);
  assign state_out_3_2_0 = (((mul2_75_port_byte_out_0 ^ mul3_75_port_byte_out_0) ^ port_state_in_1_2_0) ^ port_state_in_2_2_0);
  assign state_out_0_2_1 = (((mul2_72_port_byte_out_1 ^ mul3_72_port_byte_out_1) ^ port_state_in_2_2_1) ^ port_state_in_3_2_1);
  assign state_out_1_2_1 = (((mul2_73_port_byte_out_1 ^ mul3_73_port_byte_out_1) ^ port_state_in_0_2_1) ^ port_state_in_3_2_1);
  assign state_out_2_2_1 = (((mul2_74_port_byte_out_1 ^ mul3_74_port_byte_out_1) ^ port_state_in_0_2_1) ^ port_state_in_1_2_1);
  assign state_out_3_2_1 = (((mul2_75_port_byte_out_1 ^ mul3_75_port_byte_out_1) ^ port_state_in_1_2_1) ^ port_state_in_2_2_1);
  assign state_out_0_2_2 = (((mul2_72_port_byte_out_2 ^ mul3_72_port_byte_out_2) ^ port_state_in_2_2_2) ^ port_state_in_3_2_2);
  assign state_out_1_2_2 = (((mul2_73_port_byte_out_2 ^ mul3_73_port_byte_out_2) ^ port_state_in_0_2_2) ^ port_state_in_3_2_2);
  assign state_out_2_2_2 = (((mul2_74_port_byte_out_2 ^ mul3_74_port_byte_out_2) ^ port_state_in_0_2_2) ^ port_state_in_1_2_2);
  assign state_out_3_2_2 = (((mul2_75_port_byte_out_2 ^ mul3_75_port_byte_out_2) ^ port_state_in_1_2_2) ^ port_state_in_2_2_2);
  assign state_out_0_2_3 = (((mul2_72_port_byte_out_3 ^ mul3_72_port_byte_out_3) ^ port_state_in_2_2_3) ^ port_state_in_3_2_3);
  assign state_out_1_2_3 = (((mul2_73_port_byte_out_3 ^ mul3_73_port_byte_out_3) ^ port_state_in_0_2_3) ^ port_state_in_3_2_3);
  assign state_out_2_2_3 = (((mul2_74_port_byte_out_3 ^ mul3_74_port_byte_out_3) ^ port_state_in_0_2_3) ^ port_state_in_1_2_3);
  assign state_out_3_2_3 = (((mul2_75_port_byte_out_3 ^ mul3_75_port_byte_out_3) ^ port_state_in_1_2_3) ^ port_state_in_2_2_3);
  assign state_out_0_2_4 = (((mul2_72_port_byte_out_4 ^ mul3_72_port_byte_out_4) ^ port_state_in_2_2_4) ^ port_state_in_3_2_4);
  assign state_out_1_2_4 = (((mul2_73_port_byte_out_4 ^ mul3_73_port_byte_out_4) ^ port_state_in_0_2_4) ^ port_state_in_3_2_4);
  assign state_out_2_2_4 = (((mul2_74_port_byte_out_4 ^ mul3_74_port_byte_out_4) ^ port_state_in_0_2_4) ^ port_state_in_1_2_4);
  assign state_out_3_2_4 = (((mul2_75_port_byte_out_4 ^ mul3_75_port_byte_out_4) ^ port_state_in_1_2_4) ^ port_state_in_2_2_4);
  assign state_out_0_2_5 = (((mul2_72_port_byte_out_5 ^ mul3_72_port_byte_out_5) ^ port_state_in_2_2_5) ^ port_state_in_3_2_5);
  assign state_out_1_2_5 = (((mul2_73_port_byte_out_5 ^ mul3_73_port_byte_out_5) ^ port_state_in_0_2_5) ^ port_state_in_3_2_5);
  assign state_out_2_2_5 = (((mul2_74_port_byte_out_5 ^ mul3_74_port_byte_out_5) ^ port_state_in_0_2_5) ^ port_state_in_1_2_5);
  assign state_out_3_2_5 = (((mul2_75_port_byte_out_5 ^ mul3_75_port_byte_out_5) ^ port_state_in_1_2_5) ^ port_state_in_2_2_5);
  assign state_out_0_2_6 = (((mul2_72_port_byte_out_6 ^ mul3_72_port_byte_out_6) ^ port_state_in_2_2_6) ^ port_state_in_3_2_6);
  assign state_out_1_2_6 = (((mul2_73_port_byte_out_6 ^ mul3_73_port_byte_out_6) ^ port_state_in_0_2_6) ^ port_state_in_3_2_6);
  assign state_out_2_2_6 = (((mul2_74_port_byte_out_6 ^ mul3_74_port_byte_out_6) ^ port_state_in_0_2_6) ^ port_state_in_1_2_6);
  assign state_out_3_2_6 = (((mul2_75_port_byte_out_6 ^ mul3_75_port_byte_out_6) ^ port_state_in_1_2_6) ^ port_state_in_2_2_6);
  assign state_out_0_2_7 = (((mul2_72_port_byte_out_7 ^ mul3_72_port_byte_out_7) ^ port_state_in_2_2_7) ^ port_state_in_3_2_7);
  assign state_out_1_2_7 = (((mul2_73_port_byte_out_7 ^ mul3_73_port_byte_out_7) ^ port_state_in_0_2_7) ^ port_state_in_3_2_7);
  assign state_out_2_2_7 = (((mul2_74_port_byte_out_7 ^ mul3_74_port_byte_out_7) ^ port_state_in_0_2_7) ^ port_state_in_1_2_7);
  assign state_out_3_2_7 = (((mul2_75_port_byte_out_7 ^ mul3_75_port_byte_out_7) ^ port_state_in_1_2_7) ^ port_state_in_2_2_7);
  assign state_out_0_3_0 = (((mul2_76_port_byte_out_0 ^ mul3_76_port_byte_out_0) ^ port_state_in_2_3_0) ^ port_state_in_3_3_0);
  assign state_out_1_3_0 = (((mul2_77_port_byte_out_0 ^ mul3_77_port_byte_out_0) ^ port_state_in_0_3_0) ^ port_state_in_3_3_0);
  assign state_out_2_3_0 = (((mul2_78_port_byte_out_0 ^ mul3_78_port_byte_out_0) ^ port_state_in_0_3_0) ^ port_state_in_1_3_0);
  assign state_out_3_3_0 = (((mul2_79_port_byte_out_0 ^ mul3_79_port_byte_out_0) ^ port_state_in_1_3_0) ^ port_state_in_2_3_0);
  assign state_out_0_3_1 = (((mul2_76_port_byte_out_1 ^ mul3_76_port_byte_out_1) ^ port_state_in_2_3_1) ^ port_state_in_3_3_1);
  assign state_out_1_3_1 = (((mul2_77_port_byte_out_1 ^ mul3_77_port_byte_out_1) ^ port_state_in_0_3_1) ^ port_state_in_3_3_1);
  assign state_out_2_3_1 = (((mul2_78_port_byte_out_1 ^ mul3_78_port_byte_out_1) ^ port_state_in_0_3_1) ^ port_state_in_1_3_1);
  assign state_out_3_3_1 = (((mul2_79_port_byte_out_1 ^ mul3_79_port_byte_out_1) ^ port_state_in_1_3_1) ^ port_state_in_2_3_1);
  assign state_out_0_3_2 = (((mul2_76_port_byte_out_2 ^ mul3_76_port_byte_out_2) ^ port_state_in_2_3_2) ^ port_state_in_3_3_2);
  assign state_out_1_3_2 = (((mul2_77_port_byte_out_2 ^ mul3_77_port_byte_out_2) ^ port_state_in_0_3_2) ^ port_state_in_3_3_2);
  assign state_out_2_3_2 = (((mul2_78_port_byte_out_2 ^ mul3_78_port_byte_out_2) ^ port_state_in_0_3_2) ^ port_state_in_1_3_2);
  assign state_out_3_3_2 = (((mul2_79_port_byte_out_2 ^ mul3_79_port_byte_out_2) ^ port_state_in_1_3_2) ^ port_state_in_2_3_2);
  assign state_out_0_3_3 = (((mul2_76_port_byte_out_3 ^ mul3_76_port_byte_out_3) ^ port_state_in_2_3_3) ^ port_state_in_3_3_3);
  assign state_out_1_3_3 = (((mul2_77_port_byte_out_3 ^ mul3_77_port_byte_out_3) ^ port_state_in_0_3_3) ^ port_state_in_3_3_3);
  assign state_out_2_3_3 = (((mul2_78_port_byte_out_3 ^ mul3_78_port_byte_out_3) ^ port_state_in_0_3_3) ^ port_state_in_1_3_3);
  assign state_out_3_3_3 = (((mul2_79_port_byte_out_3 ^ mul3_79_port_byte_out_3) ^ port_state_in_1_3_3) ^ port_state_in_2_3_3);
  assign state_out_0_3_4 = (((mul2_76_port_byte_out_4 ^ mul3_76_port_byte_out_4) ^ port_state_in_2_3_4) ^ port_state_in_3_3_4);
  assign state_out_1_3_4 = (((mul2_77_port_byte_out_4 ^ mul3_77_port_byte_out_4) ^ port_state_in_0_3_4) ^ port_state_in_3_3_4);
  assign state_out_2_3_4 = (((mul2_78_port_byte_out_4 ^ mul3_78_port_byte_out_4) ^ port_state_in_0_3_4) ^ port_state_in_1_3_4);
  assign state_out_3_3_4 = (((mul2_79_port_byte_out_4 ^ mul3_79_port_byte_out_4) ^ port_state_in_1_3_4) ^ port_state_in_2_3_4);
  assign state_out_0_3_5 = (((mul2_76_port_byte_out_5 ^ mul3_76_port_byte_out_5) ^ port_state_in_2_3_5) ^ port_state_in_3_3_5);
  assign state_out_1_3_5 = (((mul2_77_port_byte_out_5 ^ mul3_77_port_byte_out_5) ^ port_state_in_0_3_5) ^ port_state_in_3_3_5);
  assign state_out_2_3_5 = (((mul2_78_port_byte_out_5 ^ mul3_78_port_byte_out_5) ^ port_state_in_0_3_5) ^ port_state_in_1_3_5);
  assign state_out_3_3_5 = (((mul2_79_port_byte_out_5 ^ mul3_79_port_byte_out_5) ^ port_state_in_1_3_5) ^ port_state_in_2_3_5);
  assign state_out_0_3_6 = (((mul2_76_port_byte_out_6 ^ mul3_76_port_byte_out_6) ^ port_state_in_2_3_6) ^ port_state_in_3_3_6);
  assign state_out_1_3_6 = (((mul2_77_port_byte_out_6 ^ mul3_77_port_byte_out_6) ^ port_state_in_0_3_6) ^ port_state_in_3_3_6);
  assign state_out_2_3_6 = (((mul2_78_port_byte_out_6 ^ mul3_78_port_byte_out_6) ^ port_state_in_0_3_6) ^ port_state_in_1_3_6);
  assign state_out_3_3_6 = (((mul2_79_port_byte_out_6 ^ mul3_79_port_byte_out_6) ^ port_state_in_1_3_6) ^ port_state_in_2_3_6);
  assign state_out_0_3_7 = (((mul2_76_port_byte_out_7 ^ mul3_76_port_byte_out_7) ^ port_state_in_2_3_7) ^ port_state_in_3_3_7);
  assign state_out_1_3_7 = (((mul2_77_port_byte_out_7 ^ mul3_77_port_byte_out_7) ^ port_state_in_0_3_7) ^ port_state_in_3_3_7);
  assign state_out_2_3_7 = (((mul2_78_port_byte_out_7 ^ mul3_78_port_byte_out_7) ^ port_state_in_0_3_7) ^ port_state_in_1_3_7);
  assign state_out_3_3_7 = (((mul2_79_port_byte_out_7 ^ mul3_79_port_byte_out_7) ^ port_state_in_1_3_7) ^ port_state_in_2_3_7);
  assign state_out_4_0_0 = (((mul2_80_port_byte_out_0 ^ mul3_80_port_byte_out_0) ^ port_state_in_6_0_0) ^ port_state_in_7_0_0);
  assign state_out_5_0_0 = (((mul2_81_port_byte_out_0 ^ mul3_81_port_byte_out_0) ^ port_state_in_4_0_0) ^ port_state_in_7_0_0);
  assign state_out_6_0_0 = (((mul2_82_port_byte_out_0 ^ mul3_82_port_byte_out_0) ^ port_state_in_4_0_0) ^ port_state_in_5_0_0);
  assign state_out_7_0_0 = (((mul2_83_port_byte_out_0 ^ mul3_83_port_byte_out_0) ^ port_state_in_5_0_0) ^ port_state_in_6_0_0);
  assign state_out_4_0_1 = (((mul2_80_port_byte_out_1 ^ mul3_80_port_byte_out_1) ^ port_state_in_6_0_1) ^ port_state_in_7_0_1);
  assign state_out_5_0_1 = (((mul2_81_port_byte_out_1 ^ mul3_81_port_byte_out_1) ^ port_state_in_4_0_1) ^ port_state_in_7_0_1);
  assign state_out_6_0_1 = (((mul2_82_port_byte_out_1 ^ mul3_82_port_byte_out_1) ^ port_state_in_4_0_1) ^ port_state_in_5_0_1);
  assign state_out_7_0_1 = (((mul2_83_port_byte_out_1 ^ mul3_83_port_byte_out_1) ^ port_state_in_5_0_1) ^ port_state_in_6_0_1);
  assign state_out_4_0_2 = (((mul2_80_port_byte_out_2 ^ mul3_80_port_byte_out_2) ^ port_state_in_6_0_2) ^ port_state_in_7_0_2);
  assign state_out_5_0_2 = (((mul2_81_port_byte_out_2 ^ mul3_81_port_byte_out_2) ^ port_state_in_4_0_2) ^ port_state_in_7_0_2);
  assign state_out_6_0_2 = (((mul2_82_port_byte_out_2 ^ mul3_82_port_byte_out_2) ^ port_state_in_4_0_2) ^ port_state_in_5_0_2);
  assign state_out_7_0_2 = (((mul2_83_port_byte_out_2 ^ mul3_83_port_byte_out_2) ^ port_state_in_5_0_2) ^ port_state_in_6_0_2);
  assign state_out_4_0_3 = (((mul2_80_port_byte_out_3 ^ mul3_80_port_byte_out_3) ^ port_state_in_6_0_3) ^ port_state_in_7_0_3);
  assign state_out_5_0_3 = (((mul2_81_port_byte_out_3 ^ mul3_81_port_byte_out_3) ^ port_state_in_4_0_3) ^ port_state_in_7_0_3);
  assign state_out_6_0_3 = (((mul2_82_port_byte_out_3 ^ mul3_82_port_byte_out_3) ^ port_state_in_4_0_3) ^ port_state_in_5_0_3);
  assign state_out_7_0_3 = (((mul2_83_port_byte_out_3 ^ mul3_83_port_byte_out_3) ^ port_state_in_5_0_3) ^ port_state_in_6_0_3);
  assign state_out_4_0_4 = (((mul2_80_port_byte_out_4 ^ mul3_80_port_byte_out_4) ^ port_state_in_6_0_4) ^ port_state_in_7_0_4);
  assign state_out_5_0_4 = (((mul2_81_port_byte_out_4 ^ mul3_81_port_byte_out_4) ^ port_state_in_4_0_4) ^ port_state_in_7_0_4);
  assign state_out_6_0_4 = (((mul2_82_port_byte_out_4 ^ mul3_82_port_byte_out_4) ^ port_state_in_4_0_4) ^ port_state_in_5_0_4);
  assign state_out_7_0_4 = (((mul2_83_port_byte_out_4 ^ mul3_83_port_byte_out_4) ^ port_state_in_5_0_4) ^ port_state_in_6_0_4);
  assign state_out_4_0_5 = (((mul2_80_port_byte_out_5 ^ mul3_80_port_byte_out_5) ^ port_state_in_6_0_5) ^ port_state_in_7_0_5);
  assign state_out_5_0_5 = (((mul2_81_port_byte_out_5 ^ mul3_81_port_byte_out_5) ^ port_state_in_4_0_5) ^ port_state_in_7_0_5);
  assign state_out_6_0_5 = (((mul2_82_port_byte_out_5 ^ mul3_82_port_byte_out_5) ^ port_state_in_4_0_5) ^ port_state_in_5_0_5);
  assign state_out_7_0_5 = (((mul2_83_port_byte_out_5 ^ mul3_83_port_byte_out_5) ^ port_state_in_5_0_5) ^ port_state_in_6_0_5);
  assign state_out_4_0_6 = (((mul2_80_port_byte_out_6 ^ mul3_80_port_byte_out_6) ^ port_state_in_6_0_6) ^ port_state_in_7_0_6);
  assign state_out_5_0_6 = (((mul2_81_port_byte_out_6 ^ mul3_81_port_byte_out_6) ^ port_state_in_4_0_6) ^ port_state_in_7_0_6);
  assign state_out_6_0_6 = (((mul2_82_port_byte_out_6 ^ mul3_82_port_byte_out_6) ^ port_state_in_4_0_6) ^ port_state_in_5_0_6);
  assign state_out_7_0_6 = (((mul2_83_port_byte_out_6 ^ mul3_83_port_byte_out_6) ^ port_state_in_5_0_6) ^ port_state_in_6_0_6);
  assign state_out_4_0_7 = (((mul2_80_port_byte_out_7 ^ mul3_80_port_byte_out_7) ^ port_state_in_6_0_7) ^ port_state_in_7_0_7);
  assign state_out_5_0_7 = (((mul2_81_port_byte_out_7 ^ mul3_81_port_byte_out_7) ^ port_state_in_4_0_7) ^ port_state_in_7_0_7);
  assign state_out_6_0_7 = (((mul2_82_port_byte_out_7 ^ mul3_82_port_byte_out_7) ^ port_state_in_4_0_7) ^ port_state_in_5_0_7);
  assign state_out_7_0_7 = (((mul2_83_port_byte_out_7 ^ mul3_83_port_byte_out_7) ^ port_state_in_5_0_7) ^ port_state_in_6_0_7);
  assign state_out_4_1_0 = (((mul2_84_port_byte_out_0 ^ mul3_84_port_byte_out_0) ^ port_state_in_6_1_0) ^ port_state_in_7_1_0);
  assign state_out_5_1_0 = (((mul2_85_port_byte_out_0 ^ mul3_85_port_byte_out_0) ^ port_state_in_4_1_0) ^ port_state_in_7_1_0);
  assign state_out_6_1_0 = (((mul2_86_port_byte_out_0 ^ mul3_86_port_byte_out_0) ^ port_state_in_4_1_0) ^ port_state_in_5_1_0);
  assign state_out_7_1_0 = (((mul2_87_port_byte_out_0 ^ mul3_87_port_byte_out_0) ^ port_state_in_5_1_0) ^ port_state_in_6_1_0);
  assign state_out_4_1_1 = (((mul2_84_port_byte_out_1 ^ mul3_84_port_byte_out_1) ^ port_state_in_6_1_1) ^ port_state_in_7_1_1);
  assign state_out_5_1_1 = (((mul2_85_port_byte_out_1 ^ mul3_85_port_byte_out_1) ^ port_state_in_4_1_1) ^ port_state_in_7_1_1);
  assign state_out_6_1_1 = (((mul2_86_port_byte_out_1 ^ mul3_86_port_byte_out_1) ^ port_state_in_4_1_1) ^ port_state_in_5_1_1);
  assign state_out_7_1_1 = (((mul2_87_port_byte_out_1 ^ mul3_87_port_byte_out_1) ^ port_state_in_5_1_1) ^ port_state_in_6_1_1);
  assign state_out_4_1_2 = (((mul2_84_port_byte_out_2 ^ mul3_84_port_byte_out_2) ^ port_state_in_6_1_2) ^ port_state_in_7_1_2);
  assign state_out_5_1_2 = (((mul2_85_port_byte_out_2 ^ mul3_85_port_byte_out_2) ^ port_state_in_4_1_2) ^ port_state_in_7_1_2);
  assign state_out_6_1_2 = (((mul2_86_port_byte_out_2 ^ mul3_86_port_byte_out_2) ^ port_state_in_4_1_2) ^ port_state_in_5_1_2);
  assign state_out_7_1_2 = (((mul2_87_port_byte_out_2 ^ mul3_87_port_byte_out_2) ^ port_state_in_5_1_2) ^ port_state_in_6_1_2);
  assign state_out_4_1_3 = (((mul2_84_port_byte_out_3 ^ mul3_84_port_byte_out_3) ^ port_state_in_6_1_3) ^ port_state_in_7_1_3);
  assign state_out_5_1_3 = (((mul2_85_port_byte_out_3 ^ mul3_85_port_byte_out_3) ^ port_state_in_4_1_3) ^ port_state_in_7_1_3);
  assign state_out_6_1_3 = (((mul2_86_port_byte_out_3 ^ mul3_86_port_byte_out_3) ^ port_state_in_4_1_3) ^ port_state_in_5_1_3);
  assign state_out_7_1_3 = (((mul2_87_port_byte_out_3 ^ mul3_87_port_byte_out_3) ^ port_state_in_5_1_3) ^ port_state_in_6_1_3);
  assign state_out_4_1_4 = (((mul2_84_port_byte_out_4 ^ mul3_84_port_byte_out_4) ^ port_state_in_6_1_4) ^ port_state_in_7_1_4);
  assign state_out_5_1_4 = (((mul2_85_port_byte_out_4 ^ mul3_85_port_byte_out_4) ^ port_state_in_4_1_4) ^ port_state_in_7_1_4);
  assign state_out_6_1_4 = (((mul2_86_port_byte_out_4 ^ mul3_86_port_byte_out_4) ^ port_state_in_4_1_4) ^ port_state_in_5_1_4);
  assign state_out_7_1_4 = (((mul2_87_port_byte_out_4 ^ mul3_87_port_byte_out_4) ^ port_state_in_5_1_4) ^ port_state_in_6_1_4);
  assign state_out_4_1_5 = (((mul2_84_port_byte_out_5 ^ mul3_84_port_byte_out_5) ^ port_state_in_6_1_5) ^ port_state_in_7_1_5);
  assign state_out_5_1_5 = (((mul2_85_port_byte_out_5 ^ mul3_85_port_byte_out_5) ^ port_state_in_4_1_5) ^ port_state_in_7_1_5);
  assign state_out_6_1_5 = (((mul2_86_port_byte_out_5 ^ mul3_86_port_byte_out_5) ^ port_state_in_4_1_5) ^ port_state_in_5_1_5);
  assign state_out_7_1_5 = (((mul2_87_port_byte_out_5 ^ mul3_87_port_byte_out_5) ^ port_state_in_5_1_5) ^ port_state_in_6_1_5);
  assign state_out_4_1_6 = (((mul2_84_port_byte_out_6 ^ mul3_84_port_byte_out_6) ^ port_state_in_6_1_6) ^ port_state_in_7_1_6);
  assign state_out_5_1_6 = (((mul2_85_port_byte_out_6 ^ mul3_85_port_byte_out_6) ^ port_state_in_4_1_6) ^ port_state_in_7_1_6);
  assign state_out_6_1_6 = (((mul2_86_port_byte_out_6 ^ mul3_86_port_byte_out_6) ^ port_state_in_4_1_6) ^ port_state_in_5_1_6);
  assign state_out_7_1_6 = (((mul2_87_port_byte_out_6 ^ mul3_87_port_byte_out_6) ^ port_state_in_5_1_6) ^ port_state_in_6_1_6);
  assign state_out_4_1_7 = (((mul2_84_port_byte_out_7 ^ mul3_84_port_byte_out_7) ^ port_state_in_6_1_7) ^ port_state_in_7_1_7);
  assign state_out_5_1_7 = (((mul2_85_port_byte_out_7 ^ mul3_85_port_byte_out_7) ^ port_state_in_4_1_7) ^ port_state_in_7_1_7);
  assign state_out_6_1_7 = (((mul2_86_port_byte_out_7 ^ mul3_86_port_byte_out_7) ^ port_state_in_4_1_7) ^ port_state_in_5_1_7);
  assign state_out_7_1_7 = (((mul2_87_port_byte_out_7 ^ mul3_87_port_byte_out_7) ^ port_state_in_5_1_7) ^ port_state_in_6_1_7);
  assign state_out_4_2_0 = (((mul2_88_port_byte_out_0 ^ mul3_88_port_byte_out_0) ^ port_state_in_6_2_0) ^ port_state_in_7_2_0);
  assign state_out_5_2_0 = (((mul2_89_port_byte_out_0 ^ mul3_89_port_byte_out_0) ^ port_state_in_4_2_0) ^ port_state_in_7_2_0);
  assign state_out_6_2_0 = (((mul2_90_port_byte_out_0 ^ mul3_90_port_byte_out_0) ^ port_state_in_4_2_0) ^ port_state_in_5_2_0);
  assign state_out_7_2_0 = (((mul2_91_port_byte_out_0 ^ mul3_91_port_byte_out_0) ^ port_state_in_5_2_0) ^ port_state_in_6_2_0);
  assign state_out_4_2_1 = (((mul2_88_port_byte_out_1 ^ mul3_88_port_byte_out_1) ^ port_state_in_6_2_1) ^ port_state_in_7_2_1);
  assign state_out_5_2_1 = (((mul2_89_port_byte_out_1 ^ mul3_89_port_byte_out_1) ^ port_state_in_4_2_1) ^ port_state_in_7_2_1);
  assign state_out_6_2_1 = (((mul2_90_port_byte_out_1 ^ mul3_90_port_byte_out_1) ^ port_state_in_4_2_1) ^ port_state_in_5_2_1);
  assign state_out_7_2_1 = (((mul2_91_port_byte_out_1 ^ mul3_91_port_byte_out_1) ^ port_state_in_5_2_1) ^ port_state_in_6_2_1);
  assign state_out_4_2_2 = (((mul2_88_port_byte_out_2 ^ mul3_88_port_byte_out_2) ^ port_state_in_6_2_2) ^ port_state_in_7_2_2);
  assign state_out_5_2_2 = (((mul2_89_port_byte_out_2 ^ mul3_89_port_byte_out_2) ^ port_state_in_4_2_2) ^ port_state_in_7_2_2);
  assign state_out_6_2_2 = (((mul2_90_port_byte_out_2 ^ mul3_90_port_byte_out_2) ^ port_state_in_4_2_2) ^ port_state_in_5_2_2);
  assign state_out_7_2_2 = (((mul2_91_port_byte_out_2 ^ mul3_91_port_byte_out_2) ^ port_state_in_5_2_2) ^ port_state_in_6_2_2);
  assign state_out_4_2_3 = (((mul2_88_port_byte_out_3 ^ mul3_88_port_byte_out_3) ^ port_state_in_6_2_3) ^ port_state_in_7_2_3);
  assign state_out_5_2_3 = (((mul2_89_port_byte_out_3 ^ mul3_89_port_byte_out_3) ^ port_state_in_4_2_3) ^ port_state_in_7_2_3);
  assign state_out_6_2_3 = (((mul2_90_port_byte_out_3 ^ mul3_90_port_byte_out_3) ^ port_state_in_4_2_3) ^ port_state_in_5_2_3);
  assign state_out_7_2_3 = (((mul2_91_port_byte_out_3 ^ mul3_91_port_byte_out_3) ^ port_state_in_5_2_3) ^ port_state_in_6_2_3);
  assign state_out_4_2_4 = (((mul2_88_port_byte_out_4 ^ mul3_88_port_byte_out_4) ^ port_state_in_6_2_4) ^ port_state_in_7_2_4);
  assign state_out_5_2_4 = (((mul2_89_port_byte_out_4 ^ mul3_89_port_byte_out_4) ^ port_state_in_4_2_4) ^ port_state_in_7_2_4);
  assign state_out_6_2_4 = (((mul2_90_port_byte_out_4 ^ mul3_90_port_byte_out_4) ^ port_state_in_4_2_4) ^ port_state_in_5_2_4);
  assign state_out_7_2_4 = (((mul2_91_port_byte_out_4 ^ mul3_91_port_byte_out_4) ^ port_state_in_5_2_4) ^ port_state_in_6_2_4);
  assign state_out_4_2_5 = (((mul2_88_port_byte_out_5 ^ mul3_88_port_byte_out_5) ^ port_state_in_6_2_5) ^ port_state_in_7_2_5);
  assign state_out_5_2_5 = (((mul2_89_port_byte_out_5 ^ mul3_89_port_byte_out_5) ^ port_state_in_4_2_5) ^ port_state_in_7_2_5);
  assign state_out_6_2_5 = (((mul2_90_port_byte_out_5 ^ mul3_90_port_byte_out_5) ^ port_state_in_4_2_5) ^ port_state_in_5_2_5);
  assign state_out_7_2_5 = (((mul2_91_port_byte_out_5 ^ mul3_91_port_byte_out_5) ^ port_state_in_5_2_5) ^ port_state_in_6_2_5);
  assign state_out_4_2_6 = (((mul2_88_port_byte_out_6 ^ mul3_88_port_byte_out_6) ^ port_state_in_6_2_6) ^ port_state_in_7_2_6);
  assign state_out_5_2_6 = (((mul2_89_port_byte_out_6 ^ mul3_89_port_byte_out_6) ^ port_state_in_4_2_6) ^ port_state_in_7_2_6);
  assign state_out_6_2_6 = (((mul2_90_port_byte_out_6 ^ mul3_90_port_byte_out_6) ^ port_state_in_4_2_6) ^ port_state_in_5_2_6);
  assign state_out_7_2_6 = (((mul2_91_port_byte_out_6 ^ mul3_91_port_byte_out_6) ^ port_state_in_5_2_6) ^ port_state_in_6_2_6);
  assign state_out_4_2_7 = (((mul2_88_port_byte_out_7 ^ mul3_88_port_byte_out_7) ^ port_state_in_6_2_7) ^ port_state_in_7_2_7);
  assign state_out_5_2_7 = (((mul2_89_port_byte_out_7 ^ mul3_89_port_byte_out_7) ^ port_state_in_4_2_7) ^ port_state_in_7_2_7);
  assign state_out_6_2_7 = (((mul2_90_port_byte_out_7 ^ mul3_90_port_byte_out_7) ^ port_state_in_4_2_7) ^ port_state_in_5_2_7);
  assign state_out_7_2_7 = (((mul2_91_port_byte_out_7 ^ mul3_91_port_byte_out_7) ^ port_state_in_5_2_7) ^ port_state_in_6_2_7);
  assign state_out_4_3_0 = (((mul2_92_port_byte_out_0 ^ mul3_92_port_byte_out_0) ^ port_state_in_6_3_0) ^ port_state_in_7_3_0);
  assign state_out_5_3_0 = (((mul2_93_port_byte_out_0 ^ mul3_93_port_byte_out_0) ^ port_state_in_4_3_0) ^ port_state_in_7_3_0);
  assign state_out_6_3_0 = (((mul2_94_port_byte_out_0 ^ mul3_94_port_byte_out_0) ^ port_state_in_4_3_0) ^ port_state_in_5_3_0);
  assign state_out_7_3_0 = (((mul2_95_port_byte_out_0 ^ mul3_95_port_byte_out_0) ^ port_state_in_5_3_0) ^ port_state_in_6_3_0);
  assign state_out_4_3_1 = (((mul2_92_port_byte_out_1 ^ mul3_92_port_byte_out_1) ^ port_state_in_6_3_1) ^ port_state_in_7_3_1);
  assign state_out_5_3_1 = (((mul2_93_port_byte_out_1 ^ mul3_93_port_byte_out_1) ^ port_state_in_4_3_1) ^ port_state_in_7_3_1);
  assign state_out_6_3_1 = (((mul2_94_port_byte_out_1 ^ mul3_94_port_byte_out_1) ^ port_state_in_4_3_1) ^ port_state_in_5_3_1);
  assign state_out_7_3_1 = (((mul2_95_port_byte_out_1 ^ mul3_95_port_byte_out_1) ^ port_state_in_5_3_1) ^ port_state_in_6_3_1);
  assign state_out_4_3_2 = (((mul2_92_port_byte_out_2 ^ mul3_92_port_byte_out_2) ^ port_state_in_6_3_2) ^ port_state_in_7_3_2);
  assign state_out_5_3_2 = (((mul2_93_port_byte_out_2 ^ mul3_93_port_byte_out_2) ^ port_state_in_4_3_2) ^ port_state_in_7_3_2);
  assign state_out_6_3_2 = (((mul2_94_port_byte_out_2 ^ mul3_94_port_byte_out_2) ^ port_state_in_4_3_2) ^ port_state_in_5_3_2);
  assign state_out_7_3_2 = (((mul2_95_port_byte_out_2 ^ mul3_95_port_byte_out_2) ^ port_state_in_5_3_2) ^ port_state_in_6_3_2);
  assign state_out_4_3_3 = (((mul2_92_port_byte_out_3 ^ mul3_92_port_byte_out_3) ^ port_state_in_6_3_3) ^ port_state_in_7_3_3);
  assign state_out_5_3_3 = (((mul2_93_port_byte_out_3 ^ mul3_93_port_byte_out_3) ^ port_state_in_4_3_3) ^ port_state_in_7_3_3);
  assign state_out_6_3_3 = (((mul2_94_port_byte_out_3 ^ mul3_94_port_byte_out_3) ^ port_state_in_4_3_3) ^ port_state_in_5_3_3);
  assign state_out_7_3_3 = (((mul2_95_port_byte_out_3 ^ mul3_95_port_byte_out_3) ^ port_state_in_5_3_3) ^ port_state_in_6_3_3);
  assign state_out_4_3_4 = (((mul2_92_port_byte_out_4 ^ mul3_92_port_byte_out_4) ^ port_state_in_6_3_4) ^ port_state_in_7_3_4);
  assign state_out_5_3_4 = (((mul2_93_port_byte_out_4 ^ mul3_93_port_byte_out_4) ^ port_state_in_4_3_4) ^ port_state_in_7_3_4);
  assign state_out_6_3_4 = (((mul2_94_port_byte_out_4 ^ mul3_94_port_byte_out_4) ^ port_state_in_4_3_4) ^ port_state_in_5_3_4);
  assign state_out_7_3_4 = (((mul2_95_port_byte_out_4 ^ mul3_95_port_byte_out_4) ^ port_state_in_5_3_4) ^ port_state_in_6_3_4);
  assign state_out_4_3_5 = (((mul2_92_port_byte_out_5 ^ mul3_92_port_byte_out_5) ^ port_state_in_6_3_5) ^ port_state_in_7_3_5);
  assign state_out_5_3_5 = (((mul2_93_port_byte_out_5 ^ mul3_93_port_byte_out_5) ^ port_state_in_4_3_5) ^ port_state_in_7_3_5);
  assign state_out_6_3_5 = (((mul2_94_port_byte_out_5 ^ mul3_94_port_byte_out_5) ^ port_state_in_4_3_5) ^ port_state_in_5_3_5);
  assign state_out_7_3_5 = (((mul2_95_port_byte_out_5 ^ mul3_95_port_byte_out_5) ^ port_state_in_5_3_5) ^ port_state_in_6_3_5);
  assign state_out_4_3_6 = (((mul2_92_port_byte_out_6 ^ mul3_92_port_byte_out_6) ^ port_state_in_6_3_6) ^ port_state_in_7_3_6);
  assign state_out_5_3_6 = (((mul2_93_port_byte_out_6 ^ mul3_93_port_byte_out_6) ^ port_state_in_4_3_6) ^ port_state_in_7_3_6);
  assign state_out_6_3_6 = (((mul2_94_port_byte_out_6 ^ mul3_94_port_byte_out_6) ^ port_state_in_4_3_6) ^ port_state_in_5_3_6);
  assign state_out_7_3_6 = (((mul2_95_port_byte_out_6 ^ mul3_95_port_byte_out_6) ^ port_state_in_5_3_6) ^ port_state_in_6_3_6);
  assign state_out_4_3_7 = (((mul2_92_port_byte_out_7 ^ mul3_92_port_byte_out_7) ^ port_state_in_6_3_7) ^ port_state_in_7_3_7);
  assign state_out_5_3_7 = (((mul2_93_port_byte_out_7 ^ mul3_93_port_byte_out_7) ^ port_state_in_4_3_7) ^ port_state_in_7_3_7);
  assign state_out_6_3_7 = (((mul2_94_port_byte_out_7 ^ mul3_94_port_byte_out_7) ^ port_state_in_4_3_7) ^ port_state_in_5_3_7);
  assign state_out_7_3_7 = (((mul2_95_port_byte_out_7 ^ mul3_95_port_byte_out_7) ^ port_state_in_5_3_7) ^ port_state_in_6_3_7);
  assign state_out_8_0_0 = (((mul2_96_port_byte_out_0 ^ mul3_96_port_byte_out_0) ^ port_state_in_10_0_0) ^ port_state_in_11_0_0);
  assign state_out_9_0_0 = (((mul2_97_port_byte_out_0 ^ mul3_97_port_byte_out_0) ^ port_state_in_8_0_0) ^ port_state_in_11_0_0);
  assign state_out_10_0_0 = (((mul2_98_port_byte_out_0 ^ mul3_98_port_byte_out_0) ^ port_state_in_8_0_0) ^ port_state_in_9_0_0);
  assign state_out_11_0_0 = (((mul2_99_port_byte_out_0 ^ mul3_99_port_byte_out_0) ^ port_state_in_9_0_0) ^ port_state_in_10_0_0);
  assign state_out_8_0_1 = (((mul2_96_port_byte_out_1 ^ mul3_96_port_byte_out_1) ^ port_state_in_10_0_1) ^ port_state_in_11_0_1);
  assign state_out_9_0_1 = (((mul2_97_port_byte_out_1 ^ mul3_97_port_byte_out_1) ^ port_state_in_8_0_1) ^ port_state_in_11_0_1);
  assign state_out_10_0_1 = (((mul2_98_port_byte_out_1 ^ mul3_98_port_byte_out_1) ^ port_state_in_8_0_1) ^ port_state_in_9_0_1);
  assign state_out_11_0_1 = (((mul2_99_port_byte_out_1 ^ mul3_99_port_byte_out_1) ^ port_state_in_9_0_1) ^ port_state_in_10_0_1);
  assign state_out_8_0_2 = (((mul2_96_port_byte_out_2 ^ mul3_96_port_byte_out_2) ^ port_state_in_10_0_2) ^ port_state_in_11_0_2);
  assign state_out_9_0_2 = (((mul2_97_port_byte_out_2 ^ mul3_97_port_byte_out_2) ^ port_state_in_8_0_2) ^ port_state_in_11_0_2);
  assign state_out_10_0_2 = (((mul2_98_port_byte_out_2 ^ mul3_98_port_byte_out_2) ^ port_state_in_8_0_2) ^ port_state_in_9_0_2);
  assign state_out_11_0_2 = (((mul2_99_port_byte_out_2 ^ mul3_99_port_byte_out_2) ^ port_state_in_9_0_2) ^ port_state_in_10_0_2);
  assign state_out_8_0_3 = (((mul2_96_port_byte_out_3 ^ mul3_96_port_byte_out_3) ^ port_state_in_10_0_3) ^ port_state_in_11_0_3);
  assign state_out_9_0_3 = (((mul2_97_port_byte_out_3 ^ mul3_97_port_byte_out_3) ^ port_state_in_8_0_3) ^ port_state_in_11_0_3);
  assign state_out_10_0_3 = (((mul2_98_port_byte_out_3 ^ mul3_98_port_byte_out_3) ^ port_state_in_8_0_3) ^ port_state_in_9_0_3);
  assign state_out_11_0_3 = (((mul2_99_port_byte_out_3 ^ mul3_99_port_byte_out_3) ^ port_state_in_9_0_3) ^ port_state_in_10_0_3);
  assign state_out_8_0_4 = (((mul2_96_port_byte_out_4 ^ mul3_96_port_byte_out_4) ^ port_state_in_10_0_4) ^ port_state_in_11_0_4);
  assign state_out_9_0_4 = (((mul2_97_port_byte_out_4 ^ mul3_97_port_byte_out_4) ^ port_state_in_8_0_4) ^ port_state_in_11_0_4);
  assign state_out_10_0_4 = (((mul2_98_port_byte_out_4 ^ mul3_98_port_byte_out_4) ^ port_state_in_8_0_4) ^ port_state_in_9_0_4);
  assign state_out_11_0_4 = (((mul2_99_port_byte_out_4 ^ mul3_99_port_byte_out_4) ^ port_state_in_9_0_4) ^ port_state_in_10_0_4);
  assign state_out_8_0_5 = (((mul2_96_port_byte_out_5 ^ mul3_96_port_byte_out_5) ^ port_state_in_10_0_5) ^ port_state_in_11_0_5);
  assign state_out_9_0_5 = (((mul2_97_port_byte_out_5 ^ mul3_97_port_byte_out_5) ^ port_state_in_8_0_5) ^ port_state_in_11_0_5);
  assign state_out_10_0_5 = (((mul2_98_port_byte_out_5 ^ mul3_98_port_byte_out_5) ^ port_state_in_8_0_5) ^ port_state_in_9_0_5);
  assign state_out_11_0_5 = (((mul2_99_port_byte_out_5 ^ mul3_99_port_byte_out_5) ^ port_state_in_9_0_5) ^ port_state_in_10_0_5);
  assign state_out_8_0_6 = (((mul2_96_port_byte_out_6 ^ mul3_96_port_byte_out_6) ^ port_state_in_10_0_6) ^ port_state_in_11_0_6);
  assign state_out_9_0_6 = (((mul2_97_port_byte_out_6 ^ mul3_97_port_byte_out_6) ^ port_state_in_8_0_6) ^ port_state_in_11_0_6);
  assign state_out_10_0_6 = (((mul2_98_port_byte_out_6 ^ mul3_98_port_byte_out_6) ^ port_state_in_8_0_6) ^ port_state_in_9_0_6);
  assign state_out_11_0_6 = (((mul2_99_port_byte_out_6 ^ mul3_99_port_byte_out_6) ^ port_state_in_9_0_6) ^ port_state_in_10_0_6);
  assign state_out_8_0_7 = (((mul2_96_port_byte_out_7 ^ mul3_96_port_byte_out_7) ^ port_state_in_10_0_7) ^ port_state_in_11_0_7);
  assign state_out_9_0_7 = (((mul2_97_port_byte_out_7 ^ mul3_97_port_byte_out_7) ^ port_state_in_8_0_7) ^ port_state_in_11_0_7);
  assign state_out_10_0_7 = (((mul2_98_port_byte_out_7 ^ mul3_98_port_byte_out_7) ^ port_state_in_8_0_7) ^ port_state_in_9_0_7);
  assign state_out_11_0_7 = (((mul2_99_port_byte_out_7 ^ mul3_99_port_byte_out_7) ^ port_state_in_9_0_7) ^ port_state_in_10_0_7);
  assign state_out_8_1_0 = (((mul2_100_port_byte_out_0 ^ mul3_100_port_byte_out_0) ^ port_state_in_10_1_0) ^ port_state_in_11_1_0);
  assign state_out_9_1_0 = (((mul2_101_port_byte_out_0 ^ mul3_101_port_byte_out_0) ^ port_state_in_8_1_0) ^ port_state_in_11_1_0);
  assign state_out_10_1_0 = (((mul2_102_port_byte_out_0 ^ mul3_102_port_byte_out_0) ^ port_state_in_8_1_0) ^ port_state_in_9_1_0);
  assign state_out_11_1_0 = (((mul2_103_port_byte_out_0 ^ mul3_103_port_byte_out_0) ^ port_state_in_9_1_0) ^ port_state_in_10_1_0);
  assign state_out_8_1_1 = (((mul2_100_port_byte_out_1 ^ mul3_100_port_byte_out_1) ^ port_state_in_10_1_1) ^ port_state_in_11_1_1);
  assign state_out_9_1_1 = (((mul2_101_port_byte_out_1 ^ mul3_101_port_byte_out_1) ^ port_state_in_8_1_1) ^ port_state_in_11_1_1);
  assign state_out_10_1_1 = (((mul2_102_port_byte_out_1 ^ mul3_102_port_byte_out_1) ^ port_state_in_8_1_1) ^ port_state_in_9_1_1);
  assign state_out_11_1_1 = (((mul2_103_port_byte_out_1 ^ mul3_103_port_byte_out_1) ^ port_state_in_9_1_1) ^ port_state_in_10_1_1);
  assign state_out_8_1_2 = (((mul2_100_port_byte_out_2 ^ mul3_100_port_byte_out_2) ^ port_state_in_10_1_2) ^ port_state_in_11_1_2);
  assign state_out_9_1_2 = (((mul2_101_port_byte_out_2 ^ mul3_101_port_byte_out_2) ^ port_state_in_8_1_2) ^ port_state_in_11_1_2);
  assign state_out_10_1_2 = (((mul2_102_port_byte_out_2 ^ mul3_102_port_byte_out_2) ^ port_state_in_8_1_2) ^ port_state_in_9_1_2);
  assign state_out_11_1_2 = (((mul2_103_port_byte_out_2 ^ mul3_103_port_byte_out_2) ^ port_state_in_9_1_2) ^ port_state_in_10_1_2);
  assign state_out_8_1_3 = (((mul2_100_port_byte_out_3 ^ mul3_100_port_byte_out_3) ^ port_state_in_10_1_3) ^ port_state_in_11_1_3);
  assign state_out_9_1_3 = (((mul2_101_port_byte_out_3 ^ mul3_101_port_byte_out_3) ^ port_state_in_8_1_3) ^ port_state_in_11_1_3);
  assign state_out_10_1_3 = (((mul2_102_port_byte_out_3 ^ mul3_102_port_byte_out_3) ^ port_state_in_8_1_3) ^ port_state_in_9_1_3);
  assign state_out_11_1_3 = (((mul2_103_port_byte_out_3 ^ mul3_103_port_byte_out_3) ^ port_state_in_9_1_3) ^ port_state_in_10_1_3);
  assign state_out_8_1_4 = (((mul2_100_port_byte_out_4 ^ mul3_100_port_byte_out_4) ^ port_state_in_10_1_4) ^ port_state_in_11_1_4);
  assign state_out_9_1_4 = (((mul2_101_port_byte_out_4 ^ mul3_101_port_byte_out_4) ^ port_state_in_8_1_4) ^ port_state_in_11_1_4);
  assign state_out_10_1_4 = (((mul2_102_port_byte_out_4 ^ mul3_102_port_byte_out_4) ^ port_state_in_8_1_4) ^ port_state_in_9_1_4);
  assign state_out_11_1_4 = (((mul2_103_port_byte_out_4 ^ mul3_103_port_byte_out_4) ^ port_state_in_9_1_4) ^ port_state_in_10_1_4);
  assign state_out_8_1_5 = (((mul2_100_port_byte_out_5 ^ mul3_100_port_byte_out_5) ^ port_state_in_10_1_5) ^ port_state_in_11_1_5);
  assign state_out_9_1_5 = (((mul2_101_port_byte_out_5 ^ mul3_101_port_byte_out_5) ^ port_state_in_8_1_5) ^ port_state_in_11_1_5);
  assign state_out_10_1_5 = (((mul2_102_port_byte_out_5 ^ mul3_102_port_byte_out_5) ^ port_state_in_8_1_5) ^ port_state_in_9_1_5);
  assign state_out_11_1_5 = (((mul2_103_port_byte_out_5 ^ mul3_103_port_byte_out_5) ^ port_state_in_9_1_5) ^ port_state_in_10_1_5);
  assign state_out_8_1_6 = (((mul2_100_port_byte_out_6 ^ mul3_100_port_byte_out_6) ^ port_state_in_10_1_6) ^ port_state_in_11_1_6);
  assign state_out_9_1_6 = (((mul2_101_port_byte_out_6 ^ mul3_101_port_byte_out_6) ^ port_state_in_8_1_6) ^ port_state_in_11_1_6);
  assign state_out_10_1_6 = (((mul2_102_port_byte_out_6 ^ mul3_102_port_byte_out_6) ^ port_state_in_8_1_6) ^ port_state_in_9_1_6);
  assign state_out_11_1_6 = (((mul2_103_port_byte_out_6 ^ mul3_103_port_byte_out_6) ^ port_state_in_9_1_6) ^ port_state_in_10_1_6);
  assign state_out_8_1_7 = (((mul2_100_port_byte_out_7 ^ mul3_100_port_byte_out_7) ^ port_state_in_10_1_7) ^ port_state_in_11_1_7);
  assign state_out_9_1_7 = (((mul2_101_port_byte_out_7 ^ mul3_101_port_byte_out_7) ^ port_state_in_8_1_7) ^ port_state_in_11_1_7);
  assign state_out_10_1_7 = (((mul2_102_port_byte_out_7 ^ mul3_102_port_byte_out_7) ^ port_state_in_8_1_7) ^ port_state_in_9_1_7);
  assign state_out_11_1_7 = (((mul2_103_port_byte_out_7 ^ mul3_103_port_byte_out_7) ^ port_state_in_9_1_7) ^ port_state_in_10_1_7);
  assign state_out_8_2_0 = (((mul2_104_port_byte_out_0 ^ mul3_104_port_byte_out_0) ^ port_state_in_10_2_0) ^ port_state_in_11_2_0);
  assign state_out_9_2_0 = (((mul2_105_port_byte_out_0 ^ mul3_105_port_byte_out_0) ^ port_state_in_8_2_0) ^ port_state_in_11_2_0);
  assign state_out_10_2_0 = (((mul2_106_port_byte_out_0 ^ mul3_106_port_byte_out_0) ^ port_state_in_8_2_0) ^ port_state_in_9_2_0);
  assign state_out_11_2_0 = (((mul2_107_port_byte_out_0 ^ mul3_107_port_byte_out_0) ^ port_state_in_9_2_0) ^ port_state_in_10_2_0);
  assign state_out_8_2_1 = (((mul2_104_port_byte_out_1 ^ mul3_104_port_byte_out_1) ^ port_state_in_10_2_1) ^ port_state_in_11_2_1);
  assign state_out_9_2_1 = (((mul2_105_port_byte_out_1 ^ mul3_105_port_byte_out_1) ^ port_state_in_8_2_1) ^ port_state_in_11_2_1);
  assign state_out_10_2_1 = (((mul2_106_port_byte_out_1 ^ mul3_106_port_byte_out_1) ^ port_state_in_8_2_1) ^ port_state_in_9_2_1);
  assign state_out_11_2_1 = (((mul2_107_port_byte_out_1 ^ mul3_107_port_byte_out_1) ^ port_state_in_9_2_1) ^ port_state_in_10_2_1);
  assign state_out_8_2_2 = (((mul2_104_port_byte_out_2 ^ mul3_104_port_byte_out_2) ^ port_state_in_10_2_2) ^ port_state_in_11_2_2);
  assign state_out_9_2_2 = (((mul2_105_port_byte_out_2 ^ mul3_105_port_byte_out_2) ^ port_state_in_8_2_2) ^ port_state_in_11_2_2);
  assign state_out_10_2_2 = (((mul2_106_port_byte_out_2 ^ mul3_106_port_byte_out_2) ^ port_state_in_8_2_2) ^ port_state_in_9_2_2);
  assign state_out_11_2_2 = (((mul2_107_port_byte_out_2 ^ mul3_107_port_byte_out_2) ^ port_state_in_9_2_2) ^ port_state_in_10_2_2);
  assign state_out_8_2_3 = (((mul2_104_port_byte_out_3 ^ mul3_104_port_byte_out_3) ^ port_state_in_10_2_3) ^ port_state_in_11_2_3);
  assign state_out_9_2_3 = (((mul2_105_port_byte_out_3 ^ mul3_105_port_byte_out_3) ^ port_state_in_8_2_3) ^ port_state_in_11_2_3);
  assign state_out_10_2_3 = (((mul2_106_port_byte_out_3 ^ mul3_106_port_byte_out_3) ^ port_state_in_8_2_3) ^ port_state_in_9_2_3);
  assign state_out_11_2_3 = (((mul2_107_port_byte_out_3 ^ mul3_107_port_byte_out_3) ^ port_state_in_9_2_3) ^ port_state_in_10_2_3);
  assign state_out_8_2_4 = (((mul2_104_port_byte_out_4 ^ mul3_104_port_byte_out_4) ^ port_state_in_10_2_4) ^ port_state_in_11_2_4);
  assign state_out_9_2_4 = (((mul2_105_port_byte_out_4 ^ mul3_105_port_byte_out_4) ^ port_state_in_8_2_4) ^ port_state_in_11_2_4);
  assign state_out_10_2_4 = (((mul2_106_port_byte_out_4 ^ mul3_106_port_byte_out_4) ^ port_state_in_8_2_4) ^ port_state_in_9_2_4);
  assign state_out_11_2_4 = (((mul2_107_port_byte_out_4 ^ mul3_107_port_byte_out_4) ^ port_state_in_9_2_4) ^ port_state_in_10_2_4);
  assign state_out_8_2_5 = (((mul2_104_port_byte_out_5 ^ mul3_104_port_byte_out_5) ^ port_state_in_10_2_5) ^ port_state_in_11_2_5);
  assign state_out_9_2_5 = (((mul2_105_port_byte_out_5 ^ mul3_105_port_byte_out_5) ^ port_state_in_8_2_5) ^ port_state_in_11_2_5);
  assign state_out_10_2_5 = (((mul2_106_port_byte_out_5 ^ mul3_106_port_byte_out_5) ^ port_state_in_8_2_5) ^ port_state_in_9_2_5);
  assign state_out_11_2_5 = (((mul2_107_port_byte_out_5 ^ mul3_107_port_byte_out_5) ^ port_state_in_9_2_5) ^ port_state_in_10_2_5);
  assign state_out_8_2_6 = (((mul2_104_port_byte_out_6 ^ mul3_104_port_byte_out_6) ^ port_state_in_10_2_6) ^ port_state_in_11_2_6);
  assign state_out_9_2_6 = (((mul2_105_port_byte_out_6 ^ mul3_105_port_byte_out_6) ^ port_state_in_8_2_6) ^ port_state_in_11_2_6);
  assign state_out_10_2_6 = (((mul2_106_port_byte_out_6 ^ mul3_106_port_byte_out_6) ^ port_state_in_8_2_6) ^ port_state_in_9_2_6);
  assign state_out_11_2_6 = (((mul2_107_port_byte_out_6 ^ mul3_107_port_byte_out_6) ^ port_state_in_9_2_6) ^ port_state_in_10_2_6);
  assign state_out_8_2_7 = (((mul2_104_port_byte_out_7 ^ mul3_104_port_byte_out_7) ^ port_state_in_10_2_7) ^ port_state_in_11_2_7);
  assign state_out_9_2_7 = (((mul2_105_port_byte_out_7 ^ mul3_105_port_byte_out_7) ^ port_state_in_8_2_7) ^ port_state_in_11_2_7);
  assign state_out_10_2_7 = (((mul2_106_port_byte_out_7 ^ mul3_106_port_byte_out_7) ^ port_state_in_8_2_7) ^ port_state_in_9_2_7);
  assign state_out_11_2_7 = (((mul2_107_port_byte_out_7 ^ mul3_107_port_byte_out_7) ^ port_state_in_9_2_7) ^ port_state_in_10_2_7);
  assign state_out_8_3_0 = (((mul2_108_port_byte_out_0 ^ mul3_108_port_byte_out_0) ^ port_state_in_10_3_0) ^ port_state_in_11_3_0);
  assign state_out_9_3_0 = (((mul2_109_port_byte_out_0 ^ mul3_109_port_byte_out_0) ^ port_state_in_8_3_0) ^ port_state_in_11_3_0);
  assign state_out_10_3_0 = (((mul2_110_port_byte_out_0 ^ mul3_110_port_byte_out_0) ^ port_state_in_8_3_0) ^ port_state_in_9_3_0);
  assign state_out_11_3_0 = (((mul2_111_port_byte_out_0 ^ mul3_111_port_byte_out_0) ^ port_state_in_9_3_0) ^ port_state_in_10_3_0);
  assign state_out_8_3_1 = (((mul2_108_port_byte_out_1 ^ mul3_108_port_byte_out_1) ^ port_state_in_10_3_1) ^ port_state_in_11_3_1);
  assign state_out_9_3_1 = (((mul2_109_port_byte_out_1 ^ mul3_109_port_byte_out_1) ^ port_state_in_8_3_1) ^ port_state_in_11_3_1);
  assign state_out_10_3_1 = (((mul2_110_port_byte_out_1 ^ mul3_110_port_byte_out_1) ^ port_state_in_8_3_1) ^ port_state_in_9_3_1);
  assign state_out_11_3_1 = (((mul2_111_port_byte_out_1 ^ mul3_111_port_byte_out_1) ^ port_state_in_9_3_1) ^ port_state_in_10_3_1);
  assign state_out_8_3_2 = (((mul2_108_port_byte_out_2 ^ mul3_108_port_byte_out_2) ^ port_state_in_10_3_2) ^ port_state_in_11_3_2);
  assign state_out_9_3_2 = (((mul2_109_port_byte_out_2 ^ mul3_109_port_byte_out_2) ^ port_state_in_8_3_2) ^ port_state_in_11_3_2);
  assign state_out_10_3_2 = (((mul2_110_port_byte_out_2 ^ mul3_110_port_byte_out_2) ^ port_state_in_8_3_2) ^ port_state_in_9_3_2);
  assign state_out_11_3_2 = (((mul2_111_port_byte_out_2 ^ mul3_111_port_byte_out_2) ^ port_state_in_9_3_2) ^ port_state_in_10_3_2);
  assign state_out_8_3_3 = (((mul2_108_port_byte_out_3 ^ mul3_108_port_byte_out_3) ^ port_state_in_10_3_3) ^ port_state_in_11_3_3);
  assign state_out_9_3_3 = (((mul2_109_port_byte_out_3 ^ mul3_109_port_byte_out_3) ^ port_state_in_8_3_3) ^ port_state_in_11_3_3);
  assign state_out_10_3_3 = (((mul2_110_port_byte_out_3 ^ mul3_110_port_byte_out_3) ^ port_state_in_8_3_3) ^ port_state_in_9_3_3);
  assign state_out_11_3_3 = (((mul2_111_port_byte_out_3 ^ mul3_111_port_byte_out_3) ^ port_state_in_9_3_3) ^ port_state_in_10_3_3);
  assign state_out_8_3_4 = (((mul2_108_port_byte_out_4 ^ mul3_108_port_byte_out_4) ^ port_state_in_10_3_4) ^ port_state_in_11_3_4);
  assign state_out_9_3_4 = (((mul2_109_port_byte_out_4 ^ mul3_109_port_byte_out_4) ^ port_state_in_8_3_4) ^ port_state_in_11_3_4);
  assign state_out_10_3_4 = (((mul2_110_port_byte_out_4 ^ mul3_110_port_byte_out_4) ^ port_state_in_8_3_4) ^ port_state_in_9_3_4);
  assign state_out_11_3_4 = (((mul2_111_port_byte_out_4 ^ mul3_111_port_byte_out_4) ^ port_state_in_9_3_4) ^ port_state_in_10_3_4);
  assign state_out_8_3_5 = (((mul2_108_port_byte_out_5 ^ mul3_108_port_byte_out_5) ^ port_state_in_10_3_5) ^ port_state_in_11_3_5);
  assign state_out_9_3_5 = (((mul2_109_port_byte_out_5 ^ mul3_109_port_byte_out_5) ^ port_state_in_8_3_5) ^ port_state_in_11_3_5);
  assign state_out_10_3_5 = (((mul2_110_port_byte_out_5 ^ mul3_110_port_byte_out_5) ^ port_state_in_8_3_5) ^ port_state_in_9_3_5);
  assign state_out_11_3_5 = (((mul2_111_port_byte_out_5 ^ mul3_111_port_byte_out_5) ^ port_state_in_9_3_5) ^ port_state_in_10_3_5);
  assign state_out_8_3_6 = (((mul2_108_port_byte_out_6 ^ mul3_108_port_byte_out_6) ^ port_state_in_10_3_6) ^ port_state_in_11_3_6);
  assign state_out_9_3_6 = (((mul2_109_port_byte_out_6 ^ mul3_109_port_byte_out_6) ^ port_state_in_8_3_6) ^ port_state_in_11_3_6);
  assign state_out_10_3_6 = (((mul2_110_port_byte_out_6 ^ mul3_110_port_byte_out_6) ^ port_state_in_8_3_6) ^ port_state_in_9_3_6);
  assign state_out_11_3_6 = (((mul2_111_port_byte_out_6 ^ mul3_111_port_byte_out_6) ^ port_state_in_9_3_6) ^ port_state_in_10_3_6);
  assign state_out_8_3_7 = (((mul2_108_port_byte_out_7 ^ mul3_108_port_byte_out_7) ^ port_state_in_10_3_7) ^ port_state_in_11_3_7);
  assign state_out_9_3_7 = (((mul2_109_port_byte_out_7 ^ mul3_109_port_byte_out_7) ^ port_state_in_8_3_7) ^ port_state_in_11_3_7);
  assign state_out_10_3_7 = (((mul2_110_port_byte_out_7 ^ mul3_110_port_byte_out_7) ^ port_state_in_8_3_7) ^ port_state_in_9_3_7);
  assign state_out_11_3_7 = (((mul2_111_port_byte_out_7 ^ mul3_111_port_byte_out_7) ^ port_state_in_9_3_7) ^ port_state_in_10_3_7);
  assign state_out_12_0_0 = (((mul2_112_port_byte_out_0 ^ mul3_112_port_byte_out_0) ^ port_state_in_14_0_0) ^ port_state_in_15_0_0);
  assign state_out_13_0_0 = (((mul2_113_port_byte_out_0 ^ mul3_113_port_byte_out_0) ^ port_state_in_12_0_0) ^ port_state_in_15_0_0);
  assign state_out_14_0_0 = (((mul2_114_port_byte_out_0 ^ mul3_114_port_byte_out_0) ^ port_state_in_12_0_0) ^ port_state_in_13_0_0);
  assign state_out_15_0_0 = (((mul2_115_port_byte_out_0 ^ mul3_115_port_byte_out_0) ^ port_state_in_13_0_0) ^ port_state_in_14_0_0);
  assign state_out_12_0_1 = (((mul2_112_port_byte_out_1 ^ mul3_112_port_byte_out_1) ^ port_state_in_14_0_1) ^ port_state_in_15_0_1);
  assign state_out_13_0_1 = (((mul2_113_port_byte_out_1 ^ mul3_113_port_byte_out_1) ^ port_state_in_12_0_1) ^ port_state_in_15_0_1);
  assign state_out_14_0_1 = (((mul2_114_port_byte_out_1 ^ mul3_114_port_byte_out_1) ^ port_state_in_12_0_1) ^ port_state_in_13_0_1);
  assign state_out_15_0_1 = (((mul2_115_port_byte_out_1 ^ mul3_115_port_byte_out_1) ^ port_state_in_13_0_1) ^ port_state_in_14_0_1);
  assign state_out_12_0_2 = (((mul2_112_port_byte_out_2 ^ mul3_112_port_byte_out_2) ^ port_state_in_14_0_2) ^ port_state_in_15_0_2);
  assign state_out_13_0_2 = (((mul2_113_port_byte_out_2 ^ mul3_113_port_byte_out_2) ^ port_state_in_12_0_2) ^ port_state_in_15_0_2);
  assign state_out_14_0_2 = (((mul2_114_port_byte_out_2 ^ mul3_114_port_byte_out_2) ^ port_state_in_12_0_2) ^ port_state_in_13_0_2);
  assign state_out_15_0_2 = (((mul2_115_port_byte_out_2 ^ mul3_115_port_byte_out_2) ^ port_state_in_13_0_2) ^ port_state_in_14_0_2);
  assign state_out_12_0_3 = (((mul2_112_port_byte_out_3 ^ mul3_112_port_byte_out_3) ^ port_state_in_14_0_3) ^ port_state_in_15_0_3);
  assign state_out_13_0_3 = (((mul2_113_port_byte_out_3 ^ mul3_113_port_byte_out_3) ^ port_state_in_12_0_3) ^ port_state_in_15_0_3);
  assign state_out_14_0_3 = (((mul2_114_port_byte_out_3 ^ mul3_114_port_byte_out_3) ^ port_state_in_12_0_3) ^ port_state_in_13_0_3);
  assign state_out_15_0_3 = (((mul2_115_port_byte_out_3 ^ mul3_115_port_byte_out_3) ^ port_state_in_13_0_3) ^ port_state_in_14_0_3);
  assign state_out_12_0_4 = (((mul2_112_port_byte_out_4 ^ mul3_112_port_byte_out_4) ^ port_state_in_14_0_4) ^ port_state_in_15_0_4);
  assign state_out_13_0_4 = (((mul2_113_port_byte_out_4 ^ mul3_113_port_byte_out_4) ^ port_state_in_12_0_4) ^ port_state_in_15_0_4);
  assign state_out_14_0_4 = (((mul2_114_port_byte_out_4 ^ mul3_114_port_byte_out_4) ^ port_state_in_12_0_4) ^ port_state_in_13_0_4);
  assign state_out_15_0_4 = (((mul2_115_port_byte_out_4 ^ mul3_115_port_byte_out_4) ^ port_state_in_13_0_4) ^ port_state_in_14_0_4);
  assign state_out_12_0_5 = (((mul2_112_port_byte_out_5 ^ mul3_112_port_byte_out_5) ^ port_state_in_14_0_5) ^ port_state_in_15_0_5);
  assign state_out_13_0_5 = (((mul2_113_port_byte_out_5 ^ mul3_113_port_byte_out_5) ^ port_state_in_12_0_5) ^ port_state_in_15_0_5);
  assign state_out_14_0_5 = (((mul2_114_port_byte_out_5 ^ mul3_114_port_byte_out_5) ^ port_state_in_12_0_5) ^ port_state_in_13_0_5);
  assign state_out_15_0_5 = (((mul2_115_port_byte_out_5 ^ mul3_115_port_byte_out_5) ^ port_state_in_13_0_5) ^ port_state_in_14_0_5);
  assign state_out_12_0_6 = (((mul2_112_port_byte_out_6 ^ mul3_112_port_byte_out_6) ^ port_state_in_14_0_6) ^ port_state_in_15_0_6);
  assign state_out_13_0_6 = (((mul2_113_port_byte_out_6 ^ mul3_113_port_byte_out_6) ^ port_state_in_12_0_6) ^ port_state_in_15_0_6);
  assign state_out_14_0_6 = (((mul2_114_port_byte_out_6 ^ mul3_114_port_byte_out_6) ^ port_state_in_12_0_6) ^ port_state_in_13_0_6);
  assign state_out_15_0_6 = (((mul2_115_port_byte_out_6 ^ mul3_115_port_byte_out_6) ^ port_state_in_13_0_6) ^ port_state_in_14_0_6);
  assign state_out_12_0_7 = (((mul2_112_port_byte_out_7 ^ mul3_112_port_byte_out_7) ^ port_state_in_14_0_7) ^ port_state_in_15_0_7);
  assign state_out_13_0_7 = (((mul2_113_port_byte_out_7 ^ mul3_113_port_byte_out_7) ^ port_state_in_12_0_7) ^ port_state_in_15_0_7);
  assign state_out_14_0_7 = (((mul2_114_port_byte_out_7 ^ mul3_114_port_byte_out_7) ^ port_state_in_12_0_7) ^ port_state_in_13_0_7);
  assign state_out_15_0_7 = (((mul2_115_port_byte_out_7 ^ mul3_115_port_byte_out_7) ^ port_state_in_13_0_7) ^ port_state_in_14_0_7);
  assign state_out_12_1_0 = (((mul2_116_port_byte_out_0 ^ mul3_116_port_byte_out_0) ^ port_state_in_14_1_0) ^ port_state_in_15_1_0);
  assign state_out_13_1_0 = (((mul2_117_port_byte_out_0 ^ mul3_117_port_byte_out_0) ^ port_state_in_12_1_0) ^ port_state_in_15_1_0);
  assign state_out_14_1_0 = (((mul2_118_port_byte_out_0 ^ mul3_118_port_byte_out_0) ^ port_state_in_12_1_0) ^ port_state_in_13_1_0);
  assign state_out_15_1_0 = (((mul2_119_port_byte_out_0 ^ mul3_119_port_byte_out_0) ^ port_state_in_13_1_0) ^ port_state_in_14_1_0);
  assign state_out_12_1_1 = (((mul2_116_port_byte_out_1 ^ mul3_116_port_byte_out_1) ^ port_state_in_14_1_1) ^ port_state_in_15_1_1);
  assign state_out_13_1_1 = (((mul2_117_port_byte_out_1 ^ mul3_117_port_byte_out_1) ^ port_state_in_12_1_1) ^ port_state_in_15_1_1);
  assign state_out_14_1_1 = (((mul2_118_port_byte_out_1 ^ mul3_118_port_byte_out_1) ^ port_state_in_12_1_1) ^ port_state_in_13_1_1);
  assign state_out_15_1_1 = (((mul2_119_port_byte_out_1 ^ mul3_119_port_byte_out_1) ^ port_state_in_13_1_1) ^ port_state_in_14_1_1);
  assign state_out_12_1_2 = (((mul2_116_port_byte_out_2 ^ mul3_116_port_byte_out_2) ^ port_state_in_14_1_2) ^ port_state_in_15_1_2);
  assign state_out_13_1_2 = (((mul2_117_port_byte_out_2 ^ mul3_117_port_byte_out_2) ^ port_state_in_12_1_2) ^ port_state_in_15_1_2);
  assign state_out_14_1_2 = (((mul2_118_port_byte_out_2 ^ mul3_118_port_byte_out_2) ^ port_state_in_12_1_2) ^ port_state_in_13_1_2);
  assign state_out_15_1_2 = (((mul2_119_port_byte_out_2 ^ mul3_119_port_byte_out_2) ^ port_state_in_13_1_2) ^ port_state_in_14_1_2);
  assign state_out_12_1_3 = (((mul2_116_port_byte_out_3 ^ mul3_116_port_byte_out_3) ^ port_state_in_14_1_3) ^ port_state_in_15_1_3);
  assign state_out_13_1_3 = (((mul2_117_port_byte_out_3 ^ mul3_117_port_byte_out_3) ^ port_state_in_12_1_3) ^ port_state_in_15_1_3);
  assign state_out_14_1_3 = (((mul2_118_port_byte_out_3 ^ mul3_118_port_byte_out_3) ^ port_state_in_12_1_3) ^ port_state_in_13_1_3);
  assign state_out_15_1_3 = (((mul2_119_port_byte_out_3 ^ mul3_119_port_byte_out_3) ^ port_state_in_13_1_3) ^ port_state_in_14_1_3);
  assign state_out_12_1_4 = (((mul2_116_port_byte_out_4 ^ mul3_116_port_byte_out_4) ^ port_state_in_14_1_4) ^ port_state_in_15_1_4);
  assign state_out_13_1_4 = (((mul2_117_port_byte_out_4 ^ mul3_117_port_byte_out_4) ^ port_state_in_12_1_4) ^ port_state_in_15_1_4);
  assign state_out_14_1_4 = (((mul2_118_port_byte_out_4 ^ mul3_118_port_byte_out_4) ^ port_state_in_12_1_4) ^ port_state_in_13_1_4);
  assign state_out_15_1_4 = (((mul2_119_port_byte_out_4 ^ mul3_119_port_byte_out_4) ^ port_state_in_13_1_4) ^ port_state_in_14_1_4);
  assign state_out_12_1_5 = (((mul2_116_port_byte_out_5 ^ mul3_116_port_byte_out_5) ^ port_state_in_14_1_5) ^ port_state_in_15_1_5);
  assign state_out_13_1_5 = (((mul2_117_port_byte_out_5 ^ mul3_117_port_byte_out_5) ^ port_state_in_12_1_5) ^ port_state_in_15_1_5);
  assign state_out_14_1_5 = (((mul2_118_port_byte_out_5 ^ mul3_118_port_byte_out_5) ^ port_state_in_12_1_5) ^ port_state_in_13_1_5);
  assign state_out_15_1_5 = (((mul2_119_port_byte_out_5 ^ mul3_119_port_byte_out_5) ^ port_state_in_13_1_5) ^ port_state_in_14_1_5);
  assign state_out_12_1_6 = (((mul2_116_port_byte_out_6 ^ mul3_116_port_byte_out_6) ^ port_state_in_14_1_6) ^ port_state_in_15_1_6);
  assign state_out_13_1_6 = (((mul2_117_port_byte_out_6 ^ mul3_117_port_byte_out_6) ^ port_state_in_12_1_6) ^ port_state_in_15_1_6);
  assign state_out_14_1_6 = (((mul2_118_port_byte_out_6 ^ mul3_118_port_byte_out_6) ^ port_state_in_12_1_6) ^ port_state_in_13_1_6);
  assign state_out_15_1_6 = (((mul2_119_port_byte_out_6 ^ mul3_119_port_byte_out_6) ^ port_state_in_13_1_6) ^ port_state_in_14_1_6);
  assign state_out_12_1_7 = (((mul2_116_port_byte_out_7 ^ mul3_116_port_byte_out_7) ^ port_state_in_14_1_7) ^ port_state_in_15_1_7);
  assign state_out_13_1_7 = (((mul2_117_port_byte_out_7 ^ mul3_117_port_byte_out_7) ^ port_state_in_12_1_7) ^ port_state_in_15_1_7);
  assign state_out_14_1_7 = (((mul2_118_port_byte_out_7 ^ mul3_118_port_byte_out_7) ^ port_state_in_12_1_7) ^ port_state_in_13_1_7);
  assign state_out_15_1_7 = (((mul2_119_port_byte_out_7 ^ mul3_119_port_byte_out_7) ^ port_state_in_13_1_7) ^ port_state_in_14_1_7);
  assign state_out_12_2_0 = (((mul2_120_port_byte_out_0 ^ mul3_120_port_byte_out_0) ^ port_state_in_14_2_0) ^ port_state_in_15_2_0);
  assign state_out_13_2_0 = (((mul2_121_port_byte_out_0 ^ mul3_121_port_byte_out_0) ^ port_state_in_12_2_0) ^ port_state_in_15_2_0);
  assign state_out_14_2_0 = (((mul2_122_port_byte_out_0 ^ mul3_122_port_byte_out_0) ^ port_state_in_12_2_0) ^ port_state_in_13_2_0);
  assign state_out_15_2_0 = (((mul2_123_port_byte_out_0 ^ mul3_123_port_byte_out_0) ^ port_state_in_13_2_0) ^ port_state_in_14_2_0);
  assign state_out_12_2_1 = (((mul2_120_port_byte_out_1 ^ mul3_120_port_byte_out_1) ^ port_state_in_14_2_1) ^ port_state_in_15_2_1);
  assign state_out_13_2_1 = (((mul2_121_port_byte_out_1 ^ mul3_121_port_byte_out_1) ^ port_state_in_12_2_1) ^ port_state_in_15_2_1);
  assign state_out_14_2_1 = (((mul2_122_port_byte_out_1 ^ mul3_122_port_byte_out_1) ^ port_state_in_12_2_1) ^ port_state_in_13_2_1);
  assign state_out_15_2_1 = (((mul2_123_port_byte_out_1 ^ mul3_123_port_byte_out_1) ^ port_state_in_13_2_1) ^ port_state_in_14_2_1);
  assign state_out_12_2_2 = (((mul2_120_port_byte_out_2 ^ mul3_120_port_byte_out_2) ^ port_state_in_14_2_2) ^ port_state_in_15_2_2);
  assign state_out_13_2_2 = (((mul2_121_port_byte_out_2 ^ mul3_121_port_byte_out_2) ^ port_state_in_12_2_2) ^ port_state_in_15_2_2);
  assign state_out_14_2_2 = (((mul2_122_port_byte_out_2 ^ mul3_122_port_byte_out_2) ^ port_state_in_12_2_2) ^ port_state_in_13_2_2);
  assign state_out_15_2_2 = (((mul2_123_port_byte_out_2 ^ mul3_123_port_byte_out_2) ^ port_state_in_13_2_2) ^ port_state_in_14_2_2);
  assign state_out_12_2_3 = (((mul2_120_port_byte_out_3 ^ mul3_120_port_byte_out_3) ^ port_state_in_14_2_3) ^ port_state_in_15_2_3);
  assign state_out_13_2_3 = (((mul2_121_port_byte_out_3 ^ mul3_121_port_byte_out_3) ^ port_state_in_12_2_3) ^ port_state_in_15_2_3);
  assign state_out_14_2_3 = (((mul2_122_port_byte_out_3 ^ mul3_122_port_byte_out_3) ^ port_state_in_12_2_3) ^ port_state_in_13_2_3);
  assign state_out_15_2_3 = (((mul2_123_port_byte_out_3 ^ mul3_123_port_byte_out_3) ^ port_state_in_13_2_3) ^ port_state_in_14_2_3);
  assign state_out_12_2_4 = (((mul2_120_port_byte_out_4 ^ mul3_120_port_byte_out_4) ^ port_state_in_14_2_4) ^ port_state_in_15_2_4);
  assign state_out_13_2_4 = (((mul2_121_port_byte_out_4 ^ mul3_121_port_byte_out_4) ^ port_state_in_12_2_4) ^ port_state_in_15_2_4);
  assign state_out_14_2_4 = (((mul2_122_port_byte_out_4 ^ mul3_122_port_byte_out_4) ^ port_state_in_12_2_4) ^ port_state_in_13_2_4);
  assign state_out_15_2_4 = (((mul2_123_port_byte_out_4 ^ mul3_123_port_byte_out_4) ^ port_state_in_13_2_4) ^ port_state_in_14_2_4);
  assign state_out_12_2_5 = (((mul2_120_port_byte_out_5 ^ mul3_120_port_byte_out_5) ^ port_state_in_14_2_5) ^ port_state_in_15_2_5);
  assign state_out_13_2_5 = (((mul2_121_port_byte_out_5 ^ mul3_121_port_byte_out_5) ^ port_state_in_12_2_5) ^ port_state_in_15_2_5);
  assign state_out_14_2_5 = (((mul2_122_port_byte_out_5 ^ mul3_122_port_byte_out_5) ^ port_state_in_12_2_5) ^ port_state_in_13_2_5);
  assign state_out_15_2_5 = (((mul2_123_port_byte_out_5 ^ mul3_123_port_byte_out_5) ^ port_state_in_13_2_5) ^ port_state_in_14_2_5);
  assign state_out_12_2_6 = (((mul2_120_port_byte_out_6 ^ mul3_120_port_byte_out_6) ^ port_state_in_14_2_6) ^ port_state_in_15_2_6);
  assign state_out_13_2_6 = (((mul2_121_port_byte_out_6 ^ mul3_121_port_byte_out_6) ^ port_state_in_12_2_6) ^ port_state_in_15_2_6);
  assign state_out_14_2_6 = (((mul2_122_port_byte_out_6 ^ mul3_122_port_byte_out_6) ^ port_state_in_12_2_6) ^ port_state_in_13_2_6);
  assign state_out_15_2_6 = (((mul2_123_port_byte_out_6 ^ mul3_123_port_byte_out_6) ^ port_state_in_13_2_6) ^ port_state_in_14_2_6);
  assign state_out_12_2_7 = (((mul2_120_port_byte_out_7 ^ mul3_120_port_byte_out_7) ^ port_state_in_14_2_7) ^ port_state_in_15_2_7);
  assign state_out_13_2_7 = (((mul2_121_port_byte_out_7 ^ mul3_121_port_byte_out_7) ^ port_state_in_12_2_7) ^ port_state_in_15_2_7);
  assign state_out_14_2_7 = (((mul2_122_port_byte_out_7 ^ mul3_122_port_byte_out_7) ^ port_state_in_12_2_7) ^ port_state_in_13_2_7);
  assign state_out_15_2_7 = (((mul2_123_port_byte_out_7 ^ mul3_123_port_byte_out_7) ^ port_state_in_13_2_7) ^ port_state_in_14_2_7);
  assign state_out_12_3_0 = (((mul2_124_port_byte_out_0 ^ mul3_124_port_byte_out_0) ^ port_state_in_14_3_0) ^ port_state_in_15_3_0);
  assign state_out_13_3_0 = (((mul2_125_port_byte_out_0 ^ mul3_125_port_byte_out_0) ^ port_state_in_12_3_0) ^ port_state_in_15_3_0);
  assign state_out_14_3_0 = (((mul2_126_port_byte_out_0 ^ mul3_126_port_byte_out_0) ^ port_state_in_12_3_0) ^ port_state_in_13_3_0);
  assign state_out_15_3_0 = (((mul2_127_port_byte_out_0 ^ mul3_127_port_byte_out_0) ^ port_state_in_13_3_0) ^ port_state_in_14_3_0);
  assign state_out_12_3_1 = (((mul2_124_port_byte_out_1 ^ mul3_124_port_byte_out_1) ^ port_state_in_14_3_1) ^ port_state_in_15_3_1);
  assign state_out_13_3_1 = (((mul2_125_port_byte_out_1 ^ mul3_125_port_byte_out_1) ^ port_state_in_12_3_1) ^ port_state_in_15_3_1);
  assign state_out_14_3_1 = (((mul2_126_port_byte_out_1 ^ mul3_126_port_byte_out_1) ^ port_state_in_12_3_1) ^ port_state_in_13_3_1);
  assign state_out_15_3_1 = (((mul2_127_port_byte_out_1 ^ mul3_127_port_byte_out_1) ^ port_state_in_13_3_1) ^ port_state_in_14_3_1);
  assign state_out_12_3_2 = (((mul2_124_port_byte_out_2 ^ mul3_124_port_byte_out_2) ^ port_state_in_14_3_2) ^ port_state_in_15_3_2);
  assign state_out_13_3_2 = (((mul2_125_port_byte_out_2 ^ mul3_125_port_byte_out_2) ^ port_state_in_12_3_2) ^ port_state_in_15_3_2);
  assign state_out_14_3_2 = (((mul2_126_port_byte_out_2 ^ mul3_126_port_byte_out_2) ^ port_state_in_12_3_2) ^ port_state_in_13_3_2);
  assign state_out_15_3_2 = (((mul2_127_port_byte_out_2 ^ mul3_127_port_byte_out_2) ^ port_state_in_13_3_2) ^ port_state_in_14_3_2);
  assign state_out_12_3_3 = (((mul2_124_port_byte_out_3 ^ mul3_124_port_byte_out_3) ^ port_state_in_14_3_3) ^ port_state_in_15_3_3);
  assign state_out_13_3_3 = (((mul2_125_port_byte_out_3 ^ mul3_125_port_byte_out_3) ^ port_state_in_12_3_3) ^ port_state_in_15_3_3);
  assign state_out_14_3_3 = (((mul2_126_port_byte_out_3 ^ mul3_126_port_byte_out_3) ^ port_state_in_12_3_3) ^ port_state_in_13_3_3);
  assign state_out_15_3_3 = (((mul2_127_port_byte_out_3 ^ mul3_127_port_byte_out_3) ^ port_state_in_13_3_3) ^ port_state_in_14_3_3);
  assign state_out_12_3_4 = (((mul2_124_port_byte_out_4 ^ mul3_124_port_byte_out_4) ^ port_state_in_14_3_4) ^ port_state_in_15_3_4);
  assign state_out_13_3_4 = (((mul2_125_port_byte_out_4 ^ mul3_125_port_byte_out_4) ^ port_state_in_12_3_4) ^ port_state_in_15_3_4);
  assign state_out_14_3_4 = (((mul2_126_port_byte_out_4 ^ mul3_126_port_byte_out_4) ^ port_state_in_12_3_4) ^ port_state_in_13_3_4);
  assign state_out_15_3_4 = (((mul2_127_port_byte_out_4 ^ mul3_127_port_byte_out_4) ^ port_state_in_13_3_4) ^ port_state_in_14_3_4);
  assign state_out_12_3_5 = (((mul2_124_port_byte_out_5 ^ mul3_124_port_byte_out_5) ^ port_state_in_14_3_5) ^ port_state_in_15_3_5);
  assign state_out_13_3_5 = (((mul2_125_port_byte_out_5 ^ mul3_125_port_byte_out_5) ^ port_state_in_12_3_5) ^ port_state_in_15_3_5);
  assign state_out_14_3_5 = (((mul2_126_port_byte_out_5 ^ mul3_126_port_byte_out_5) ^ port_state_in_12_3_5) ^ port_state_in_13_3_5);
  assign state_out_15_3_5 = (((mul2_127_port_byte_out_5 ^ mul3_127_port_byte_out_5) ^ port_state_in_13_3_5) ^ port_state_in_14_3_5);
  assign state_out_12_3_6 = (((mul2_124_port_byte_out_6 ^ mul3_124_port_byte_out_6) ^ port_state_in_14_3_6) ^ port_state_in_15_3_6);
  assign state_out_13_3_6 = (((mul2_125_port_byte_out_6 ^ mul3_125_port_byte_out_6) ^ port_state_in_12_3_6) ^ port_state_in_15_3_6);
  assign state_out_14_3_6 = (((mul2_126_port_byte_out_6 ^ mul3_126_port_byte_out_6) ^ port_state_in_12_3_6) ^ port_state_in_13_3_6);
  assign state_out_15_3_6 = (((mul2_127_port_byte_out_6 ^ mul3_127_port_byte_out_6) ^ port_state_in_13_3_6) ^ port_state_in_14_3_6);
  assign state_out_12_3_7 = (((mul2_124_port_byte_out_7 ^ mul3_124_port_byte_out_7) ^ port_state_in_14_3_7) ^ port_state_in_15_3_7);
  assign state_out_13_3_7 = (((mul2_125_port_byte_out_7 ^ mul3_125_port_byte_out_7) ^ port_state_in_12_3_7) ^ port_state_in_15_3_7);
  assign state_out_14_3_7 = (((mul2_126_port_byte_out_7 ^ mul3_126_port_byte_out_7) ^ port_state_in_12_3_7) ^ port_state_in_13_3_7);
  assign state_out_15_3_7 = (((mul2_127_port_byte_out_7 ^ mul3_127_port_byte_out_7) ^ port_state_in_13_3_7) ^ port_state_in_14_3_7);
  assign port_state_out_0_0_0 = state_out_0_0_0;
  assign port_state_out_0_0_1 = state_out_0_0_1;
  assign port_state_out_0_0_2 = state_out_0_0_2;
  assign port_state_out_0_0_3 = state_out_0_0_3;
  assign port_state_out_0_0_4 = state_out_0_0_4;
  assign port_state_out_0_0_5 = state_out_0_0_5;
  assign port_state_out_0_0_6 = state_out_0_0_6;
  assign port_state_out_0_0_7 = state_out_0_0_7;
  assign port_state_out_0_1_0 = state_out_0_1_0;
  assign port_state_out_0_1_1 = state_out_0_1_1;
  assign port_state_out_0_1_2 = state_out_0_1_2;
  assign port_state_out_0_1_3 = state_out_0_1_3;
  assign port_state_out_0_1_4 = state_out_0_1_4;
  assign port_state_out_0_1_5 = state_out_0_1_5;
  assign port_state_out_0_1_6 = state_out_0_1_6;
  assign port_state_out_0_1_7 = state_out_0_1_7;
  assign port_state_out_0_2_0 = state_out_0_2_0;
  assign port_state_out_0_2_1 = state_out_0_2_1;
  assign port_state_out_0_2_2 = state_out_0_2_2;
  assign port_state_out_0_2_3 = state_out_0_2_3;
  assign port_state_out_0_2_4 = state_out_0_2_4;
  assign port_state_out_0_2_5 = state_out_0_2_5;
  assign port_state_out_0_2_6 = state_out_0_2_6;
  assign port_state_out_0_2_7 = state_out_0_2_7;
  assign port_state_out_0_3_0 = state_out_0_3_0;
  assign port_state_out_0_3_1 = state_out_0_3_1;
  assign port_state_out_0_3_2 = state_out_0_3_2;
  assign port_state_out_0_3_3 = state_out_0_3_3;
  assign port_state_out_0_3_4 = state_out_0_3_4;
  assign port_state_out_0_3_5 = state_out_0_3_5;
  assign port_state_out_0_3_6 = state_out_0_3_6;
  assign port_state_out_0_3_7 = state_out_0_3_7;
  assign port_state_out_1_0_0 = state_out_1_0_0;
  assign port_state_out_1_0_1 = state_out_1_0_1;
  assign port_state_out_1_0_2 = state_out_1_0_2;
  assign port_state_out_1_0_3 = state_out_1_0_3;
  assign port_state_out_1_0_4 = state_out_1_0_4;
  assign port_state_out_1_0_5 = state_out_1_0_5;
  assign port_state_out_1_0_6 = state_out_1_0_6;
  assign port_state_out_1_0_7 = state_out_1_0_7;
  assign port_state_out_1_1_0 = state_out_1_1_0;
  assign port_state_out_1_1_1 = state_out_1_1_1;
  assign port_state_out_1_1_2 = state_out_1_1_2;
  assign port_state_out_1_1_3 = state_out_1_1_3;
  assign port_state_out_1_1_4 = state_out_1_1_4;
  assign port_state_out_1_1_5 = state_out_1_1_5;
  assign port_state_out_1_1_6 = state_out_1_1_6;
  assign port_state_out_1_1_7 = state_out_1_1_7;
  assign port_state_out_1_2_0 = state_out_1_2_0;
  assign port_state_out_1_2_1 = state_out_1_2_1;
  assign port_state_out_1_2_2 = state_out_1_2_2;
  assign port_state_out_1_2_3 = state_out_1_2_3;
  assign port_state_out_1_2_4 = state_out_1_2_4;
  assign port_state_out_1_2_5 = state_out_1_2_5;
  assign port_state_out_1_2_6 = state_out_1_2_6;
  assign port_state_out_1_2_7 = state_out_1_2_7;
  assign port_state_out_1_3_0 = state_out_1_3_0;
  assign port_state_out_1_3_1 = state_out_1_3_1;
  assign port_state_out_1_3_2 = state_out_1_3_2;
  assign port_state_out_1_3_3 = state_out_1_3_3;
  assign port_state_out_1_3_4 = state_out_1_3_4;
  assign port_state_out_1_3_5 = state_out_1_3_5;
  assign port_state_out_1_3_6 = state_out_1_3_6;
  assign port_state_out_1_3_7 = state_out_1_3_7;
  assign port_state_out_2_0_0 = state_out_2_0_0;
  assign port_state_out_2_0_1 = state_out_2_0_1;
  assign port_state_out_2_0_2 = state_out_2_0_2;
  assign port_state_out_2_0_3 = state_out_2_0_3;
  assign port_state_out_2_0_4 = state_out_2_0_4;
  assign port_state_out_2_0_5 = state_out_2_0_5;
  assign port_state_out_2_0_6 = state_out_2_0_6;
  assign port_state_out_2_0_7 = state_out_2_0_7;
  assign port_state_out_2_1_0 = state_out_2_1_0;
  assign port_state_out_2_1_1 = state_out_2_1_1;
  assign port_state_out_2_1_2 = state_out_2_1_2;
  assign port_state_out_2_1_3 = state_out_2_1_3;
  assign port_state_out_2_1_4 = state_out_2_1_4;
  assign port_state_out_2_1_5 = state_out_2_1_5;
  assign port_state_out_2_1_6 = state_out_2_1_6;
  assign port_state_out_2_1_7 = state_out_2_1_7;
  assign port_state_out_2_2_0 = state_out_2_2_0;
  assign port_state_out_2_2_1 = state_out_2_2_1;
  assign port_state_out_2_2_2 = state_out_2_2_2;
  assign port_state_out_2_2_3 = state_out_2_2_3;
  assign port_state_out_2_2_4 = state_out_2_2_4;
  assign port_state_out_2_2_5 = state_out_2_2_5;
  assign port_state_out_2_2_6 = state_out_2_2_6;
  assign port_state_out_2_2_7 = state_out_2_2_7;
  assign port_state_out_2_3_0 = state_out_2_3_0;
  assign port_state_out_2_3_1 = state_out_2_3_1;
  assign port_state_out_2_3_2 = state_out_2_3_2;
  assign port_state_out_2_3_3 = state_out_2_3_3;
  assign port_state_out_2_3_4 = state_out_2_3_4;
  assign port_state_out_2_3_5 = state_out_2_3_5;
  assign port_state_out_2_3_6 = state_out_2_3_6;
  assign port_state_out_2_3_7 = state_out_2_3_7;
  assign port_state_out_3_0_0 = state_out_3_0_0;
  assign port_state_out_3_0_1 = state_out_3_0_1;
  assign port_state_out_3_0_2 = state_out_3_0_2;
  assign port_state_out_3_0_3 = state_out_3_0_3;
  assign port_state_out_3_0_4 = state_out_3_0_4;
  assign port_state_out_3_0_5 = state_out_3_0_5;
  assign port_state_out_3_0_6 = state_out_3_0_6;
  assign port_state_out_3_0_7 = state_out_3_0_7;
  assign port_state_out_3_1_0 = state_out_3_1_0;
  assign port_state_out_3_1_1 = state_out_3_1_1;
  assign port_state_out_3_1_2 = state_out_3_1_2;
  assign port_state_out_3_1_3 = state_out_3_1_3;
  assign port_state_out_3_1_4 = state_out_3_1_4;
  assign port_state_out_3_1_5 = state_out_3_1_5;
  assign port_state_out_3_1_6 = state_out_3_1_6;
  assign port_state_out_3_1_7 = state_out_3_1_7;
  assign port_state_out_3_2_0 = state_out_3_2_0;
  assign port_state_out_3_2_1 = state_out_3_2_1;
  assign port_state_out_3_2_2 = state_out_3_2_2;
  assign port_state_out_3_2_3 = state_out_3_2_3;
  assign port_state_out_3_2_4 = state_out_3_2_4;
  assign port_state_out_3_2_5 = state_out_3_2_5;
  assign port_state_out_3_2_6 = state_out_3_2_6;
  assign port_state_out_3_2_7 = state_out_3_2_7;
  assign port_state_out_3_3_0 = state_out_3_3_0;
  assign port_state_out_3_3_1 = state_out_3_3_1;
  assign port_state_out_3_3_2 = state_out_3_3_2;
  assign port_state_out_3_3_3 = state_out_3_3_3;
  assign port_state_out_3_3_4 = state_out_3_3_4;
  assign port_state_out_3_3_5 = state_out_3_3_5;
  assign port_state_out_3_3_6 = state_out_3_3_6;
  assign port_state_out_3_3_7 = state_out_3_3_7;
  assign port_state_out_4_0_0 = state_out_4_0_0;
  assign port_state_out_4_0_1 = state_out_4_0_1;
  assign port_state_out_4_0_2 = state_out_4_0_2;
  assign port_state_out_4_0_3 = state_out_4_0_3;
  assign port_state_out_4_0_4 = state_out_4_0_4;
  assign port_state_out_4_0_5 = state_out_4_0_5;
  assign port_state_out_4_0_6 = state_out_4_0_6;
  assign port_state_out_4_0_7 = state_out_4_0_7;
  assign port_state_out_4_1_0 = state_out_4_1_0;
  assign port_state_out_4_1_1 = state_out_4_1_1;
  assign port_state_out_4_1_2 = state_out_4_1_2;
  assign port_state_out_4_1_3 = state_out_4_1_3;
  assign port_state_out_4_1_4 = state_out_4_1_4;
  assign port_state_out_4_1_5 = state_out_4_1_5;
  assign port_state_out_4_1_6 = state_out_4_1_6;
  assign port_state_out_4_1_7 = state_out_4_1_7;
  assign port_state_out_4_2_0 = state_out_4_2_0;
  assign port_state_out_4_2_1 = state_out_4_2_1;
  assign port_state_out_4_2_2 = state_out_4_2_2;
  assign port_state_out_4_2_3 = state_out_4_2_3;
  assign port_state_out_4_2_4 = state_out_4_2_4;
  assign port_state_out_4_2_5 = state_out_4_2_5;
  assign port_state_out_4_2_6 = state_out_4_2_6;
  assign port_state_out_4_2_7 = state_out_4_2_7;
  assign port_state_out_4_3_0 = state_out_4_3_0;
  assign port_state_out_4_3_1 = state_out_4_3_1;
  assign port_state_out_4_3_2 = state_out_4_3_2;
  assign port_state_out_4_3_3 = state_out_4_3_3;
  assign port_state_out_4_3_4 = state_out_4_3_4;
  assign port_state_out_4_3_5 = state_out_4_3_5;
  assign port_state_out_4_3_6 = state_out_4_3_6;
  assign port_state_out_4_3_7 = state_out_4_3_7;
  assign port_state_out_5_0_0 = state_out_5_0_0;
  assign port_state_out_5_0_1 = state_out_5_0_1;
  assign port_state_out_5_0_2 = state_out_5_0_2;
  assign port_state_out_5_0_3 = state_out_5_0_3;
  assign port_state_out_5_0_4 = state_out_5_0_4;
  assign port_state_out_5_0_5 = state_out_5_0_5;
  assign port_state_out_5_0_6 = state_out_5_0_6;
  assign port_state_out_5_0_7 = state_out_5_0_7;
  assign port_state_out_5_1_0 = state_out_5_1_0;
  assign port_state_out_5_1_1 = state_out_5_1_1;
  assign port_state_out_5_1_2 = state_out_5_1_2;
  assign port_state_out_5_1_3 = state_out_5_1_3;
  assign port_state_out_5_1_4 = state_out_5_1_4;
  assign port_state_out_5_1_5 = state_out_5_1_5;
  assign port_state_out_5_1_6 = state_out_5_1_6;
  assign port_state_out_5_1_7 = state_out_5_1_7;
  assign port_state_out_5_2_0 = state_out_5_2_0;
  assign port_state_out_5_2_1 = state_out_5_2_1;
  assign port_state_out_5_2_2 = state_out_5_2_2;
  assign port_state_out_5_2_3 = state_out_5_2_3;
  assign port_state_out_5_2_4 = state_out_5_2_4;
  assign port_state_out_5_2_5 = state_out_5_2_5;
  assign port_state_out_5_2_6 = state_out_5_2_6;
  assign port_state_out_5_2_7 = state_out_5_2_7;
  assign port_state_out_5_3_0 = state_out_5_3_0;
  assign port_state_out_5_3_1 = state_out_5_3_1;
  assign port_state_out_5_3_2 = state_out_5_3_2;
  assign port_state_out_5_3_3 = state_out_5_3_3;
  assign port_state_out_5_3_4 = state_out_5_3_4;
  assign port_state_out_5_3_5 = state_out_5_3_5;
  assign port_state_out_5_3_6 = state_out_5_3_6;
  assign port_state_out_5_3_7 = state_out_5_3_7;
  assign port_state_out_6_0_0 = state_out_6_0_0;
  assign port_state_out_6_0_1 = state_out_6_0_1;
  assign port_state_out_6_0_2 = state_out_6_0_2;
  assign port_state_out_6_0_3 = state_out_6_0_3;
  assign port_state_out_6_0_4 = state_out_6_0_4;
  assign port_state_out_6_0_5 = state_out_6_0_5;
  assign port_state_out_6_0_6 = state_out_6_0_6;
  assign port_state_out_6_0_7 = state_out_6_0_7;
  assign port_state_out_6_1_0 = state_out_6_1_0;
  assign port_state_out_6_1_1 = state_out_6_1_1;
  assign port_state_out_6_1_2 = state_out_6_1_2;
  assign port_state_out_6_1_3 = state_out_6_1_3;
  assign port_state_out_6_1_4 = state_out_6_1_4;
  assign port_state_out_6_1_5 = state_out_6_1_5;
  assign port_state_out_6_1_6 = state_out_6_1_6;
  assign port_state_out_6_1_7 = state_out_6_1_7;
  assign port_state_out_6_2_0 = state_out_6_2_0;
  assign port_state_out_6_2_1 = state_out_6_2_1;
  assign port_state_out_6_2_2 = state_out_6_2_2;
  assign port_state_out_6_2_3 = state_out_6_2_3;
  assign port_state_out_6_2_4 = state_out_6_2_4;
  assign port_state_out_6_2_5 = state_out_6_2_5;
  assign port_state_out_6_2_6 = state_out_6_2_6;
  assign port_state_out_6_2_7 = state_out_6_2_7;
  assign port_state_out_6_3_0 = state_out_6_3_0;
  assign port_state_out_6_3_1 = state_out_6_3_1;
  assign port_state_out_6_3_2 = state_out_6_3_2;
  assign port_state_out_6_3_3 = state_out_6_3_3;
  assign port_state_out_6_3_4 = state_out_6_3_4;
  assign port_state_out_6_3_5 = state_out_6_3_5;
  assign port_state_out_6_3_6 = state_out_6_3_6;
  assign port_state_out_6_3_7 = state_out_6_3_7;
  assign port_state_out_7_0_0 = state_out_7_0_0;
  assign port_state_out_7_0_1 = state_out_7_0_1;
  assign port_state_out_7_0_2 = state_out_7_0_2;
  assign port_state_out_7_0_3 = state_out_7_0_3;
  assign port_state_out_7_0_4 = state_out_7_0_4;
  assign port_state_out_7_0_5 = state_out_7_0_5;
  assign port_state_out_7_0_6 = state_out_7_0_6;
  assign port_state_out_7_0_7 = state_out_7_0_7;
  assign port_state_out_7_1_0 = state_out_7_1_0;
  assign port_state_out_7_1_1 = state_out_7_1_1;
  assign port_state_out_7_1_2 = state_out_7_1_2;
  assign port_state_out_7_1_3 = state_out_7_1_3;
  assign port_state_out_7_1_4 = state_out_7_1_4;
  assign port_state_out_7_1_5 = state_out_7_1_5;
  assign port_state_out_7_1_6 = state_out_7_1_6;
  assign port_state_out_7_1_7 = state_out_7_1_7;
  assign port_state_out_7_2_0 = state_out_7_2_0;
  assign port_state_out_7_2_1 = state_out_7_2_1;
  assign port_state_out_7_2_2 = state_out_7_2_2;
  assign port_state_out_7_2_3 = state_out_7_2_3;
  assign port_state_out_7_2_4 = state_out_7_2_4;
  assign port_state_out_7_2_5 = state_out_7_2_5;
  assign port_state_out_7_2_6 = state_out_7_2_6;
  assign port_state_out_7_2_7 = state_out_7_2_7;
  assign port_state_out_7_3_0 = state_out_7_3_0;
  assign port_state_out_7_3_1 = state_out_7_3_1;
  assign port_state_out_7_3_2 = state_out_7_3_2;
  assign port_state_out_7_3_3 = state_out_7_3_3;
  assign port_state_out_7_3_4 = state_out_7_3_4;
  assign port_state_out_7_3_5 = state_out_7_3_5;
  assign port_state_out_7_3_6 = state_out_7_3_6;
  assign port_state_out_7_3_7 = state_out_7_3_7;
  assign port_state_out_8_0_0 = state_out_8_0_0;
  assign port_state_out_8_0_1 = state_out_8_0_1;
  assign port_state_out_8_0_2 = state_out_8_0_2;
  assign port_state_out_8_0_3 = state_out_8_0_3;
  assign port_state_out_8_0_4 = state_out_8_0_4;
  assign port_state_out_8_0_5 = state_out_8_0_5;
  assign port_state_out_8_0_6 = state_out_8_0_6;
  assign port_state_out_8_0_7 = state_out_8_0_7;
  assign port_state_out_8_1_0 = state_out_8_1_0;
  assign port_state_out_8_1_1 = state_out_8_1_1;
  assign port_state_out_8_1_2 = state_out_8_1_2;
  assign port_state_out_8_1_3 = state_out_8_1_3;
  assign port_state_out_8_1_4 = state_out_8_1_4;
  assign port_state_out_8_1_5 = state_out_8_1_5;
  assign port_state_out_8_1_6 = state_out_8_1_6;
  assign port_state_out_8_1_7 = state_out_8_1_7;
  assign port_state_out_8_2_0 = state_out_8_2_0;
  assign port_state_out_8_2_1 = state_out_8_2_1;
  assign port_state_out_8_2_2 = state_out_8_2_2;
  assign port_state_out_8_2_3 = state_out_8_2_3;
  assign port_state_out_8_2_4 = state_out_8_2_4;
  assign port_state_out_8_2_5 = state_out_8_2_5;
  assign port_state_out_8_2_6 = state_out_8_2_6;
  assign port_state_out_8_2_7 = state_out_8_2_7;
  assign port_state_out_8_3_0 = state_out_8_3_0;
  assign port_state_out_8_3_1 = state_out_8_3_1;
  assign port_state_out_8_3_2 = state_out_8_3_2;
  assign port_state_out_8_3_3 = state_out_8_3_3;
  assign port_state_out_8_3_4 = state_out_8_3_4;
  assign port_state_out_8_3_5 = state_out_8_3_5;
  assign port_state_out_8_3_6 = state_out_8_3_6;
  assign port_state_out_8_3_7 = state_out_8_3_7;
  assign port_state_out_9_0_0 = state_out_9_0_0;
  assign port_state_out_9_0_1 = state_out_9_0_1;
  assign port_state_out_9_0_2 = state_out_9_0_2;
  assign port_state_out_9_0_3 = state_out_9_0_3;
  assign port_state_out_9_0_4 = state_out_9_0_4;
  assign port_state_out_9_0_5 = state_out_9_0_5;
  assign port_state_out_9_0_6 = state_out_9_0_6;
  assign port_state_out_9_0_7 = state_out_9_0_7;
  assign port_state_out_9_1_0 = state_out_9_1_0;
  assign port_state_out_9_1_1 = state_out_9_1_1;
  assign port_state_out_9_1_2 = state_out_9_1_2;
  assign port_state_out_9_1_3 = state_out_9_1_3;
  assign port_state_out_9_1_4 = state_out_9_1_4;
  assign port_state_out_9_1_5 = state_out_9_1_5;
  assign port_state_out_9_1_6 = state_out_9_1_6;
  assign port_state_out_9_1_7 = state_out_9_1_7;
  assign port_state_out_9_2_0 = state_out_9_2_0;
  assign port_state_out_9_2_1 = state_out_9_2_1;
  assign port_state_out_9_2_2 = state_out_9_2_2;
  assign port_state_out_9_2_3 = state_out_9_2_3;
  assign port_state_out_9_2_4 = state_out_9_2_4;
  assign port_state_out_9_2_5 = state_out_9_2_5;
  assign port_state_out_9_2_6 = state_out_9_2_6;
  assign port_state_out_9_2_7 = state_out_9_2_7;
  assign port_state_out_9_3_0 = state_out_9_3_0;
  assign port_state_out_9_3_1 = state_out_9_3_1;
  assign port_state_out_9_3_2 = state_out_9_3_2;
  assign port_state_out_9_3_3 = state_out_9_3_3;
  assign port_state_out_9_3_4 = state_out_9_3_4;
  assign port_state_out_9_3_5 = state_out_9_3_5;
  assign port_state_out_9_3_6 = state_out_9_3_6;
  assign port_state_out_9_3_7 = state_out_9_3_7;
  assign port_state_out_10_0_0 = state_out_10_0_0;
  assign port_state_out_10_0_1 = state_out_10_0_1;
  assign port_state_out_10_0_2 = state_out_10_0_2;
  assign port_state_out_10_0_3 = state_out_10_0_3;
  assign port_state_out_10_0_4 = state_out_10_0_4;
  assign port_state_out_10_0_5 = state_out_10_0_5;
  assign port_state_out_10_0_6 = state_out_10_0_6;
  assign port_state_out_10_0_7 = state_out_10_0_7;
  assign port_state_out_10_1_0 = state_out_10_1_0;
  assign port_state_out_10_1_1 = state_out_10_1_1;
  assign port_state_out_10_1_2 = state_out_10_1_2;
  assign port_state_out_10_1_3 = state_out_10_1_3;
  assign port_state_out_10_1_4 = state_out_10_1_4;
  assign port_state_out_10_1_5 = state_out_10_1_5;
  assign port_state_out_10_1_6 = state_out_10_1_6;
  assign port_state_out_10_1_7 = state_out_10_1_7;
  assign port_state_out_10_2_0 = state_out_10_2_0;
  assign port_state_out_10_2_1 = state_out_10_2_1;
  assign port_state_out_10_2_2 = state_out_10_2_2;
  assign port_state_out_10_2_3 = state_out_10_2_3;
  assign port_state_out_10_2_4 = state_out_10_2_4;
  assign port_state_out_10_2_5 = state_out_10_2_5;
  assign port_state_out_10_2_6 = state_out_10_2_6;
  assign port_state_out_10_2_7 = state_out_10_2_7;
  assign port_state_out_10_3_0 = state_out_10_3_0;
  assign port_state_out_10_3_1 = state_out_10_3_1;
  assign port_state_out_10_3_2 = state_out_10_3_2;
  assign port_state_out_10_3_3 = state_out_10_3_3;
  assign port_state_out_10_3_4 = state_out_10_3_4;
  assign port_state_out_10_3_5 = state_out_10_3_5;
  assign port_state_out_10_3_6 = state_out_10_3_6;
  assign port_state_out_10_3_7 = state_out_10_3_7;
  assign port_state_out_11_0_0 = state_out_11_0_0;
  assign port_state_out_11_0_1 = state_out_11_0_1;
  assign port_state_out_11_0_2 = state_out_11_0_2;
  assign port_state_out_11_0_3 = state_out_11_0_3;
  assign port_state_out_11_0_4 = state_out_11_0_4;
  assign port_state_out_11_0_5 = state_out_11_0_5;
  assign port_state_out_11_0_6 = state_out_11_0_6;
  assign port_state_out_11_0_7 = state_out_11_0_7;
  assign port_state_out_11_1_0 = state_out_11_1_0;
  assign port_state_out_11_1_1 = state_out_11_1_1;
  assign port_state_out_11_1_2 = state_out_11_1_2;
  assign port_state_out_11_1_3 = state_out_11_1_3;
  assign port_state_out_11_1_4 = state_out_11_1_4;
  assign port_state_out_11_1_5 = state_out_11_1_5;
  assign port_state_out_11_1_6 = state_out_11_1_6;
  assign port_state_out_11_1_7 = state_out_11_1_7;
  assign port_state_out_11_2_0 = state_out_11_2_0;
  assign port_state_out_11_2_1 = state_out_11_2_1;
  assign port_state_out_11_2_2 = state_out_11_2_2;
  assign port_state_out_11_2_3 = state_out_11_2_3;
  assign port_state_out_11_2_4 = state_out_11_2_4;
  assign port_state_out_11_2_5 = state_out_11_2_5;
  assign port_state_out_11_2_6 = state_out_11_2_6;
  assign port_state_out_11_2_7 = state_out_11_2_7;
  assign port_state_out_11_3_0 = state_out_11_3_0;
  assign port_state_out_11_3_1 = state_out_11_3_1;
  assign port_state_out_11_3_2 = state_out_11_3_2;
  assign port_state_out_11_3_3 = state_out_11_3_3;
  assign port_state_out_11_3_4 = state_out_11_3_4;
  assign port_state_out_11_3_5 = state_out_11_3_5;
  assign port_state_out_11_3_6 = state_out_11_3_6;
  assign port_state_out_11_3_7 = state_out_11_3_7;
  assign port_state_out_12_0_0 = state_out_12_0_0;
  assign port_state_out_12_0_1 = state_out_12_0_1;
  assign port_state_out_12_0_2 = state_out_12_0_2;
  assign port_state_out_12_0_3 = state_out_12_0_3;
  assign port_state_out_12_0_4 = state_out_12_0_4;
  assign port_state_out_12_0_5 = state_out_12_0_5;
  assign port_state_out_12_0_6 = state_out_12_0_6;
  assign port_state_out_12_0_7 = state_out_12_0_7;
  assign port_state_out_12_1_0 = state_out_12_1_0;
  assign port_state_out_12_1_1 = state_out_12_1_1;
  assign port_state_out_12_1_2 = state_out_12_1_2;
  assign port_state_out_12_1_3 = state_out_12_1_3;
  assign port_state_out_12_1_4 = state_out_12_1_4;
  assign port_state_out_12_1_5 = state_out_12_1_5;
  assign port_state_out_12_1_6 = state_out_12_1_6;
  assign port_state_out_12_1_7 = state_out_12_1_7;
  assign port_state_out_12_2_0 = state_out_12_2_0;
  assign port_state_out_12_2_1 = state_out_12_2_1;
  assign port_state_out_12_2_2 = state_out_12_2_2;
  assign port_state_out_12_2_3 = state_out_12_2_3;
  assign port_state_out_12_2_4 = state_out_12_2_4;
  assign port_state_out_12_2_5 = state_out_12_2_5;
  assign port_state_out_12_2_6 = state_out_12_2_6;
  assign port_state_out_12_2_7 = state_out_12_2_7;
  assign port_state_out_12_3_0 = state_out_12_3_0;
  assign port_state_out_12_3_1 = state_out_12_3_1;
  assign port_state_out_12_3_2 = state_out_12_3_2;
  assign port_state_out_12_3_3 = state_out_12_3_3;
  assign port_state_out_12_3_4 = state_out_12_3_4;
  assign port_state_out_12_3_5 = state_out_12_3_5;
  assign port_state_out_12_3_6 = state_out_12_3_6;
  assign port_state_out_12_3_7 = state_out_12_3_7;
  assign port_state_out_13_0_0 = state_out_13_0_0;
  assign port_state_out_13_0_1 = state_out_13_0_1;
  assign port_state_out_13_0_2 = state_out_13_0_2;
  assign port_state_out_13_0_3 = state_out_13_0_3;
  assign port_state_out_13_0_4 = state_out_13_0_4;
  assign port_state_out_13_0_5 = state_out_13_0_5;
  assign port_state_out_13_0_6 = state_out_13_0_6;
  assign port_state_out_13_0_7 = state_out_13_0_7;
  assign port_state_out_13_1_0 = state_out_13_1_0;
  assign port_state_out_13_1_1 = state_out_13_1_1;
  assign port_state_out_13_1_2 = state_out_13_1_2;
  assign port_state_out_13_1_3 = state_out_13_1_3;
  assign port_state_out_13_1_4 = state_out_13_1_4;
  assign port_state_out_13_1_5 = state_out_13_1_5;
  assign port_state_out_13_1_6 = state_out_13_1_6;
  assign port_state_out_13_1_7 = state_out_13_1_7;
  assign port_state_out_13_2_0 = state_out_13_2_0;
  assign port_state_out_13_2_1 = state_out_13_2_1;
  assign port_state_out_13_2_2 = state_out_13_2_2;
  assign port_state_out_13_2_3 = state_out_13_2_3;
  assign port_state_out_13_2_4 = state_out_13_2_4;
  assign port_state_out_13_2_5 = state_out_13_2_5;
  assign port_state_out_13_2_6 = state_out_13_2_6;
  assign port_state_out_13_2_7 = state_out_13_2_7;
  assign port_state_out_13_3_0 = state_out_13_3_0;
  assign port_state_out_13_3_1 = state_out_13_3_1;
  assign port_state_out_13_3_2 = state_out_13_3_2;
  assign port_state_out_13_3_3 = state_out_13_3_3;
  assign port_state_out_13_3_4 = state_out_13_3_4;
  assign port_state_out_13_3_5 = state_out_13_3_5;
  assign port_state_out_13_3_6 = state_out_13_3_6;
  assign port_state_out_13_3_7 = state_out_13_3_7;
  assign port_state_out_14_0_0 = state_out_14_0_0;
  assign port_state_out_14_0_1 = state_out_14_0_1;
  assign port_state_out_14_0_2 = state_out_14_0_2;
  assign port_state_out_14_0_3 = state_out_14_0_3;
  assign port_state_out_14_0_4 = state_out_14_0_4;
  assign port_state_out_14_0_5 = state_out_14_0_5;
  assign port_state_out_14_0_6 = state_out_14_0_6;
  assign port_state_out_14_0_7 = state_out_14_0_7;
  assign port_state_out_14_1_0 = state_out_14_1_0;
  assign port_state_out_14_1_1 = state_out_14_1_1;
  assign port_state_out_14_1_2 = state_out_14_1_2;
  assign port_state_out_14_1_3 = state_out_14_1_3;
  assign port_state_out_14_1_4 = state_out_14_1_4;
  assign port_state_out_14_1_5 = state_out_14_1_5;
  assign port_state_out_14_1_6 = state_out_14_1_6;
  assign port_state_out_14_1_7 = state_out_14_1_7;
  assign port_state_out_14_2_0 = state_out_14_2_0;
  assign port_state_out_14_2_1 = state_out_14_2_1;
  assign port_state_out_14_2_2 = state_out_14_2_2;
  assign port_state_out_14_2_3 = state_out_14_2_3;
  assign port_state_out_14_2_4 = state_out_14_2_4;
  assign port_state_out_14_2_5 = state_out_14_2_5;
  assign port_state_out_14_2_6 = state_out_14_2_6;
  assign port_state_out_14_2_7 = state_out_14_2_7;
  assign port_state_out_14_3_0 = state_out_14_3_0;
  assign port_state_out_14_3_1 = state_out_14_3_1;
  assign port_state_out_14_3_2 = state_out_14_3_2;
  assign port_state_out_14_3_3 = state_out_14_3_3;
  assign port_state_out_14_3_4 = state_out_14_3_4;
  assign port_state_out_14_3_5 = state_out_14_3_5;
  assign port_state_out_14_3_6 = state_out_14_3_6;
  assign port_state_out_14_3_7 = state_out_14_3_7;
  assign port_state_out_15_0_0 = state_out_15_0_0;
  assign port_state_out_15_0_1 = state_out_15_0_1;
  assign port_state_out_15_0_2 = state_out_15_0_2;
  assign port_state_out_15_0_3 = state_out_15_0_3;
  assign port_state_out_15_0_4 = state_out_15_0_4;
  assign port_state_out_15_0_5 = state_out_15_0_5;
  assign port_state_out_15_0_6 = state_out_15_0_6;
  assign port_state_out_15_0_7 = state_out_15_0_7;
  assign port_state_out_15_1_0 = state_out_15_1_0;
  assign port_state_out_15_1_1 = state_out_15_1_1;
  assign port_state_out_15_1_2 = state_out_15_1_2;
  assign port_state_out_15_1_3 = state_out_15_1_3;
  assign port_state_out_15_1_4 = state_out_15_1_4;
  assign port_state_out_15_1_5 = state_out_15_1_5;
  assign port_state_out_15_1_6 = state_out_15_1_6;
  assign port_state_out_15_1_7 = state_out_15_1_7;
  assign port_state_out_15_2_0 = state_out_15_2_0;
  assign port_state_out_15_2_1 = state_out_15_2_1;
  assign port_state_out_15_2_2 = state_out_15_2_2;
  assign port_state_out_15_2_3 = state_out_15_2_3;
  assign port_state_out_15_2_4 = state_out_15_2_4;
  assign port_state_out_15_2_5 = state_out_15_2_5;
  assign port_state_out_15_2_6 = state_out_15_2_6;
  assign port_state_out_15_2_7 = state_out_15_2_7;
  assign port_state_out_15_3_0 = state_out_15_3_0;
  assign port_state_out_15_3_1 = state_out_15_3_1;
  assign port_state_out_15_3_2 = state_out_15_3_2;
  assign port_state_out_15_3_3 = state_out_15_3_3;
  assign port_state_out_15_3_4 = state_out_15_3_4;
  assign port_state_out_15_3_5 = state_out_15_3_5;
  assign port_state_out_15_3_6 = state_out_15_3_6;
  assign port_state_out_15_3_7 = state_out_15_3_7;

endmodule

module AES_ShiftRows (
  input      [2:0]    port_state_in_0_0_0,
  input      [2:0]    port_state_in_0_0_1,
  input      [2:0]    port_state_in_0_0_2,
  input      [2:0]    port_state_in_0_0_3,
  input      [2:0]    port_state_in_0_0_4,
  input      [2:0]    port_state_in_0_0_5,
  input      [2:0]    port_state_in_0_0_6,
  input      [2:0]    port_state_in_0_0_7,
  input      [2:0]    port_state_in_0_1_0,
  input      [2:0]    port_state_in_0_1_1,
  input      [2:0]    port_state_in_0_1_2,
  input      [2:0]    port_state_in_0_1_3,
  input      [2:0]    port_state_in_0_1_4,
  input      [2:0]    port_state_in_0_1_5,
  input      [2:0]    port_state_in_0_1_6,
  input      [2:0]    port_state_in_0_1_7,
  input      [2:0]    port_state_in_0_2_0,
  input      [2:0]    port_state_in_0_2_1,
  input      [2:0]    port_state_in_0_2_2,
  input      [2:0]    port_state_in_0_2_3,
  input      [2:0]    port_state_in_0_2_4,
  input      [2:0]    port_state_in_0_2_5,
  input      [2:0]    port_state_in_0_2_6,
  input      [2:0]    port_state_in_0_2_7,
  input      [2:0]    port_state_in_0_3_0,
  input      [2:0]    port_state_in_0_3_1,
  input      [2:0]    port_state_in_0_3_2,
  input      [2:0]    port_state_in_0_3_3,
  input      [2:0]    port_state_in_0_3_4,
  input      [2:0]    port_state_in_0_3_5,
  input      [2:0]    port_state_in_0_3_6,
  input      [2:0]    port_state_in_0_3_7,
  input      [2:0]    port_state_in_1_0_0,
  input      [2:0]    port_state_in_1_0_1,
  input      [2:0]    port_state_in_1_0_2,
  input      [2:0]    port_state_in_1_0_3,
  input      [2:0]    port_state_in_1_0_4,
  input      [2:0]    port_state_in_1_0_5,
  input      [2:0]    port_state_in_1_0_6,
  input      [2:0]    port_state_in_1_0_7,
  input      [2:0]    port_state_in_1_1_0,
  input      [2:0]    port_state_in_1_1_1,
  input      [2:0]    port_state_in_1_1_2,
  input      [2:0]    port_state_in_1_1_3,
  input      [2:0]    port_state_in_1_1_4,
  input      [2:0]    port_state_in_1_1_5,
  input      [2:0]    port_state_in_1_1_6,
  input      [2:0]    port_state_in_1_1_7,
  input      [2:0]    port_state_in_1_2_0,
  input      [2:0]    port_state_in_1_2_1,
  input      [2:0]    port_state_in_1_2_2,
  input      [2:0]    port_state_in_1_2_3,
  input      [2:0]    port_state_in_1_2_4,
  input      [2:0]    port_state_in_1_2_5,
  input      [2:0]    port_state_in_1_2_6,
  input      [2:0]    port_state_in_1_2_7,
  input      [2:0]    port_state_in_1_3_0,
  input      [2:0]    port_state_in_1_3_1,
  input      [2:0]    port_state_in_1_3_2,
  input      [2:0]    port_state_in_1_3_3,
  input      [2:0]    port_state_in_1_3_4,
  input      [2:0]    port_state_in_1_3_5,
  input      [2:0]    port_state_in_1_3_6,
  input      [2:0]    port_state_in_1_3_7,
  input      [2:0]    port_state_in_2_0_0,
  input      [2:0]    port_state_in_2_0_1,
  input      [2:0]    port_state_in_2_0_2,
  input      [2:0]    port_state_in_2_0_3,
  input      [2:0]    port_state_in_2_0_4,
  input      [2:0]    port_state_in_2_0_5,
  input      [2:0]    port_state_in_2_0_6,
  input      [2:0]    port_state_in_2_0_7,
  input      [2:0]    port_state_in_2_1_0,
  input      [2:0]    port_state_in_2_1_1,
  input      [2:0]    port_state_in_2_1_2,
  input      [2:0]    port_state_in_2_1_3,
  input      [2:0]    port_state_in_2_1_4,
  input      [2:0]    port_state_in_2_1_5,
  input      [2:0]    port_state_in_2_1_6,
  input      [2:0]    port_state_in_2_1_7,
  input      [2:0]    port_state_in_2_2_0,
  input      [2:0]    port_state_in_2_2_1,
  input      [2:0]    port_state_in_2_2_2,
  input      [2:0]    port_state_in_2_2_3,
  input      [2:0]    port_state_in_2_2_4,
  input      [2:0]    port_state_in_2_2_5,
  input      [2:0]    port_state_in_2_2_6,
  input      [2:0]    port_state_in_2_2_7,
  input      [2:0]    port_state_in_2_3_0,
  input      [2:0]    port_state_in_2_3_1,
  input      [2:0]    port_state_in_2_3_2,
  input      [2:0]    port_state_in_2_3_3,
  input      [2:0]    port_state_in_2_3_4,
  input      [2:0]    port_state_in_2_3_5,
  input      [2:0]    port_state_in_2_3_6,
  input      [2:0]    port_state_in_2_3_7,
  input      [2:0]    port_state_in_3_0_0,
  input      [2:0]    port_state_in_3_0_1,
  input      [2:0]    port_state_in_3_0_2,
  input      [2:0]    port_state_in_3_0_3,
  input      [2:0]    port_state_in_3_0_4,
  input      [2:0]    port_state_in_3_0_5,
  input      [2:0]    port_state_in_3_0_6,
  input      [2:0]    port_state_in_3_0_7,
  input      [2:0]    port_state_in_3_1_0,
  input      [2:0]    port_state_in_3_1_1,
  input      [2:0]    port_state_in_3_1_2,
  input      [2:0]    port_state_in_3_1_3,
  input      [2:0]    port_state_in_3_1_4,
  input      [2:0]    port_state_in_3_1_5,
  input      [2:0]    port_state_in_3_1_6,
  input      [2:0]    port_state_in_3_1_7,
  input      [2:0]    port_state_in_3_2_0,
  input      [2:0]    port_state_in_3_2_1,
  input      [2:0]    port_state_in_3_2_2,
  input      [2:0]    port_state_in_3_2_3,
  input      [2:0]    port_state_in_3_2_4,
  input      [2:0]    port_state_in_3_2_5,
  input      [2:0]    port_state_in_3_2_6,
  input      [2:0]    port_state_in_3_2_7,
  input      [2:0]    port_state_in_3_3_0,
  input      [2:0]    port_state_in_3_3_1,
  input      [2:0]    port_state_in_3_3_2,
  input      [2:0]    port_state_in_3_3_3,
  input      [2:0]    port_state_in_3_3_4,
  input      [2:0]    port_state_in_3_3_5,
  input      [2:0]    port_state_in_3_3_6,
  input      [2:0]    port_state_in_3_3_7,
  input      [2:0]    port_state_in_4_0_0,
  input      [2:0]    port_state_in_4_0_1,
  input      [2:0]    port_state_in_4_0_2,
  input      [2:0]    port_state_in_4_0_3,
  input      [2:0]    port_state_in_4_0_4,
  input      [2:0]    port_state_in_4_0_5,
  input      [2:0]    port_state_in_4_0_6,
  input      [2:0]    port_state_in_4_0_7,
  input      [2:0]    port_state_in_4_1_0,
  input      [2:0]    port_state_in_4_1_1,
  input      [2:0]    port_state_in_4_1_2,
  input      [2:0]    port_state_in_4_1_3,
  input      [2:0]    port_state_in_4_1_4,
  input      [2:0]    port_state_in_4_1_5,
  input      [2:0]    port_state_in_4_1_6,
  input      [2:0]    port_state_in_4_1_7,
  input      [2:0]    port_state_in_4_2_0,
  input      [2:0]    port_state_in_4_2_1,
  input      [2:0]    port_state_in_4_2_2,
  input      [2:0]    port_state_in_4_2_3,
  input      [2:0]    port_state_in_4_2_4,
  input      [2:0]    port_state_in_4_2_5,
  input      [2:0]    port_state_in_4_2_6,
  input      [2:0]    port_state_in_4_2_7,
  input      [2:0]    port_state_in_4_3_0,
  input      [2:0]    port_state_in_4_3_1,
  input      [2:0]    port_state_in_4_3_2,
  input      [2:0]    port_state_in_4_3_3,
  input      [2:0]    port_state_in_4_3_4,
  input      [2:0]    port_state_in_4_3_5,
  input      [2:0]    port_state_in_4_3_6,
  input      [2:0]    port_state_in_4_3_7,
  input      [2:0]    port_state_in_5_0_0,
  input      [2:0]    port_state_in_5_0_1,
  input      [2:0]    port_state_in_5_0_2,
  input      [2:0]    port_state_in_5_0_3,
  input      [2:0]    port_state_in_5_0_4,
  input      [2:0]    port_state_in_5_0_5,
  input      [2:0]    port_state_in_5_0_6,
  input      [2:0]    port_state_in_5_0_7,
  input      [2:0]    port_state_in_5_1_0,
  input      [2:0]    port_state_in_5_1_1,
  input      [2:0]    port_state_in_5_1_2,
  input      [2:0]    port_state_in_5_1_3,
  input      [2:0]    port_state_in_5_1_4,
  input      [2:0]    port_state_in_5_1_5,
  input      [2:0]    port_state_in_5_1_6,
  input      [2:0]    port_state_in_5_1_7,
  input      [2:0]    port_state_in_5_2_0,
  input      [2:0]    port_state_in_5_2_1,
  input      [2:0]    port_state_in_5_2_2,
  input      [2:0]    port_state_in_5_2_3,
  input      [2:0]    port_state_in_5_2_4,
  input      [2:0]    port_state_in_5_2_5,
  input      [2:0]    port_state_in_5_2_6,
  input      [2:0]    port_state_in_5_2_7,
  input      [2:0]    port_state_in_5_3_0,
  input      [2:0]    port_state_in_5_3_1,
  input      [2:0]    port_state_in_5_3_2,
  input      [2:0]    port_state_in_5_3_3,
  input      [2:0]    port_state_in_5_3_4,
  input      [2:0]    port_state_in_5_3_5,
  input      [2:0]    port_state_in_5_3_6,
  input      [2:0]    port_state_in_5_3_7,
  input      [2:0]    port_state_in_6_0_0,
  input      [2:0]    port_state_in_6_0_1,
  input      [2:0]    port_state_in_6_0_2,
  input      [2:0]    port_state_in_6_0_3,
  input      [2:0]    port_state_in_6_0_4,
  input      [2:0]    port_state_in_6_0_5,
  input      [2:0]    port_state_in_6_0_6,
  input      [2:0]    port_state_in_6_0_7,
  input      [2:0]    port_state_in_6_1_0,
  input      [2:0]    port_state_in_6_1_1,
  input      [2:0]    port_state_in_6_1_2,
  input      [2:0]    port_state_in_6_1_3,
  input      [2:0]    port_state_in_6_1_4,
  input      [2:0]    port_state_in_6_1_5,
  input      [2:0]    port_state_in_6_1_6,
  input      [2:0]    port_state_in_6_1_7,
  input      [2:0]    port_state_in_6_2_0,
  input      [2:0]    port_state_in_6_2_1,
  input      [2:0]    port_state_in_6_2_2,
  input      [2:0]    port_state_in_6_2_3,
  input      [2:0]    port_state_in_6_2_4,
  input      [2:0]    port_state_in_6_2_5,
  input      [2:0]    port_state_in_6_2_6,
  input      [2:0]    port_state_in_6_2_7,
  input      [2:0]    port_state_in_6_3_0,
  input      [2:0]    port_state_in_6_3_1,
  input      [2:0]    port_state_in_6_3_2,
  input      [2:0]    port_state_in_6_3_3,
  input      [2:0]    port_state_in_6_3_4,
  input      [2:0]    port_state_in_6_3_5,
  input      [2:0]    port_state_in_6_3_6,
  input      [2:0]    port_state_in_6_3_7,
  input      [2:0]    port_state_in_7_0_0,
  input      [2:0]    port_state_in_7_0_1,
  input      [2:0]    port_state_in_7_0_2,
  input      [2:0]    port_state_in_7_0_3,
  input      [2:0]    port_state_in_7_0_4,
  input      [2:0]    port_state_in_7_0_5,
  input      [2:0]    port_state_in_7_0_6,
  input      [2:0]    port_state_in_7_0_7,
  input      [2:0]    port_state_in_7_1_0,
  input      [2:0]    port_state_in_7_1_1,
  input      [2:0]    port_state_in_7_1_2,
  input      [2:0]    port_state_in_7_1_3,
  input      [2:0]    port_state_in_7_1_4,
  input      [2:0]    port_state_in_7_1_5,
  input      [2:0]    port_state_in_7_1_6,
  input      [2:0]    port_state_in_7_1_7,
  input      [2:0]    port_state_in_7_2_0,
  input      [2:0]    port_state_in_7_2_1,
  input      [2:0]    port_state_in_7_2_2,
  input      [2:0]    port_state_in_7_2_3,
  input      [2:0]    port_state_in_7_2_4,
  input      [2:0]    port_state_in_7_2_5,
  input      [2:0]    port_state_in_7_2_6,
  input      [2:0]    port_state_in_7_2_7,
  input      [2:0]    port_state_in_7_3_0,
  input      [2:0]    port_state_in_7_3_1,
  input      [2:0]    port_state_in_7_3_2,
  input      [2:0]    port_state_in_7_3_3,
  input      [2:0]    port_state_in_7_3_4,
  input      [2:0]    port_state_in_7_3_5,
  input      [2:0]    port_state_in_7_3_6,
  input      [2:0]    port_state_in_7_3_7,
  input      [2:0]    port_state_in_8_0_0,
  input      [2:0]    port_state_in_8_0_1,
  input      [2:0]    port_state_in_8_0_2,
  input      [2:0]    port_state_in_8_0_3,
  input      [2:0]    port_state_in_8_0_4,
  input      [2:0]    port_state_in_8_0_5,
  input      [2:0]    port_state_in_8_0_6,
  input      [2:0]    port_state_in_8_0_7,
  input      [2:0]    port_state_in_8_1_0,
  input      [2:0]    port_state_in_8_1_1,
  input      [2:0]    port_state_in_8_1_2,
  input      [2:0]    port_state_in_8_1_3,
  input      [2:0]    port_state_in_8_1_4,
  input      [2:0]    port_state_in_8_1_5,
  input      [2:0]    port_state_in_8_1_6,
  input      [2:0]    port_state_in_8_1_7,
  input      [2:0]    port_state_in_8_2_0,
  input      [2:0]    port_state_in_8_2_1,
  input      [2:0]    port_state_in_8_2_2,
  input      [2:0]    port_state_in_8_2_3,
  input      [2:0]    port_state_in_8_2_4,
  input      [2:0]    port_state_in_8_2_5,
  input      [2:0]    port_state_in_8_2_6,
  input      [2:0]    port_state_in_8_2_7,
  input      [2:0]    port_state_in_8_3_0,
  input      [2:0]    port_state_in_8_3_1,
  input      [2:0]    port_state_in_8_3_2,
  input      [2:0]    port_state_in_8_3_3,
  input      [2:0]    port_state_in_8_3_4,
  input      [2:0]    port_state_in_8_3_5,
  input      [2:0]    port_state_in_8_3_6,
  input      [2:0]    port_state_in_8_3_7,
  input      [2:0]    port_state_in_9_0_0,
  input      [2:0]    port_state_in_9_0_1,
  input      [2:0]    port_state_in_9_0_2,
  input      [2:0]    port_state_in_9_0_3,
  input      [2:0]    port_state_in_9_0_4,
  input      [2:0]    port_state_in_9_0_5,
  input      [2:0]    port_state_in_9_0_6,
  input      [2:0]    port_state_in_9_0_7,
  input      [2:0]    port_state_in_9_1_0,
  input      [2:0]    port_state_in_9_1_1,
  input      [2:0]    port_state_in_9_1_2,
  input      [2:0]    port_state_in_9_1_3,
  input      [2:0]    port_state_in_9_1_4,
  input      [2:0]    port_state_in_9_1_5,
  input      [2:0]    port_state_in_9_1_6,
  input      [2:0]    port_state_in_9_1_7,
  input      [2:0]    port_state_in_9_2_0,
  input      [2:0]    port_state_in_9_2_1,
  input      [2:0]    port_state_in_9_2_2,
  input      [2:0]    port_state_in_9_2_3,
  input      [2:0]    port_state_in_9_2_4,
  input      [2:0]    port_state_in_9_2_5,
  input      [2:0]    port_state_in_9_2_6,
  input      [2:0]    port_state_in_9_2_7,
  input      [2:0]    port_state_in_9_3_0,
  input      [2:0]    port_state_in_9_3_1,
  input      [2:0]    port_state_in_9_3_2,
  input      [2:0]    port_state_in_9_3_3,
  input      [2:0]    port_state_in_9_3_4,
  input      [2:0]    port_state_in_9_3_5,
  input      [2:0]    port_state_in_9_3_6,
  input      [2:0]    port_state_in_9_3_7,
  input      [2:0]    port_state_in_10_0_0,
  input      [2:0]    port_state_in_10_0_1,
  input      [2:0]    port_state_in_10_0_2,
  input      [2:0]    port_state_in_10_0_3,
  input      [2:0]    port_state_in_10_0_4,
  input      [2:0]    port_state_in_10_0_5,
  input      [2:0]    port_state_in_10_0_6,
  input      [2:0]    port_state_in_10_0_7,
  input      [2:0]    port_state_in_10_1_0,
  input      [2:0]    port_state_in_10_1_1,
  input      [2:0]    port_state_in_10_1_2,
  input      [2:0]    port_state_in_10_1_3,
  input      [2:0]    port_state_in_10_1_4,
  input      [2:0]    port_state_in_10_1_5,
  input      [2:0]    port_state_in_10_1_6,
  input      [2:0]    port_state_in_10_1_7,
  input      [2:0]    port_state_in_10_2_0,
  input      [2:0]    port_state_in_10_2_1,
  input      [2:0]    port_state_in_10_2_2,
  input      [2:0]    port_state_in_10_2_3,
  input      [2:0]    port_state_in_10_2_4,
  input      [2:0]    port_state_in_10_2_5,
  input      [2:0]    port_state_in_10_2_6,
  input      [2:0]    port_state_in_10_2_7,
  input      [2:0]    port_state_in_10_3_0,
  input      [2:0]    port_state_in_10_3_1,
  input      [2:0]    port_state_in_10_3_2,
  input      [2:0]    port_state_in_10_3_3,
  input      [2:0]    port_state_in_10_3_4,
  input      [2:0]    port_state_in_10_3_5,
  input      [2:0]    port_state_in_10_3_6,
  input      [2:0]    port_state_in_10_3_7,
  input      [2:0]    port_state_in_11_0_0,
  input      [2:0]    port_state_in_11_0_1,
  input      [2:0]    port_state_in_11_0_2,
  input      [2:0]    port_state_in_11_0_3,
  input      [2:0]    port_state_in_11_0_4,
  input      [2:0]    port_state_in_11_0_5,
  input      [2:0]    port_state_in_11_0_6,
  input      [2:0]    port_state_in_11_0_7,
  input      [2:0]    port_state_in_11_1_0,
  input      [2:0]    port_state_in_11_1_1,
  input      [2:0]    port_state_in_11_1_2,
  input      [2:0]    port_state_in_11_1_3,
  input      [2:0]    port_state_in_11_1_4,
  input      [2:0]    port_state_in_11_1_5,
  input      [2:0]    port_state_in_11_1_6,
  input      [2:0]    port_state_in_11_1_7,
  input      [2:0]    port_state_in_11_2_0,
  input      [2:0]    port_state_in_11_2_1,
  input      [2:0]    port_state_in_11_2_2,
  input      [2:0]    port_state_in_11_2_3,
  input      [2:0]    port_state_in_11_2_4,
  input      [2:0]    port_state_in_11_2_5,
  input      [2:0]    port_state_in_11_2_6,
  input      [2:0]    port_state_in_11_2_7,
  input      [2:0]    port_state_in_11_3_0,
  input      [2:0]    port_state_in_11_3_1,
  input      [2:0]    port_state_in_11_3_2,
  input      [2:0]    port_state_in_11_3_3,
  input      [2:0]    port_state_in_11_3_4,
  input      [2:0]    port_state_in_11_3_5,
  input      [2:0]    port_state_in_11_3_6,
  input      [2:0]    port_state_in_11_3_7,
  input      [2:0]    port_state_in_12_0_0,
  input      [2:0]    port_state_in_12_0_1,
  input      [2:0]    port_state_in_12_0_2,
  input      [2:0]    port_state_in_12_0_3,
  input      [2:0]    port_state_in_12_0_4,
  input      [2:0]    port_state_in_12_0_5,
  input      [2:0]    port_state_in_12_0_6,
  input      [2:0]    port_state_in_12_0_7,
  input      [2:0]    port_state_in_12_1_0,
  input      [2:0]    port_state_in_12_1_1,
  input      [2:0]    port_state_in_12_1_2,
  input      [2:0]    port_state_in_12_1_3,
  input      [2:0]    port_state_in_12_1_4,
  input      [2:0]    port_state_in_12_1_5,
  input      [2:0]    port_state_in_12_1_6,
  input      [2:0]    port_state_in_12_1_7,
  input      [2:0]    port_state_in_12_2_0,
  input      [2:0]    port_state_in_12_2_1,
  input      [2:0]    port_state_in_12_2_2,
  input      [2:0]    port_state_in_12_2_3,
  input      [2:0]    port_state_in_12_2_4,
  input      [2:0]    port_state_in_12_2_5,
  input      [2:0]    port_state_in_12_2_6,
  input      [2:0]    port_state_in_12_2_7,
  input      [2:0]    port_state_in_12_3_0,
  input      [2:0]    port_state_in_12_3_1,
  input      [2:0]    port_state_in_12_3_2,
  input      [2:0]    port_state_in_12_3_3,
  input      [2:0]    port_state_in_12_3_4,
  input      [2:0]    port_state_in_12_3_5,
  input      [2:0]    port_state_in_12_3_6,
  input      [2:0]    port_state_in_12_3_7,
  input      [2:0]    port_state_in_13_0_0,
  input      [2:0]    port_state_in_13_0_1,
  input      [2:0]    port_state_in_13_0_2,
  input      [2:0]    port_state_in_13_0_3,
  input      [2:0]    port_state_in_13_0_4,
  input      [2:0]    port_state_in_13_0_5,
  input      [2:0]    port_state_in_13_0_6,
  input      [2:0]    port_state_in_13_0_7,
  input      [2:0]    port_state_in_13_1_0,
  input      [2:0]    port_state_in_13_1_1,
  input      [2:0]    port_state_in_13_1_2,
  input      [2:0]    port_state_in_13_1_3,
  input      [2:0]    port_state_in_13_1_4,
  input      [2:0]    port_state_in_13_1_5,
  input      [2:0]    port_state_in_13_1_6,
  input      [2:0]    port_state_in_13_1_7,
  input      [2:0]    port_state_in_13_2_0,
  input      [2:0]    port_state_in_13_2_1,
  input      [2:0]    port_state_in_13_2_2,
  input      [2:0]    port_state_in_13_2_3,
  input      [2:0]    port_state_in_13_2_4,
  input      [2:0]    port_state_in_13_2_5,
  input      [2:0]    port_state_in_13_2_6,
  input      [2:0]    port_state_in_13_2_7,
  input      [2:0]    port_state_in_13_3_0,
  input      [2:0]    port_state_in_13_3_1,
  input      [2:0]    port_state_in_13_3_2,
  input      [2:0]    port_state_in_13_3_3,
  input      [2:0]    port_state_in_13_3_4,
  input      [2:0]    port_state_in_13_3_5,
  input      [2:0]    port_state_in_13_3_6,
  input      [2:0]    port_state_in_13_3_7,
  input      [2:0]    port_state_in_14_0_0,
  input      [2:0]    port_state_in_14_0_1,
  input      [2:0]    port_state_in_14_0_2,
  input      [2:0]    port_state_in_14_0_3,
  input      [2:0]    port_state_in_14_0_4,
  input      [2:0]    port_state_in_14_0_5,
  input      [2:0]    port_state_in_14_0_6,
  input      [2:0]    port_state_in_14_0_7,
  input      [2:0]    port_state_in_14_1_0,
  input      [2:0]    port_state_in_14_1_1,
  input      [2:0]    port_state_in_14_1_2,
  input      [2:0]    port_state_in_14_1_3,
  input      [2:0]    port_state_in_14_1_4,
  input      [2:0]    port_state_in_14_1_5,
  input      [2:0]    port_state_in_14_1_6,
  input      [2:0]    port_state_in_14_1_7,
  input      [2:0]    port_state_in_14_2_0,
  input      [2:0]    port_state_in_14_2_1,
  input      [2:0]    port_state_in_14_2_2,
  input      [2:0]    port_state_in_14_2_3,
  input      [2:0]    port_state_in_14_2_4,
  input      [2:0]    port_state_in_14_2_5,
  input      [2:0]    port_state_in_14_2_6,
  input      [2:0]    port_state_in_14_2_7,
  input      [2:0]    port_state_in_14_3_0,
  input      [2:0]    port_state_in_14_3_1,
  input      [2:0]    port_state_in_14_3_2,
  input      [2:0]    port_state_in_14_3_3,
  input      [2:0]    port_state_in_14_3_4,
  input      [2:0]    port_state_in_14_3_5,
  input      [2:0]    port_state_in_14_3_6,
  input      [2:0]    port_state_in_14_3_7,
  input      [2:0]    port_state_in_15_0_0,
  input      [2:0]    port_state_in_15_0_1,
  input      [2:0]    port_state_in_15_0_2,
  input      [2:0]    port_state_in_15_0_3,
  input      [2:0]    port_state_in_15_0_4,
  input      [2:0]    port_state_in_15_0_5,
  input      [2:0]    port_state_in_15_0_6,
  input      [2:0]    port_state_in_15_0_7,
  input      [2:0]    port_state_in_15_1_0,
  input      [2:0]    port_state_in_15_1_1,
  input      [2:0]    port_state_in_15_1_2,
  input      [2:0]    port_state_in_15_1_3,
  input      [2:0]    port_state_in_15_1_4,
  input      [2:0]    port_state_in_15_1_5,
  input      [2:0]    port_state_in_15_1_6,
  input      [2:0]    port_state_in_15_1_7,
  input      [2:0]    port_state_in_15_2_0,
  input      [2:0]    port_state_in_15_2_1,
  input      [2:0]    port_state_in_15_2_2,
  input      [2:0]    port_state_in_15_2_3,
  input      [2:0]    port_state_in_15_2_4,
  input      [2:0]    port_state_in_15_2_5,
  input      [2:0]    port_state_in_15_2_6,
  input      [2:0]    port_state_in_15_2_7,
  input      [2:0]    port_state_in_15_3_0,
  input      [2:0]    port_state_in_15_3_1,
  input      [2:0]    port_state_in_15_3_2,
  input      [2:0]    port_state_in_15_3_3,
  input      [2:0]    port_state_in_15_3_4,
  input      [2:0]    port_state_in_15_3_5,
  input      [2:0]    port_state_in_15_3_6,
  input      [2:0]    port_state_in_15_3_7,
  output     [2:0]    port_state_out_0_0_0,
  output     [2:0]    port_state_out_0_0_1,
  output     [2:0]    port_state_out_0_0_2,
  output     [2:0]    port_state_out_0_0_3,
  output     [2:0]    port_state_out_0_0_4,
  output     [2:0]    port_state_out_0_0_5,
  output     [2:0]    port_state_out_0_0_6,
  output     [2:0]    port_state_out_0_0_7,
  output     [2:0]    port_state_out_0_1_0,
  output     [2:0]    port_state_out_0_1_1,
  output     [2:0]    port_state_out_0_1_2,
  output     [2:0]    port_state_out_0_1_3,
  output     [2:0]    port_state_out_0_1_4,
  output     [2:0]    port_state_out_0_1_5,
  output     [2:0]    port_state_out_0_1_6,
  output     [2:0]    port_state_out_0_1_7,
  output     [2:0]    port_state_out_0_2_0,
  output     [2:0]    port_state_out_0_2_1,
  output     [2:0]    port_state_out_0_2_2,
  output     [2:0]    port_state_out_0_2_3,
  output     [2:0]    port_state_out_0_2_4,
  output     [2:0]    port_state_out_0_2_5,
  output     [2:0]    port_state_out_0_2_6,
  output     [2:0]    port_state_out_0_2_7,
  output     [2:0]    port_state_out_0_3_0,
  output     [2:0]    port_state_out_0_3_1,
  output     [2:0]    port_state_out_0_3_2,
  output     [2:0]    port_state_out_0_3_3,
  output     [2:0]    port_state_out_0_3_4,
  output     [2:0]    port_state_out_0_3_5,
  output     [2:0]    port_state_out_0_3_6,
  output     [2:0]    port_state_out_0_3_7,
  output     [2:0]    port_state_out_1_0_0,
  output     [2:0]    port_state_out_1_0_1,
  output     [2:0]    port_state_out_1_0_2,
  output     [2:0]    port_state_out_1_0_3,
  output     [2:0]    port_state_out_1_0_4,
  output     [2:0]    port_state_out_1_0_5,
  output     [2:0]    port_state_out_1_0_6,
  output     [2:0]    port_state_out_1_0_7,
  output     [2:0]    port_state_out_1_1_0,
  output     [2:0]    port_state_out_1_1_1,
  output     [2:0]    port_state_out_1_1_2,
  output     [2:0]    port_state_out_1_1_3,
  output     [2:0]    port_state_out_1_1_4,
  output     [2:0]    port_state_out_1_1_5,
  output     [2:0]    port_state_out_1_1_6,
  output     [2:0]    port_state_out_1_1_7,
  output     [2:0]    port_state_out_1_2_0,
  output     [2:0]    port_state_out_1_2_1,
  output     [2:0]    port_state_out_1_2_2,
  output     [2:0]    port_state_out_1_2_3,
  output     [2:0]    port_state_out_1_2_4,
  output     [2:0]    port_state_out_1_2_5,
  output     [2:0]    port_state_out_1_2_6,
  output     [2:0]    port_state_out_1_2_7,
  output     [2:0]    port_state_out_1_3_0,
  output     [2:0]    port_state_out_1_3_1,
  output     [2:0]    port_state_out_1_3_2,
  output     [2:0]    port_state_out_1_3_3,
  output     [2:0]    port_state_out_1_3_4,
  output     [2:0]    port_state_out_1_3_5,
  output     [2:0]    port_state_out_1_3_6,
  output     [2:0]    port_state_out_1_3_7,
  output     [2:0]    port_state_out_2_0_0,
  output     [2:0]    port_state_out_2_0_1,
  output     [2:0]    port_state_out_2_0_2,
  output     [2:0]    port_state_out_2_0_3,
  output     [2:0]    port_state_out_2_0_4,
  output     [2:0]    port_state_out_2_0_5,
  output     [2:0]    port_state_out_2_0_6,
  output     [2:0]    port_state_out_2_0_7,
  output     [2:0]    port_state_out_2_1_0,
  output     [2:0]    port_state_out_2_1_1,
  output     [2:0]    port_state_out_2_1_2,
  output     [2:0]    port_state_out_2_1_3,
  output     [2:0]    port_state_out_2_1_4,
  output     [2:0]    port_state_out_2_1_5,
  output     [2:0]    port_state_out_2_1_6,
  output     [2:0]    port_state_out_2_1_7,
  output     [2:0]    port_state_out_2_2_0,
  output     [2:0]    port_state_out_2_2_1,
  output     [2:0]    port_state_out_2_2_2,
  output     [2:0]    port_state_out_2_2_3,
  output     [2:0]    port_state_out_2_2_4,
  output     [2:0]    port_state_out_2_2_5,
  output     [2:0]    port_state_out_2_2_6,
  output     [2:0]    port_state_out_2_2_7,
  output     [2:0]    port_state_out_2_3_0,
  output     [2:0]    port_state_out_2_3_1,
  output     [2:0]    port_state_out_2_3_2,
  output     [2:0]    port_state_out_2_3_3,
  output     [2:0]    port_state_out_2_3_4,
  output     [2:0]    port_state_out_2_3_5,
  output     [2:0]    port_state_out_2_3_6,
  output     [2:0]    port_state_out_2_3_7,
  output     [2:0]    port_state_out_3_0_0,
  output     [2:0]    port_state_out_3_0_1,
  output     [2:0]    port_state_out_3_0_2,
  output     [2:0]    port_state_out_3_0_3,
  output     [2:0]    port_state_out_3_0_4,
  output     [2:0]    port_state_out_3_0_5,
  output     [2:0]    port_state_out_3_0_6,
  output     [2:0]    port_state_out_3_0_7,
  output     [2:0]    port_state_out_3_1_0,
  output     [2:0]    port_state_out_3_1_1,
  output     [2:0]    port_state_out_3_1_2,
  output     [2:0]    port_state_out_3_1_3,
  output     [2:0]    port_state_out_3_1_4,
  output     [2:0]    port_state_out_3_1_5,
  output     [2:0]    port_state_out_3_1_6,
  output     [2:0]    port_state_out_3_1_7,
  output     [2:0]    port_state_out_3_2_0,
  output     [2:0]    port_state_out_3_2_1,
  output     [2:0]    port_state_out_3_2_2,
  output     [2:0]    port_state_out_3_2_3,
  output     [2:0]    port_state_out_3_2_4,
  output     [2:0]    port_state_out_3_2_5,
  output     [2:0]    port_state_out_3_2_6,
  output     [2:0]    port_state_out_3_2_7,
  output     [2:0]    port_state_out_3_3_0,
  output     [2:0]    port_state_out_3_3_1,
  output     [2:0]    port_state_out_3_3_2,
  output     [2:0]    port_state_out_3_3_3,
  output     [2:0]    port_state_out_3_3_4,
  output     [2:0]    port_state_out_3_3_5,
  output     [2:0]    port_state_out_3_3_6,
  output     [2:0]    port_state_out_3_3_7,
  output     [2:0]    port_state_out_4_0_0,
  output     [2:0]    port_state_out_4_0_1,
  output     [2:0]    port_state_out_4_0_2,
  output     [2:0]    port_state_out_4_0_3,
  output     [2:0]    port_state_out_4_0_4,
  output     [2:0]    port_state_out_4_0_5,
  output     [2:0]    port_state_out_4_0_6,
  output     [2:0]    port_state_out_4_0_7,
  output     [2:0]    port_state_out_4_1_0,
  output     [2:0]    port_state_out_4_1_1,
  output     [2:0]    port_state_out_4_1_2,
  output     [2:0]    port_state_out_4_1_3,
  output     [2:0]    port_state_out_4_1_4,
  output     [2:0]    port_state_out_4_1_5,
  output     [2:0]    port_state_out_4_1_6,
  output     [2:0]    port_state_out_4_1_7,
  output     [2:0]    port_state_out_4_2_0,
  output     [2:0]    port_state_out_4_2_1,
  output     [2:0]    port_state_out_4_2_2,
  output     [2:0]    port_state_out_4_2_3,
  output     [2:0]    port_state_out_4_2_4,
  output     [2:0]    port_state_out_4_2_5,
  output     [2:0]    port_state_out_4_2_6,
  output     [2:0]    port_state_out_4_2_7,
  output     [2:0]    port_state_out_4_3_0,
  output     [2:0]    port_state_out_4_3_1,
  output     [2:0]    port_state_out_4_3_2,
  output     [2:0]    port_state_out_4_3_3,
  output     [2:0]    port_state_out_4_3_4,
  output     [2:0]    port_state_out_4_3_5,
  output     [2:0]    port_state_out_4_3_6,
  output     [2:0]    port_state_out_4_3_7,
  output     [2:0]    port_state_out_5_0_0,
  output     [2:0]    port_state_out_5_0_1,
  output     [2:0]    port_state_out_5_0_2,
  output     [2:0]    port_state_out_5_0_3,
  output     [2:0]    port_state_out_5_0_4,
  output     [2:0]    port_state_out_5_0_5,
  output     [2:0]    port_state_out_5_0_6,
  output     [2:0]    port_state_out_5_0_7,
  output     [2:0]    port_state_out_5_1_0,
  output     [2:0]    port_state_out_5_1_1,
  output     [2:0]    port_state_out_5_1_2,
  output     [2:0]    port_state_out_5_1_3,
  output     [2:0]    port_state_out_5_1_4,
  output     [2:0]    port_state_out_5_1_5,
  output     [2:0]    port_state_out_5_1_6,
  output     [2:0]    port_state_out_5_1_7,
  output     [2:0]    port_state_out_5_2_0,
  output     [2:0]    port_state_out_5_2_1,
  output     [2:0]    port_state_out_5_2_2,
  output     [2:0]    port_state_out_5_2_3,
  output     [2:0]    port_state_out_5_2_4,
  output     [2:0]    port_state_out_5_2_5,
  output     [2:0]    port_state_out_5_2_6,
  output     [2:0]    port_state_out_5_2_7,
  output     [2:0]    port_state_out_5_3_0,
  output     [2:0]    port_state_out_5_3_1,
  output     [2:0]    port_state_out_5_3_2,
  output     [2:0]    port_state_out_5_3_3,
  output     [2:0]    port_state_out_5_3_4,
  output     [2:0]    port_state_out_5_3_5,
  output     [2:0]    port_state_out_5_3_6,
  output     [2:0]    port_state_out_5_3_7,
  output     [2:0]    port_state_out_6_0_0,
  output     [2:0]    port_state_out_6_0_1,
  output     [2:0]    port_state_out_6_0_2,
  output     [2:0]    port_state_out_6_0_3,
  output     [2:0]    port_state_out_6_0_4,
  output     [2:0]    port_state_out_6_0_5,
  output     [2:0]    port_state_out_6_0_6,
  output     [2:0]    port_state_out_6_0_7,
  output     [2:0]    port_state_out_6_1_0,
  output     [2:0]    port_state_out_6_1_1,
  output     [2:0]    port_state_out_6_1_2,
  output     [2:0]    port_state_out_6_1_3,
  output     [2:0]    port_state_out_6_1_4,
  output     [2:0]    port_state_out_6_1_5,
  output     [2:0]    port_state_out_6_1_6,
  output     [2:0]    port_state_out_6_1_7,
  output     [2:0]    port_state_out_6_2_0,
  output     [2:0]    port_state_out_6_2_1,
  output     [2:0]    port_state_out_6_2_2,
  output     [2:0]    port_state_out_6_2_3,
  output     [2:0]    port_state_out_6_2_4,
  output     [2:0]    port_state_out_6_2_5,
  output     [2:0]    port_state_out_6_2_6,
  output     [2:0]    port_state_out_6_2_7,
  output     [2:0]    port_state_out_6_3_0,
  output     [2:0]    port_state_out_6_3_1,
  output     [2:0]    port_state_out_6_3_2,
  output     [2:0]    port_state_out_6_3_3,
  output     [2:0]    port_state_out_6_3_4,
  output     [2:0]    port_state_out_6_3_5,
  output     [2:0]    port_state_out_6_3_6,
  output     [2:0]    port_state_out_6_3_7,
  output     [2:0]    port_state_out_7_0_0,
  output     [2:0]    port_state_out_7_0_1,
  output     [2:0]    port_state_out_7_0_2,
  output     [2:0]    port_state_out_7_0_3,
  output     [2:0]    port_state_out_7_0_4,
  output     [2:0]    port_state_out_7_0_5,
  output     [2:0]    port_state_out_7_0_6,
  output     [2:0]    port_state_out_7_0_7,
  output     [2:0]    port_state_out_7_1_0,
  output     [2:0]    port_state_out_7_1_1,
  output     [2:0]    port_state_out_7_1_2,
  output     [2:0]    port_state_out_7_1_3,
  output     [2:0]    port_state_out_7_1_4,
  output     [2:0]    port_state_out_7_1_5,
  output     [2:0]    port_state_out_7_1_6,
  output     [2:0]    port_state_out_7_1_7,
  output     [2:0]    port_state_out_7_2_0,
  output     [2:0]    port_state_out_7_2_1,
  output     [2:0]    port_state_out_7_2_2,
  output     [2:0]    port_state_out_7_2_3,
  output     [2:0]    port_state_out_7_2_4,
  output     [2:0]    port_state_out_7_2_5,
  output     [2:0]    port_state_out_7_2_6,
  output     [2:0]    port_state_out_7_2_7,
  output     [2:0]    port_state_out_7_3_0,
  output     [2:0]    port_state_out_7_3_1,
  output     [2:0]    port_state_out_7_3_2,
  output     [2:0]    port_state_out_7_3_3,
  output     [2:0]    port_state_out_7_3_4,
  output     [2:0]    port_state_out_7_3_5,
  output     [2:0]    port_state_out_7_3_6,
  output     [2:0]    port_state_out_7_3_7,
  output     [2:0]    port_state_out_8_0_0,
  output     [2:0]    port_state_out_8_0_1,
  output     [2:0]    port_state_out_8_0_2,
  output     [2:0]    port_state_out_8_0_3,
  output     [2:0]    port_state_out_8_0_4,
  output     [2:0]    port_state_out_8_0_5,
  output     [2:0]    port_state_out_8_0_6,
  output     [2:0]    port_state_out_8_0_7,
  output     [2:0]    port_state_out_8_1_0,
  output     [2:0]    port_state_out_8_1_1,
  output     [2:0]    port_state_out_8_1_2,
  output     [2:0]    port_state_out_8_1_3,
  output     [2:0]    port_state_out_8_1_4,
  output     [2:0]    port_state_out_8_1_5,
  output     [2:0]    port_state_out_8_1_6,
  output     [2:0]    port_state_out_8_1_7,
  output     [2:0]    port_state_out_8_2_0,
  output     [2:0]    port_state_out_8_2_1,
  output     [2:0]    port_state_out_8_2_2,
  output     [2:0]    port_state_out_8_2_3,
  output     [2:0]    port_state_out_8_2_4,
  output     [2:0]    port_state_out_8_2_5,
  output     [2:0]    port_state_out_8_2_6,
  output     [2:0]    port_state_out_8_2_7,
  output     [2:0]    port_state_out_8_3_0,
  output     [2:0]    port_state_out_8_3_1,
  output     [2:0]    port_state_out_8_3_2,
  output     [2:0]    port_state_out_8_3_3,
  output     [2:0]    port_state_out_8_3_4,
  output     [2:0]    port_state_out_8_3_5,
  output     [2:0]    port_state_out_8_3_6,
  output     [2:0]    port_state_out_8_3_7,
  output     [2:0]    port_state_out_9_0_0,
  output     [2:0]    port_state_out_9_0_1,
  output     [2:0]    port_state_out_9_0_2,
  output     [2:0]    port_state_out_9_0_3,
  output     [2:0]    port_state_out_9_0_4,
  output     [2:0]    port_state_out_9_0_5,
  output     [2:0]    port_state_out_9_0_6,
  output     [2:0]    port_state_out_9_0_7,
  output     [2:0]    port_state_out_9_1_0,
  output     [2:0]    port_state_out_9_1_1,
  output     [2:0]    port_state_out_9_1_2,
  output     [2:0]    port_state_out_9_1_3,
  output     [2:0]    port_state_out_9_1_4,
  output     [2:0]    port_state_out_9_1_5,
  output     [2:0]    port_state_out_9_1_6,
  output     [2:0]    port_state_out_9_1_7,
  output     [2:0]    port_state_out_9_2_0,
  output     [2:0]    port_state_out_9_2_1,
  output     [2:0]    port_state_out_9_2_2,
  output     [2:0]    port_state_out_9_2_3,
  output     [2:0]    port_state_out_9_2_4,
  output     [2:0]    port_state_out_9_2_5,
  output     [2:0]    port_state_out_9_2_6,
  output     [2:0]    port_state_out_9_2_7,
  output     [2:0]    port_state_out_9_3_0,
  output     [2:0]    port_state_out_9_3_1,
  output     [2:0]    port_state_out_9_3_2,
  output     [2:0]    port_state_out_9_3_3,
  output     [2:0]    port_state_out_9_3_4,
  output     [2:0]    port_state_out_9_3_5,
  output     [2:0]    port_state_out_9_3_6,
  output     [2:0]    port_state_out_9_3_7,
  output     [2:0]    port_state_out_10_0_0,
  output     [2:0]    port_state_out_10_0_1,
  output     [2:0]    port_state_out_10_0_2,
  output     [2:0]    port_state_out_10_0_3,
  output     [2:0]    port_state_out_10_0_4,
  output     [2:0]    port_state_out_10_0_5,
  output     [2:0]    port_state_out_10_0_6,
  output     [2:0]    port_state_out_10_0_7,
  output     [2:0]    port_state_out_10_1_0,
  output     [2:0]    port_state_out_10_1_1,
  output     [2:0]    port_state_out_10_1_2,
  output     [2:0]    port_state_out_10_1_3,
  output     [2:0]    port_state_out_10_1_4,
  output     [2:0]    port_state_out_10_1_5,
  output     [2:0]    port_state_out_10_1_6,
  output     [2:0]    port_state_out_10_1_7,
  output     [2:0]    port_state_out_10_2_0,
  output     [2:0]    port_state_out_10_2_1,
  output     [2:0]    port_state_out_10_2_2,
  output     [2:0]    port_state_out_10_2_3,
  output     [2:0]    port_state_out_10_2_4,
  output     [2:0]    port_state_out_10_2_5,
  output     [2:0]    port_state_out_10_2_6,
  output     [2:0]    port_state_out_10_2_7,
  output     [2:0]    port_state_out_10_3_0,
  output     [2:0]    port_state_out_10_3_1,
  output     [2:0]    port_state_out_10_3_2,
  output     [2:0]    port_state_out_10_3_3,
  output     [2:0]    port_state_out_10_3_4,
  output     [2:0]    port_state_out_10_3_5,
  output     [2:0]    port_state_out_10_3_6,
  output     [2:0]    port_state_out_10_3_7,
  output     [2:0]    port_state_out_11_0_0,
  output     [2:0]    port_state_out_11_0_1,
  output     [2:0]    port_state_out_11_0_2,
  output     [2:0]    port_state_out_11_0_3,
  output     [2:0]    port_state_out_11_0_4,
  output     [2:0]    port_state_out_11_0_5,
  output     [2:0]    port_state_out_11_0_6,
  output     [2:0]    port_state_out_11_0_7,
  output     [2:0]    port_state_out_11_1_0,
  output     [2:0]    port_state_out_11_1_1,
  output     [2:0]    port_state_out_11_1_2,
  output     [2:0]    port_state_out_11_1_3,
  output     [2:0]    port_state_out_11_1_4,
  output     [2:0]    port_state_out_11_1_5,
  output     [2:0]    port_state_out_11_1_6,
  output     [2:0]    port_state_out_11_1_7,
  output     [2:0]    port_state_out_11_2_0,
  output     [2:0]    port_state_out_11_2_1,
  output     [2:0]    port_state_out_11_2_2,
  output     [2:0]    port_state_out_11_2_3,
  output     [2:0]    port_state_out_11_2_4,
  output     [2:0]    port_state_out_11_2_5,
  output     [2:0]    port_state_out_11_2_6,
  output     [2:0]    port_state_out_11_2_7,
  output     [2:0]    port_state_out_11_3_0,
  output     [2:0]    port_state_out_11_3_1,
  output     [2:0]    port_state_out_11_3_2,
  output     [2:0]    port_state_out_11_3_3,
  output     [2:0]    port_state_out_11_3_4,
  output     [2:0]    port_state_out_11_3_5,
  output     [2:0]    port_state_out_11_3_6,
  output     [2:0]    port_state_out_11_3_7,
  output     [2:0]    port_state_out_12_0_0,
  output     [2:0]    port_state_out_12_0_1,
  output     [2:0]    port_state_out_12_0_2,
  output     [2:0]    port_state_out_12_0_3,
  output     [2:0]    port_state_out_12_0_4,
  output     [2:0]    port_state_out_12_0_5,
  output     [2:0]    port_state_out_12_0_6,
  output     [2:0]    port_state_out_12_0_7,
  output     [2:0]    port_state_out_12_1_0,
  output     [2:0]    port_state_out_12_1_1,
  output     [2:0]    port_state_out_12_1_2,
  output     [2:0]    port_state_out_12_1_3,
  output     [2:0]    port_state_out_12_1_4,
  output     [2:0]    port_state_out_12_1_5,
  output     [2:0]    port_state_out_12_1_6,
  output     [2:0]    port_state_out_12_1_7,
  output     [2:0]    port_state_out_12_2_0,
  output     [2:0]    port_state_out_12_2_1,
  output     [2:0]    port_state_out_12_2_2,
  output     [2:0]    port_state_out_12_2_3,
  output     [2:0]    port_state_out_12_2_4,
  output     [2:0]    port_state_out_12_2_5,
  output     [2:0]    port_state_out_12_2_6,
  output     [2:0]    port_state_out_12_2_7,
  output     [2:0]    port_state_out_12_3_0,
  output     [2:0]    port_state_out_12_3_1,
  output     [2:0]    port_state_out_12_3_2,
  output     [2:0]    port_state_out_12_3_3,
  output     [2:0]    port_state_out_12_3_4,
  output     [2:0]    port_state_out_12_3_5,
  output     [2:0]    port_state_out_12_3_6,
  output     [2:0]    port_state_out_12_3_7,
  output     [2:0]    port_state_out_13_0_0,
  output     [2:0]    port_state_out_13_0_1,
  output     [2:0]    port_state_out_13_0_2,
  output     [2:0]    port_state_out_13_0_3,
  output     [2:0]    port_state_out_13_0_4,
  output     [2:0]    port_state_out_13_0_5,
  output     [2:0]    port_state_out_13_0_6,
  output     [2:0]    port_state_out_13_0_7,
  output     [2:0]    port_state_out_13_1_0,
  output     [2:0]    port_state_out_13_1_1,
  output     [2:0]    port_state_out_13_1_2,
  output     [2:0]    port_state_out_13_1_3,
  output     [2:0]    port_state_out_13_1_4,
  output     [2:0]    port_state_out_13_1_5,
  output     [2:0]    port_state_out_13_1_6,
  output     [2:0]    port_state_out_13_1_7,
  output     [2:0]    port_state_out_13_2_0,
  output     [2:0]    port_state_out_13_2_1,
  output     [2:0]    port_state_out_13_2_2,
  output     [2:0]    port_state_out_13_2_3,
  output     [2:0]    port_state_out_13_2_4,
  output     [2:0]    port_state_out_13_2_5,
  output     [2:0]    port_state_out_13_2_6,
  output     [2:0]    port_state_out_13_2_7,
  output     [2:0]    port_state_out_13_3_0,
  output     [2:0]    port_state_out_13_3_1,
  output     [2:0]    port_state_out_13_3_2,
  output     [2:0]    port_state_out_13_3_3,
  output     [2:0]    port_state_out_13_3_4,
  output     [2:0]    port_state_out_13_3_5,
  output     [2:0]    port_state_out_13_3_6,
  output     [2:0]    port_state_out_13_3_7,
  output     [2:0]    port_state_out_14_0_0,
  output     [2:0]    port_state_out_14_0_1,
  output     [2:0]    port_state_out_14_0_2,
  output     [2:0]    port_state_out_14_0_3,
  output     [2:0]    port_state_out_14_0_4,
  output     [2:0]    port_state_out_14_0_5,
  output     [2:0]    port_state_out_14_0_6,
  output     [2:0]    port_state_out_14_0_7,
  output     [2:0]    port_state_out_14_1_0,
  output     [2:0]    port_state_out_14_1_1,
  output     [2:0]    port_state_out_14_1_2,
  output     [2:0]    port_state_out_14_1_3,
  output     [2:0]    port_state_out_14_1_4,
  output     [2:0]    port_state_out_14_1_5,
  output     [2:0]    port_state_out_14_1_6,
  output     [2:0]    port_state_out_14_1_7,
  output     [2:0]    port_state_out_14_2_0,
  output     [2:0]    port_state_out_14_2_1,
  output     [2:0]    port_state_out_14_2_2,
  output     [2:0]    port_state_out_14_2_3,
  output     [2:0]    port_state_out_14_2_4,
  output     [2:0]    port_state_out_14_2_5,
  output     [2:0]    port_state_out_14_2_6,
  output     [2:0]    port_state_out_14_2_7,
  output     [2:0]    port_state_out_14_3_0,
  output     [2:0]    port_state_out_14_3_1,
  output     [2:0]    port_state_out_14_3_2,
  output     [2:0]    port_state_out_14_3_3,
  output     [2:0]    port_state_out_14_3_4,
  output     [2:0]    port_state_out_14_3_5,
  output     [2:0]    port_state_out_14_3_6,
  output     [2:0]    port_state_out_14_3_7,
  output     [2:0]    port_state_out_15_0_0,
  output     [2:0]    port_state_out_15_0_1,
  output     [2:0]    port_state_out_15_0_2,
  output     [2:0]    port_state_out_15_0_3,
  output     [2:0]    port_state_out_15_0_4,
  output     [2:0]    port_state_out_15_0_5,
  output     [2:0]    port_state_out_15_0_6,
  output     [2:0]    port_state_out_15_0_7,
  output     [2:0]    port_state_out_15_1_0,
  output     [2:0]    port_state_out_15_1_1,
  output     [2:0]    port_state_out_15_1_2,
  output     [2:0]    port_state_out_15_1_3,
  output     [2:0]    port_state_out_15_1_4,
  output     [2:0]    port_state_out_15_1_5,
  output     [2:0]    port_state_out_15_1_6,
  output     [2:0]    port_state_out_15_1_7,
  output     [2:0]    port_state_out_15_2_0,
  output     [2:0]    port_state_out_15_2_1,
  output     [2:0]    port_state_out_15_2_2,
  output     [2:0]    port_state_out_15_2_3,
  output     [2:0]    port_state_out_15_2_4,
  output     [2:0]    port_state_out_15_2_5,
  output     [2:0]    port_state_out_15_2_6,
  output     [2:0]    port_state_out_15_2_7,
  output     [2:0]    port_state_out_15_3_0,
  output     [2:0]    port_state_out_15_3_1,
  output     [2:0]    port_state_out_15_3_2,
  output     [2:0]    port_state_out_15_3_3,
  output     [2:0]    port_state_out_15_3_4,
  output     [2:0]    port_state_out_15_3_5,
  output     [2:0]    port_state_out_15_3_6,
  output     [2:0]    port_state_out_15_3_7
);


  assign port_state_out_0_0_0 = port_state_in_0_0_0;
  assign port_state_out_0_0_1 = port_state_in_0_0_1;
  assign port_state_out_0_0_2 = port_state_in_0_0_2;
  assign port_state_out_0_0_3 = port_state_in_0_0_3;
  assign port_state_out_0_0_4 = port_state_in_0_0_4;
  assign port_state_out_0_0_5 = port_state_in_0_0_5;
  assign port_state_out_0_0_6 = port_state_in_0_0_6;
  assign port_state_out_0_0_7 = port_state_in_0_0_7;
  assign port_state_out_0_1_0 = port_state_in_0_1_0;
  assign port_state_out_0_1_1 = port_state_in_0_1_1;
  assign port_state_out_0_1_2 = port_state_in_0_1_2;
  assign port_state_out_0_1_3 = port_state_in_0_1_3;
  assign port_state_out_0_1_4 = port_state_in_0_1_4;
  assign port_state_out_0_1_5 = port_state_in_0_1_5;
  assign port_state_out_0_1_6 = port_state_in_0_1_6;
  assign port_state_out_0_1_7 = port_state_in_0_1_7;
  assign port_state_out_0_2_0 = port_state_in_0_2_0;
  assign port_state_out_0_2_1 = port_state_in_0_2_1;
  assign port_state_out_0_2_2 = port_state_in_0_2_2;
  assign port_state_out_0_2_3 = port_state_in_0_2_3;
  assign port_state_out_0_2_4 = port_state_in_0_2_4;
  assign port_state_out_0_2_5 = port_state_in_0_2_5;
  assign port_state_out_0_2_6 = port_state_in_0_2_6;
  assign port_state_out_0_2_7 = port_state_in_0_2_7;
  assign port_state_out_0_3_0 = port_state_in_0_3_0;
  assign port_state_out_0_3_1 = port_state_in_0_3_1;
  assign port_state_out_0_3_2 = port_state_in_0_3_2;
  assign port_state_out_0_3_3 = port_state_in_0_3_3;
  assign port_state_out_0_3_4 = port_state_in_0_3_4;
  assign port_state_out_0_3_5 = port_state_in_0_3_5;
  assign port_state_out_0_3_6 = port_state_in_0_3_6;
  assign port_state_out_0_3_7 = port_state_in_0_3_7;
  assign port_state_out_1_0_0 = port_state_in_5_0_0;
  assign port_state_out_1_0_1 = port_state_in_5_0_1;
  assign port_state_out_1_0_2 = port_state_in_5_0_2;
  assign port_state_out_1_0_3 = port_state_in_5_0_3;
  assign port_state_out_1_0_4 = port_state_in_5_0_4;
  assign port_state_out_1_0_5 = port_state_in_5_0_5;
  assign port_state_out_1_0_6 = port_state_in_5_0_6;
  assign port_state_out_1_0_7 = port_state_in_5_0_7;
  assign port_state_out_1_1_0 = port_state_in_5_1_0;
  assign port_state_out_1_1_1 = port_state_in_5_1_1;
  assign port_state_out_1_1_2 = port_state_in_5_1_2;
  assign port_state_out_1_1_3 = port_state_in_5_1_3;
  assign port_state_out_1_1_4 = port_state_in_5_1_4;
  assign port_state_out_1_1_5 = port_state_in_5_1_5;
  assign port_state_out_1_1_6 = port_state_in_5_1_6;
  assign port_state_out_1_1_7 = port_state_in_5_1_7;
  assign port_state_out_1_2_0 = port_state_in_5_2_0;
  assign port_state_out_1_2_1 = port_state_in_5_2_1;
  assign port_state_out_1_2_2 = port_state_in_5_2_2;
  assign port_state_out_1_2_3 = port_state_in_5_2_3;
  assign port_state_out_1_2_4 = port_state_in_5_2_4;
  assign port_state_out_1_2_5 = port_state_in_5_2_5;
  assign port_state_out_1_2_6 = port_state_in_5_2_6;
  assign port_state_out_1_2_7 = port_state_in_5_2_7;
  assign port_state_out_1_3_0 = port_state_in_5_3_0;
  assign port_state_out_1_3_1 = port_state_in_5_3_1;
  assign port_state_out_1_3_2 = port_state_in_5_3_2;
  assign port_state_out_1_3_3 = port_state_in_5_3_3;
  assign port_state_out_1_3_4 = port_state_in_5_3_4;
  assign port_state_out_1_3_5 = port_state_in_5_3_5;
  assign port_state_out_1_3_6 = port_state_in_5_3_6;
  assign port_state_out_1_3_7 = port_state_in_5_3_7;
  assign port_state_out_2_0_0 = port_state_in_10_0_0;
  assign port_state_out_2_0_1 = port_state_in_10_0_1;
  assign port_state_out_2_0_2 = port_state_in_10_0_2;
  assign port_state_out_2_0_3 = port_state_in_10_0_3;
  assign port_state_out_2_0_4 = port_state_in_10_0_4;
  assign port_state_out_2_0_5 = port_state_in_10_0_5;
  assign port_state_out_2_0_6 = port_state_in_10_0_6;
  assign port_state_out_2_0_7 = port_state_in_10_0_7;
  assign port_state_out_2_1_0 = port_state_in_10_1_0;
  assign port_state_out_2_1_1 = port_state_in_10_1_1;
  assign port_state_out_2_1_2 = port_state_in_10_1_2;
  assign port_state_out_2_1_3 = port_state_in_10_1_3;
  assign port_state_out_2_1_4 = port_state_in_10_1_4;
  assign port_state_out_2_1_5 = port_state_in_10_1_5;
  assign port_state_out_2_1_6 = port_state_in_10_1_6;
  assign port_state_out_2_1_7 = port_state_in_10_1_7;
  assign port_state_out_2_2_0 = port_state_in_10_2_0;
  assign port_state_out_2_2_1 = port_state_in_10_2_1;
  assign port_state_out_2_2_2 = port_state_in_10_2_2;
  assign port_state_out_2_2_3 = port_state_in_10_2_3;
  assign port_state_out_2_2_4 = port_state_in_10_2_4;
  assign port_state_out_2_2_5 = port_state_in_10_2_5;
  assign port_state_out_2_2_6 = port_state_in_10_2_6;
  assign port_state_out_2_2_7 = port_state_in_10_2_7;
  assign port_state_out_2_3_0 = port_state_in_10_3_0;
  assign port_state_out_2_3_1 = port_state_in_10_3_1;
  assign port_state_out_2_3_2 = port_state_in_10_3_2;
  assign port_state_out_2_3_3 = port_state_in_10_3_3;
  assign port_state_out_2_3_4 = port_state_in_10_3_4;
  assign port_state_out_2_3_5 = port_state_in_10_3_5;
  assign port_state_out_2_3_6 = port_state_in_10_3_6;
  assign port_state_out_2_3_7 = port_state_in_10_3_7;
  assign port_state_out_3_0_0 = port_state_in_15_0_0;
  assign port_state_out_3_0_1 = port_state_in_15_0_1;
  assign port_state_out_3_0_2 = port_state_in_15_0_2;
  assign port_state_out_3_0_3 = port_state_in_15_0_3;
  assign port_state_out_3_0_4 = port_state_in_15_0_4;
  assign port_state_out_3_0_5 = port_state_in_15_0_5;
  assign port_state_out_3_0_6 = port_state_in_15_0_6;
  assign port_state_out_3_0_7 = port_state_in_15_0_7;
  assign port_state_out_3_1_0 = port_state_in_15_1_0;
  assign port_state_out_3_1_1 = port_state_in_15_1_1;
  assign port_state_out_3_1_2 = port_state_in_15_1_2;
  assign port_state_out_3_1_3 = port_state_in_15_1_3;
  assign port_state_out_3_1_4 = port_state_in_15_1_4;
  assign port_state_out_3_1_5 = port_state_in_15_1_5;
  assign port_state_out_3_1_6 = port_state_in_15_1_6;
  assign port_state_out_3_1_7 = port_state_in_15_1_7;
  assign port_state_out_3_2_0 = port_state_in_15_2_0;
  assign port_state_out_3_2_1 = port_state_in_15_2_1;
  assign port_state_out_3_2_2 = port_state_in_15_2_2;
  assign port_state_out_3_2_3 = port_state_in_15_2_3;
  assign port_state_out_3_2_4 = port_state_in_15_2_4;
  assign port_state_out_3_2_5 = port_state_in_15_2_5;
  assign port_state_out_3_2_6 = port_state_in_15_2_6;
  assign port_state_out_3_2_7 = port_state_in_15_2_7;
  assign port_state_out_3_3_0 = port_state_in_15_3_0;
  assign port_state_out_3_3_1 = port_state_in_15_3_1;
  assign port_state_out_3_3_2 = port_state_in_15_3_2;
  assign port_state_out_3_3_3 = port_state_in_15_3_3;
  assign port_state_out_3_3_4 = port_state_in_15_3_4;
  assign port_state_out_3_3_5 = port_state_in_15_3_5;
  assign port_state_out_3_3_6 = port_state_in_15_3_6;
  assign port_state_out_3_3_7 = port_state_in_15_3_7;
  assign port_state_out_4_0_0 = port_state_in_4_0_0;
  assign port_state_out_4_0_1 = port_state_in_4_0_1;
  assign port_state_out_4_0_2 = port_state_in_4_0_2;
  assign port_state_out_4_0_3 = port_state_in_4_0_3;
  assign port_state_out_4_0_4 = port_state_in_4_0_4;
  assign port_state_out_4_0_5 = port_state_in_4_0_5;
  assign port_state_out_4_0_6 = port_state_in_4_0_6;
  assign port_state_out_4_0_7 = port_state_in_4_0_7;
  assign port_state_out_4_1_0 = port_state_in_4_1_0;
  assign port_state_out_4_1_1 = port_state_in_4_1_1;
  assign port_state_out_4_1_2 = port_state_in_4_1_2;
  assign port_state_out_4_1_3 = port_state_in_4_1_3;
  assign port_state_out_4_1_4 = port_state_in_4_1_4;
  assign port_state_out_4_1_5 = port_state_in_4_1_5;
  assign port_state_out_4_1_6 = port_state_in_4_1_6;
  assign port_state_out_4_1_7 = port_state_in_4_1_7;
  assign port_state_out_4_2_0 = port_state_in_4_2_0;
  assign port_state_out_4_2_1 = port_state_in_4_2_1;
  assign port_state_out_4_2_2 = port_state_in_4_2_2;
  assign port_state_out_4_2_3 = port_state_in_4_2_3;
  assign port_state_out_4_2_4 = port_state_in_4_2_4;
  assign port_state_out_4_2_5 = port_state_in_4_2_5;
  assign port_state_out_4_2_6 = port_state_in_4_2_6;
  assign port_state_out_4_2_7 = port_state_in_4_2_7;
  assign port_state_out_4_3_0 = port_state_in_4_3_0;
  assign port_state_out_4_3_1 = port_state_in_4_3_1;
  assign port_state_out_4_3_2 = port_state_in_4_3_2;
  assign port_state_out_4_3_3 = port_state_in_4_3_3;
  assign port_state_out_4_3_4 = port_state_in_4_3_4;
  assign port_state_out_4_3_5 = port_state_in_4_3_5;
  assign port_state_out_4_3_6 = port_state_in_4_3_6;
  assign port_state_out_4_3_7 = port_state_in_4_3_7;
  assign port_state_out_5_0_0 = port_state_in_9_0_0;
  assign port_state_out_5_0_1 = port_state_in_9_0_1;
  assign port_state_out_5_0_2 = port_state_in_9_0_2;
  assign port_state_out_5_0_3 = port_state_in_9_0_3;
  assign port_state_out_5_0_4 = port_state_in_9_0_4;
  assign port_state_out_5_0_5 = port_state_in_9_0_5;
  assign port_state_out_5_0_6 = port_state_in_9_0_6;
  assign port_state_out_5_0_7 = port_state_in_9_0_7;
  assign port_state_out_5_1_0 = port_state_in_9_1_0;
  assign port_state_out_5_1_1 = port_state_in_9_1_1;
  assign port_state_out_5_1_2 = port_state_in_9_1_2;
  assign port_state_out_5_1_3 = port_state_in_9_1_3;
  assign port_state_out_5_1_4 = port_state_in_9_1_4;
  assign port_state_out_5_1_5 = port_state_in_9_1_5;
  assign port_state_out_5_1_6 = port_state_in_9_1_6;
  assign port_state_out_5_1_7 = port_state_in_9_1_7;
  assign port_state_out_5_2_0 = port_state_in_9_2_0;
  assign port_state_out_5_2_1 = port_state_in_9_2_1;
  assign port_state_out_5_2_2 = port_state_in_9_2_2;
  assign port_state_out_5_2_3 = port_state_in_9_2_3;
  assign port_state_out_5_2_4 = port_state_in_9_2_4;
  assign port_state_out_5_2_5 = port_state_in_9_2_5;
  assign port_state_out_5_2_6 = port_state_in_9_2_6;
  assign port_state_out_5_2_7 = port_state_in_9_2_7;
  assign port_state_out_5_3_0 = port_state_in_9_3_0;
  assign port_state_out_5_3_1 = port_state_in_9_3_1;
  assign port_state_out_5_3_2 = port_state_in_9_3_2;
  assign port_state_out_5_3_3 = port_state_in_9_3_3;
  assign port_state_out_5_3_4 = port_state_in_9_3_4;
  assign port_state_out_5_3_5 = port_state_in_9_3_5;
  assign port_state_out_5_3_6 = port_state_in_9_3_6;
  assign port_state_out_5_3_7 = port_state_in_9_3_7;
  assign port_state_out_6_0_0 = port_state_in_14_0_0;
  assign port_state_out_6_0_1 = port_state_in_14_0_1;
  assign port_state_out_6_0_2 = port_state_in_14_0_2;
  assign port_state_out_6_0_3 = port_state_in_14_0_3;
  assign port_state_out_6_0_4 = port_state_in_14_0_4;
  assign port_state_out_6_0_5 = port_state_in_14_0_5;
  assign port_state_out_6_0_6 = port_state_in_14_0_6;
  assign port_state_out_6_0_7 = port_state_in_14_0_7;
  assign port_state_out_6_1_0 = port_state_in_14_1_0;
  assign port_state_out_6_1_1 = port_state_in_14_1_1;
  assign port_state_out_6_1_2 = port_state_in_14_1_2;
  assign port_state_out_6_1_3 = port_state_in_14_1_3;
  assign port_state_out_6_1_4 = port_state_in_14_1_4;
  assign port_state_out_6_1_5 = port_state_in_14_1_5;
  assign port_state_out_6_1_6 = port_state_in_14_1_6;
  assign port_state_out_6_1_7 = port_state_in_14_1_7;
  assign port_state_out_6_2_0 = port_state_in_14_2_0;
  assign port_state_out_6_2_1 = port_state_in_14_2_1;
  assign port_state_out_6_2_2 = port_state_in_14_2_2;
  assign port_state_out_6_2_3 = port_state_in_14_2_3;
  assign port_state_out_6_2_4 = port_state_in_14_2_4;
  assign port_state_out_6_2_5 = port_state_in_14_2_5;
  assign port_state_out_6_2_6 = port_state_in_14_2_6;
  assign port_state_out_6_2_7 = port_state_in_14_2_7;
  assign port_state_out_6_3_0 = port_state_in_14_3_0;
  assign port_state_out_6_3_1 = port_state_in_14_3_1;
  assign port_state_out_6_3_2 = port_state_in_14_3_2;
  assign port_state_out_6_3_3 = port_state_in_14_3_3;
  assign port_state_out_6_3_4 = port_state_in_14_3_4;
  assign port_state_out_6_3_5 = port_state_in_14_3_5;
  assign port_state_out_6_3_6 = port_state_in_14_3_6;
  assign port_state_out_6_3_7 = port_state_in_14_3_7;
  assign port_state_out_7_0_0 = port_state_in_3_0_0;
  assign port_state_out_7_0_1 = port_state_in_3_0_1;
  assign port_state_out_7_0_2 = port_state_in_3_0_2;
  assign port_state_out_7_0_3 = port_state_in_3_0_3;
  assign port_state_out_7_0_4 = port_state_in_3_0_4;
  assign port_state_out_7_0_5 = port_state_in_3_0_5;
  assign port_state_out_7_0_6 = port_state_in_3_0_6;
  assign port_state_out_7_0_7 = port_state_in_3_0_7;
  assign port_state_out_7_1_0 = port_state_in_3_1_0;
  assign port_state_out_7_1_1 = port_state_in_3_1_1;
  assign port_state_out_7_1_2 = port_state_in_3_1_2;
  assign port_state_out_7_1_3 = port_state_in_3_1_3;
  assign port_state_out_7_1_4 = port_state_in_3_1_4;
  assign port_state_out_7_1_5 = port_state_in_3_1_5;
  assign port_state_out_7_1_6 = port_state_in_3_1_6;
  assign port_state_out_7_1_7 = port_state_in_3_1_7;
  assign port_state_out_7_2_0 = port_state_in_3_2_0;
  assign port_state_out_7_2_1 = port_state_in_3_2_1;
  assign port_state_out_7_2_2 = port_state_in_3_2_2;
  assign port_state_out_7_2_3 = port_state_in_3_2_3;
  assign port_state_out_7_2_4 = port_state_in_3_2_4;
  assign port_state_out_7_2_5 = port_state_in_3_2_5;
  assign port_state_out_7_2_6 = port_state_in_3_2_6;
  assign port_state_out_7_2_7 = port_state_in_3_2_7;
  assign port_state_out_7_3_0 = port_state_in_3_3_0;
  assign port_state_out_7_3_1 = port_state_in_3_3_1;
  assign port_state_out_7_3_2 = port_state_in_3_3_2;
  assign port_state_out_7_3_3 = port_state_in_3_3_3;
  assign port_state_out_7_3_4 = port_state_in_3_3_4;
  assign port_state_out_7_3_5 = port_state_in_3_3_5;
  assign port_state_out_7_3_6 = port_state_in_3_3_6;
  assign port_state_out_7_3_7 = port_state_in_3_3_7;
  assign port_state_out_8_0_0 = port_state_in_8_0_0;
  assign port_state_out_8_0_1 = port_state_in_8_0_1;
  assign port_state_out_8_0_2 = port_state_in_8_0_2;
  assign port_state_out_8_0_3 = port_state_in_8_0_3;
  assign port_state_out_8_0_4 = port_state_in_8_0_4;
  assign port_state_out_8_0_5 = port_state_in_8_0_5;
  assign port_state_out_8_0_6 = port_state_in_8_0_6;
  assign port_state_out_8_0_7 = port_state_in_8_0_7;
  assign port_state_out_8_1_0 = port_state_in_8_1_0;
  assign port_state_out_8_1_1 = port_state_in_8_1_1;
  assign port_state_out_8_1_2 = port_state_in_8_1_2;
  assign port_state_out_8_1_3 = port_state_in_8_1_3;
  assign port_state_out_8_1_4 = port_state_in_8_1_4;
  assign port_state_out_8_1_5 = port_state_in_8_1_5;
  assign port_state_out_8_1_6 = port_state_in_8_1_6;
  assign port_state_out_8_1_7 = port_state_in_8_1_7;
  assign port_state_out_8_2_0 = port_state_in_8_2_0;
  assign port_state_out_8_2_1 = port_state_in_8_2_1;
  assign port_state_out_8_2_2 = port_state_in_8_2_2;
  assign port_state_out_8_2_3 = port_state_in_8_2_3;
  assign port_state_out_8_2_4 = port_state_in_8_2_4;
  assign port_state_out_8_2_5 = port_state_in_8_2_5;
  assign port_state_out_8_2_6 = port_state_in_8_2_6;
  assign port_state_out_8_2_7 = port_state_in_8_2_7;
  assign port_state_out_8_3_0 = port_state_in_8_3_0;
  assign port_state_out_8_3_1 = port_state_in_8_3_1;
  assign port_state_out_8_3_2 = port_state_in_8_3_2;
  assign port_state_out_8_3_3 = port_state_in_8_3_3;
  assign port_state_out_8_3_4 = port_state_in_8_3_4;
  assign port_state_out_8_3_5 = port_state_in_8_3_5;
  assign port_state_out_8_3_6 = port_state_in_8_3_6;
  assign port_state_out_8_3_7 = port_state_in_8_3_7;
  assign port_state_out_9_0_0 = port_state_in_13_0_0;
  assign port_state_out_9_0_1 = port_state_in_13_0_1;
  assign port_state_out_9_0_2 = port_state_in_13_0_2;
  assign port_state_out_9_0_3 = port_state_in_13_0_3;
  assign port_state_out_9_0_4 = port_state_in_13_0_4;
  assign port_state_out_9_0_5 = port_state_in_13_0_5;
  assign port_state_out_9_0_6 = port_state_in_13_0_6;
  assign port_state_out_9_0_7 = port_state_in_13_0_7;
  assign port_state_out_9_1_0 = port_state_in_13_1_0;
  assign port_state_out_9_1_1 = port_state_in_13_1_1;
  assign port_state_out_9_1_2 = port_state_in_13_1_2;
  assign port_state_out_9_1_3 = port_state_in_13_1_3;
  assign port_state_out_9_1_4 = port_state_in_13_1_4;
  assign port_state_out_9_1_5 = port_state_in_13_1_5;
  assign port_state_out_9_1_6 = port_state_in_13_1_6;
  assign port_state_out_9_1_7 = port_state_in_13_1_7;
  assign port_state_out_9_2_0 = port_state_in_13_2_0;
  assign port_state_out_9_2_1 = port_state_in_13_2_1;
  assign port_state_out_9_2_2 = port_state_in_13_2_2;
  assign port_state_out_9_2_3 = port_state_in_13_2_3;
  assign port_state_out_9_2_4 = port_state_in_13_2_4;
  assign port_state_out_9_2_5 = port_state_in_13_2_5;
  assign port_state_out_9_2_6 = port_state_in_13_2_6;
  assign port_state_out_9_2_7 = port_state_in_13_2_7;
  assign port_state_out_9_3_0 = port_state_in_13_3_0;
  assign port_state_out_9_3_1 = port_state_in_13_3_1;
  assign port_state_out_9_3_2 = port_state_in_13_3_2;
  assign port_state_out_9_3_3 = port_state_in_13_3_3;
  assign port_state_out_9_3_4 = port_state_in_13_3_4;
  assign port_state_out_9_3_5 = port_state_in_13_3_5;
  assign port_state_out_9_3_6 = port_state_in_13_3_6;
  assign port_state_out_9_3_7 = port_state_in_13_3_7;
  assign port_state_out_10_0_0 = port_state_in_2_0_0;
  assign port_state_out_10_0_1 = port_state_in_2_0_1;
  assign port_state_out_10_0_2 = port_state_in_2_0_2;
  assign port_state_out_10_0_3 = port_state_in_2_0_3;
  assign port_state_out_10_0_4 = port_state_in_2_0_4;
  assign port_state_out_10_0_5 = port_state_in_2_0_5;
  assign port_state_out_10_0_6 = port_state_in_2_0_6;
  assign port_state_out_10_0_7 = port_state_in_2_0_7;
  assign port_state_out_10_1_0 = port_state_in_2_1_0;
  assign port_state_out_10_1_1 = port_state_in_2_1_1;
  assign port_state_out_10_1_2 = port_state_in_2_1_2;
  assign port_state_out_10_1_3 = port_state_in_2_1_3;
  assign port_state_out_10_1_4 = port_state_in_2_1_4;
  assign port_state_out_10_1_5 = port_state_in_2_1_5;
  assign port_state_out_10_1_6 = port_state_in_2_1_6;
  assign port_state_out_10_1_7 = port_state_in_2_1_7;
  assign port_state_out_10_2_0 = port_state_in_2_2_0;
  assign port_state_out_10_2_1 = port_state_in_2_2_1;
  assign port_state_out_10_2_2 = port_state_in_2_2_2;
  assign port_state_out_10_2_3 = port_state_in_2_2_3;
  assign port_state_out_10_2_4 = port_state_in_2_2_4;
  assign port_state_out_10_2_5 = port_state_in_2_2_5;
  assign port_state_out_10_2_6 = port_state_in_2_2_6;
  assign port_state_out_10_2_7 = port_state_in_2_2_7;
  assign port_state_out_10_3_0 = port_state_in_2_3_0;
  assign port_state_out_10_3_1 = port_state_in_2_3_1;
  assign port_state_out_10_3_2 = port_state_in_2_3_2;
  assign port_state_out_10_3_3 = port_state_in_2_3_3;
  assign port_state_out_10_3_4 = port_state_in_2_3_4;
  assign port_state_out_10_3_5 = port_state_in_2_3_5;
  assign port_state_out_10_3_6 = port_state_in_2_3_6;
  assign port_state_out_10_3_7 = port_state_in_2_3_7;
  assign port_state_out_11_0_0 = port_state_in_7_0_0;
  assign port_state_out_11_0_1 = port_state_in_7_0_1;
  assign port_state_out_11_0_2 = port_state_in_7_0_2;
  assign port_state_out_11_0_3 = port_state_in_7_0_3;
  assign port_state_out_11_0_4 = port_state_in_7_0_4;
  assign port_state_out_11_0_5 = port_state_in_7_0_5;
  assign port_state_out_11_0_6 = port_state_in_7_0_6;
  assign port_state_out_11_0_7 = port_state_in_7_0_7;
  assign port_state_out_11_1_0 = port_state_in_7_1_0;
  assign port_state_out_11_1_1 = port_state_in_7_1_1;
  assign port_state_out_11_1_2 = port_state_in_7_1_2;
  assign port_state_out_11_1_3 = port_state_in_7_1_3;
  assign port_state_out_11_1_4 = port_state_in_7_1_4;
  assign port_state_out_11_1_5 = port_state_in_7_1_5;
  assign port_state_out_11_1_6 = port_state_in_7_1_6;
  assign port_state_out_11_1_7 = port_state_in_7_1_7;
  assign port_state_out_11_2_0 = port_state_in_7_2_0;
  assign port_state_out_11_2_1 = port_state_in_7_2_1;
  assign port_state_out_11_2_2 = port_state_in_7_2_2;
  assign port_state_out_11_2_3 = port_state_in_7_2_3;
  assign port_state_out_11_2_4 = port_state_in_7_2_4;
  assign port_state_out_11_2_5 = port_state_in_7_2_5;
  assign port_state_out_11_2_6 = port_state_in_7_2_6;
  assign port_state_out_11_2_7 = port_state_in_7_2_7;
  assign port_state_out_11_3_0 = port_state_in_7_3_0;
  assign port_state_out_11_3_1 = port_state_in_7_3_1;
  assign port_state_out_11_3_2 = port_state_in_7_3_2;
  assign port_state_out_11_3_3 = port_state_in_7_3_3;
  assign port_state_out_11_3_4 = port_state_in_7_3_4;
  assign port_state_out_11_3_5 = port_state_in_7_3_5;
  assign port_state_out_11_3_6 = port_state_in_7_3_6;
  assign port_state_out_11_3_7 = port_state_in_7_3_7;
  assign port_state_out_12_0_0 = port_state_in_12_0_0;
  assign port_state_out_12_0_1 = port_state_in_12_0_1;
  assign port_state_out_12_0_2 = port_state_in_12_0_2;
  assign port_state_out_12_0_3 = port_state_in_12_0_3;
  assign port_state_out_12_0_4 = port_state_in_12_0_4;
  assign port_state_out_12_0_5 = port_state_in_12_0_5;
  assign port_state_out_12_0_6 = port_state_in_12_0_6;
  assign port_state_out_12_0_7 = port_state_in_12_0_7;
  assign port_state_out_12_1_0 = port_state_in_12_1_0;
  assign port_state_out_12_1_1 = port_state_in_12_1_1;
  assign port_state_out_12_1_2 = port_state_in_12_1_2;
  assign port_state_out_12_1_3 = port_state_in_12_1_3;
  assign port_state_out_12_1_4 = port_state_in_12_1_4;
  assign port_state_out_12_1_5 = port_state_in_12_1_5;
  assign port_state_out_12_1_6 = port_state_in_12_1_6;
  assign port_state_out_12_1_7 = port_state_in_12_1_7;
  assign port_state_out_12_2_0 = port_state_in_12_2_0;
  assign port_state_out_12_2_1 = port_state_in_12_2_1;
  assign port_state_out_12_2_2 = port_state_in_12_2_2;
  assign port_state_out_12_2_3 = port_state_in_12_2_3;
  assign port_state_out_12_2_4 = port_state_in_12_2_4;
  assign port_state_out_12_2_5 = port_state_in_12_2_5;
  assign port_state_out_12_2_6 = port_state_in_12_2_6;
  assign port_state_out_12_2_7 = port_state_in_12_2_7;
  assign port_state_out_12_3_0 = port_state_in_12_3_0;
  assign port_state_out_12_3_1 = port_state_in_12_3_1;
  assign port_state_out_12_3_2 = port_state_in_12_3_2;
  assign port_state_out_12_3_3 = port_state_in_12_3_3;
  assign port_state_out_12_3_4 = port_state_in_12_3_4;
  assign port_state_out_12_3_5 = port_state_in_12_3_5;
  assign port_state_out_12_3_6 = port_state_in_12_3_6;
  assign port_state_out_12_3_7 = port_state_in_12_3_7;
  assign port_state_out_13_0_0 = port_state_in_1_0_0;
  assign port_state_out_13_0_1 = port_state_in_1_0_1;
  assign port_state_out_13_0_2 = port_state_in_1_0_2;
  assign port_state_out_13_0_3 = port_state_in_1_0_3;
  assign port_state_out_13_0_4 = port_state_in_1_0_4;
  assign port_state_out_13_0_5 = port_state_in_1_0_5;
  assign port_state_out_13_0_6 = port_state_in_1_0_6;
  assign port_state_out_13_0_7 = port_state_in_1_0_7;
  assign port_state_out_13_1_0 = port_state_in_1_1_0;
  assign port_state_out_13_1_1 = port_state_in_1_1_1;
  assign port_state_out_13_1_2 = port_state_in_1_1_2;
  assign port_state_out_13_1_3 = port_state_in_1_1_3;
  assign port_state_out_13_1_4 = port_state_in_1_1_4;
  assign port_state_out_13_1_5 = port_state_in_1_1_5;
  assign port_state_out_13_1_6 = port_state_in_1_1_6;
  assign port_state_out_13_1_7 = port_state_in_1_1_7;
  assign port_state_out_13_2_0 = port_state_in_1_2_0;
  assign port_state_out_13_2_1 = port_state_in_1_2_1;
  assign port_state_out_13_2_2 = port_state_in_1_2_2;
  assign port_state_out_13_2_3 = port_state_in_1_2_3;
  assign port_state_out_13_2_4 = port_state_in_1_2_4;
  assign port_state_out_13_2_5 = port_state_in_1_2_5;
  assign port_state_out_13_2_6 = port_state_in_1_2_6;
  assign port_state_out_13_2_7 = port_state_in_1_2_7;
  assign port_state_out_13_3_0 = port_state_in_1_3_0;
  assign port_state_out_13_3_1 = port_state_in_1_3_1;
  assign port_state_out_13_3_2 = port_state_in_1_3_2;
  assign port_state_out_13_3_3 = port_state_in_1_3_3;
  assign port_state_out_13_3_4 = port_state_in_1_3_4;
  assign port_state_out_13_3_5 = port_state_in_1_3_5;
  assign port_state_out_13_3_6 = port_state_in_1_3_6;
  assign port_state_out_13_3_7 = port_state_in_1_3_7;
  assign port_state_out_14_0_0 = port_state_in_6_0_0;
  assign port_state_out_14_0_1 = port_state_in_6_0_1;
  assign port_state_out_14_0_2 = port_state_in_6_0_2;
  assign port_state_out_14_0_3 = port_state_in_6_0_3;
  assign port_state_out_14_0_4 = port_state_in_6_0_4;
  assign port_state_out_14_0_5 = port_state_in_6_0_5;
  assign port_state_out_14_0_6 = port_state_in_6_0_6;
  assign port_state_out_14_0_7 = port_state_in_6_0_7;
  assign port_state_out_14_1_0 = port_state_in_6_1_0;
  assign port_state_out_14_1_1 = port_state_in_6_1_1;
  assign port_state_out_14_1_2 = port_state_in_6_1_2;
  assign port_state_out_14_1_3 = port_state_in_6_1_3;
  assign port_state_out_14_1_4 = port_state_in_6_1_4;
  assign port_state_out_14_1_5 = port_state_in_6_1_5;
  assign port_state_out_14_1_6 = port_state_in_6_1_6;
  assign port_state_out_14_1_7 = port_state_in_6_1_7;
  assign port_state_out_14_2_0 = port_state_in_6_2_0;
  assign port_state_out_14_2_1 = port_state_in_6_2_1;
  assign port_state_out_14_2_2 = port_state_in_6_2_2;
  assign port_state_out_14_2_3 = port_state_in_6_2_3;
  assign port_state_out_14_2_4 = port_state_in_6_2_4;
  assign port_state_out_14_2_5 = port_state_in_6_2_5;
  assign port_state_out_14_2_6 = port_state_in_6_2_6;
  assign port_state_out_14_2_7 = port_state_in_6_2_7;
  assign port_state_out_14_3_0 = port_state_in_6_3_0;
  assign port_state_out_14_3_1 = port_state_in_6_3_1;
  assign port_state_out_14_3_2 = port_state_in_6_3_2;
  assign port_state_out_14_3_3 = port_state_in_6_3_3;
  assign port_state_out_14_3_4 = port_state_in_6_3_4;
  assign port_state_out_14_3_5 = port_state_in_6_3_5;
  assign port_state_out_14_3_6 = port_state_in_6_3_6;
  assign port_state_out_14_3_7 = port_state_in_6_3_7;
  assign port_state_out_15_0_0 = port_state_in_11_0_0;
  assign port_state_out_15_0_1 = port_state_in_11_0_1;
  assign port_state_out_15_0_2 = port_state_in_11_0_2;
  assign port_state_out_15_0_3 = port_state_in_11_0_3;
  assign port_state_out_15_0_4 = port_state_in_11_0_4;
  assign port_state_out_15_0_5 = port_state_in_11_0_5;
  assign port_state_out_15_0_6 = port_state_in_11_0_6;
  assign port_state_out_15_0_7 = port_state_in_11_0_7;
  assign port_state_out_15_1_0 = port_state_in_11_1_0;
  assign port_state_out_15_1_1 = port_state_in_11_1_1;
  assign port_state_out_15_1_2 = port_state_in_11_1_2;
  assign port_state_out_15_1_3 = port_state_in_11_1_3;
  assign port_state_out_15_1_4 = port_state_in_11_1_4;
  assign port_state_out_15_1_5 = port_state_in_11_1_5;
  assign port_state_out_15_1_6 = port_state_in_11_1_6;
  assign port_state_out_15_1_7 = port_state_in_11_1_7;
  assign port_state_out_15_2_0 = port_state_in_11_2_0;
  assign port_state_out_15_2_1 = port_state_in_11_2_1;
  assign port_state_out_15_2_2 = port_state_in_11_2_2;
  assign port_state_out_15_2_3 = port_state_in_11_2_3;
  assign port_state_out_15_2_4 = port_state_in_11_2_4;
  assign port_state_out_15_2_5 = port_state_in_11_2_5;
  assign port_state_out_15_2_6 = port_state_in_11_2_6;
  assign port_state_out_15_2_7 = port_state_in_11_2_7;
  assign port_state_out_15_3_0 = port_state_in_11_3_0;
  assign port_state_out_15_3_1 = port_state_in_11_3_1;
  assign port_state_out_15_3_2 = port_state_in_11_3_2;
  assign port_state_out_15_3_3 = port_state_in_11_3_3;
  assign port_state_out_15_3_4 = port_state_in_11_3_4;
  assign port_state_out_15_3_5 = port_state_in_11_3_5;
  assign port_state_out_15_3_6 = port_state_in_11_3_6;
  assign port_state_out_15_3_7 = port_state_in_11_3_7;

endmodule

//Sbox_AES_BoyarPeralta replaced by Sbox_AES_BoyarPeralta

//Sbox_AES_BoyarPeralta replaced by Sbox_AES_BoyarPeralta

//Sbox_AES_BoyarPeralta replaced by Sbox_AES_BoyarPeralta

//Sbox_AES_BoyarPeralta replaced by Sbox_AES_BoyarPeralta

//Sbox_AES_BoyarPeralta replaced by Sbox_AES_BoyarPeralta

//Sbox_AES_BoyarPeralta replaced by Sbox_AES_BoyarPeralta

//Sbox_AES_BoyarPeralta replaced by Sbox_AES_BoyarPeralta

//Sbox_AES_BoyarPeralta replaced by Sbox_AES_BoyarPeralta

//Sbox_AES_BoyarPeralta replaced by Sbox_AES_BoyarPeralta

//Sbox_AES_BoyarPeralta replaced by Sbox_AES_BoyarPeralta

//Sbox_AES_BoyarPeralta replaced by Sbox_AES_BoyarPeralta

//Sbox_AES_BoyarPeralta replaced by Sbox_AES_BoyarPeralta

//Sbox_AES_BoyarPeralta replaced by Sbox_AES_BoyarPeralta

//Sbox_AES_BoyarPeralta replaced by Sbox_AES_BoyarPeralta

//Sbox_AES_BoyarPeralta replaced by Sbox_AES_BoyarPeralta

module Sbox_AES_BoyarPeralta (
  input      [2:0]    port_i_0_0,
  input      [2:0]    port_i_0_1,
  input      [2:0]    port_i_0_2,
  input      [2:0]    port_i_0_3,
  input      [2:0]    port_i_0_4,
  input      [2:0]    port_i_0_5,
  input      [2:0]    port_i_0_6,
  input      [2:0]    port_i_0_7,
  input      [2:0]    port_i_1_0,
  input      [2:0]    port_i_1_1,
  input      [2:0]    port_i_1_2,
  input      [2:0]    port_i_1_3,
  input      [2:0]    port_i_1_4,
  input      [2:0]    port_i_1_5,
  input      [2:0]    port_i_1_6,
  input      [2:0]    port_i_1_7,
  input      [2:0]    port_i_2_0,
  input      [2:0]    port_i_2_1,
  input      [2:0]    port_i_2_2,
  input      [2:0]    port_i_2_3,
  input      [2:0]    port_i_2_4,
  input      [2:0]    port_i_2_5,
  input      [2:0]    port_i_2_6,
  input      [2:0]    port_i_2_7,
  input      [2:0]    port_i_3_0,
  input      [2:0]    port_i_3_1,
  input      [2:0]    port_i_3_2,
  input      [2:0]    port_i_3_3,
  input      [2:0]    port_i_3_4,
  input      [2:0]    port_i_3_5,
  input      [2:0]    port_i_3_6,
  input      [2:0]    port_i_3_7,
  output     [2:0]    port_o_0_0,
  output     [2:0]    port_o_0_1,
  output     [2:0]    port_o_0_2,
  output     [2:0]    port_o_0_3,
  output     [2:0]    port_o_0_4,
  output     [2:0]    port_o_0_5,
  output     [2:0]    port_o_0_6,
  output     [2:0]    port_o_0_7,
  output     [2:0]    port_o_1_0,
  output     [2:0]    port_o_1_1,
  output     [2:0]    port_o_1_2,
  output     [2:0]    port_o_1_3,
  output     [2:0]    port_o_1_4,
  output     [2:0]    port_o_1_5,
  output     [2:0]    port_o_1_6,
  output     [2:0]    port_o_1_7,
  output     [2:0]    port_o_2_0,
  output     [2:0]    port_o_2_1,
  output     [2:0]    port_o_2_2,
  output     [2:0]    port_o_2_3,
  output     [2:0]    port_o_2_4,
  output     [2:0]    port_o_2_5,
  output     [2:0]    port_o_2_6,
  output     [2:0]    port_o_2_7,
  output     [2:0]    port_o_3_0,
  output     [2:0]    port_o_3_1,
  output     [2:0]    port_o_3_2,
  output     [2:0]    port_o_3_3,
  output     [2:0]    port_o_3_4,
  output     [2:0]    port_o_3_5,
  output     [2:0]    port_o_3_6,
  output     [2:0]    port_o_3_7,
  input               clk,
  input               reset
);

  wire       [2:0]    t1_xor_port_y_0;
  wire       [2:0]    t1_xor_port_y_1;
  wire       [2:0]    t1_xor_port_y_2;
  wire       [2:0]    t1_xor_port_y_3;
  wire       [2:0]    t2_xor_port_y_0;
  wire       [2:0]    t2_xor_port_y_1;
  wire       [2:0]    t2_xor_port_y_2;
  wire       [2:0]    t2_xor_port_y_3;
  wire       [2:0]    t3_xor_port_y_0;
  wire       [2:0]    t3_xor_port_y_1;
  wire       [2:0]    t3_xor_port_y_2;
  wire       [2:0]    t3_xor_port_y_3;
  wire       [2:0]    t4_xor_port_y_0;
  wire       [2:0]    t4_xor_port_y_1;
  wire       [2:0]    t4_xor_port_y_2;
  wire       [2:0]    t4_xor_port_y_3;
  wire       [2:0]    t5_xor_port_y_0;
  wire       [2:0]    t5_xor_port_y_1;
  wire       [2:0]    t5_xor_port_y_2;
  wire       [2:0]    t5_xor_port_y_3;
  wire       [2:0]    t6_xor_port_y_0;
  wire       [2:0]    t6_xor_port_y_1;
  wire       [2:0]    t6_xor_port_y_2;
  wire       [2:0]    t6_xor_port_y_3;
  wire       [2:0]    t7_xor_port_y_0;
  wire       [2:0]    t7_xor_port_y_1;
  wire       [2:0]    t7_xor_port_y_2;
  wire       [2:0]    t7_xor_port_y_3;
  wire       [2:0]    t8_xor_port_y_0;
  wire       [2:0]    t8_xor_port_y_1;
  wire       [2:0]    t8_xor_port_y_2;
  wire       [2:0]    t8_xor_port_y_3;
  wire       [2:0]    t9_xor_port_y_0;
  wire       [2:0]    t9_xor_port_y_1;
  wire       [2:0]    t9_xor_port_y_2;
  wire       [2:0]    t9_xor_port_y_3;
  wire       [2:0]    t10_xor_port_y_0;
  wire       [2:0]    t10_xor_port_y_1;
  wire       [2:0]    t10_xor_port_y_2;
  wire       [2:0]    t10_xor_port_y_3;
  wire       [2:0]    t11_xor_port_y_0;
  wire       [2:0]    t11_xor_port_y_1;
  wire       [2:0]    t11_xor_port_y_2;
  wire       [2:0]    t11_xor_port_y_3;
  wire       [2:0]    t12_xor_port_y_0;
  wire       [2:0]    t12_xor_port_y_1;
  wire       [2:0]    t12_xor_port_y_2;
  wire       [2:0]    t12_xor_port_y_3;
  wire       [2:0]    t13_xor_port_y_0;
  wire       [2:0]    t13_xor_port_y_1;
  wire       [2:0]    t13_xor_port_y_2;
  wire       [2:0]    t13_xor_port_y_3;
  wire       [2:0]    t14_xor_port_y_0;
  wire       [2:0]    t14_xor_port_y_1;
  wire       [2:0]    t14_xor_port_y_2;
  wire       [2:0]    t14_xor_port_y_3;
  wire       [2:0]    t15_xor_port_y_0;
  wire       [2:0]    t15_xor_port_y_1;
  wire       [2:0]    t15_xor_port_y_2;
  wire       [2:0]    t15_xor_port_y_3;
  wire       [2:0]    t16_xor_port_y_0;
  wire       [2:0]    t16_xor_port_y_1;
  wire       [2:0]    t16_xor_port_y_2;
  wire       [2:0]    t16_xor_port_y_3;
  wire       [2:0]    t17_xor_port_y_0;
  wire       [2:0]    t17_xor_port_y_1;
  wire       [2:0]    t17_xor_port_y_2;
  wire       [2:0]    t17_xor_port_y_3;
  wire       [2:0]    t18_xor_port_y_0;
  wire       [2:0]    t18_xor_port_y_1;
  wire       [2:0]    t18_xor_port_y_2;
  wire       [2:0]    t18_xor_port_y_3;
  wire       [2:0]    t19_xor_port_y_0;
  wire       [2:0]    t19_xor_port_y_1;
  wire       [2:0]    t19_xor_port_y_2;
  wire       [2:0]    t19_xor_port_y_3;
  wire       [2:0]    t20_xor_port_y_0;
  wire       [2:0]    t20_xor_port_y_1;
  wire       [2:0]    t20_xor_port_y_2;
  wire       [2:0]    t20_xor_port_y_3;
  wire       [2:0]    t21_xor_port_y_0;
  wire       [2:0]    t21_xor_port_y_1;
  wire       [2:0]    t21_xor_port_y_2;
  wire       [2:0]    t21_xor_port_y_3;
  wire       [2:0]    t22_xor_port_y_0;
  wire       [2:0]    t22_xor_port_y_1;
  wire       [2:0]    t22_xor_port_y_2;
  wire       [2:0]    t22_xor_port_y_3;
  wire       [2:0]    t23_xor_port_y_0;
  wire       [2:0]    t23_xor_port_y_1;
  wire       [2:0]    t23_xor_port_y_2;
  wire       [2:0]    t23_xor_port_y_3;
  wire       [2:0]    t24_xor_port_y_0;
  wire       [2:0]    t24_xor_port_y_1;
  wire       [2:0]    t24_xor_port_y_2;
  wire       [2:0]    t24_xor_port_y_3;
  wire       [2:0]    t25_xor_port_y_0;
  wire       [2:0]    t25_xor_port_y_1;
  wire       [2:0]    t25_xor_port_y_2;
  wire       [2:0]    t25_xor_port_y_3;
  wire       [2:0]    t26_xor_port_y_0;
  wire       [2:0]    t26_xor_port_y_1;
  wire       [2:0]    t26_xor_port_y_2;
  wire       [2:0]    t26_xor_port_y_3;
  wire       [2:0]    t27_xor_port_y_0;
  wire       [2:0]    t27_xor_port_y_1;
  wire       [2:0]    t27_xor_port_y_2;
  wire       [2:0]    t27_xor_port_y_3;
  wire       [2:0]    m1_port_y_0;
  wire       [2:0]    m1_port_y_1;
  wire       [2:0]    m1_port_y_2;
  wire       [2:0]    m1_port_y_3;
  wire       [2:0]    m2_port_y_0;
  wire       [2:0]    m2_port_y_1;
  wire       [2:0]    m2_port_y_2;
  wire       [2:0]    m2_port_y_3;
  wire       [2:0]    m4_port_y_0;
  wire       [2:0]    m4_port_y_1;
  wire       [2:0]    m4_port_y_2;
  wire       [2:0]    m4_port_y_3;
  wire       [2:0]    m6_port_y_0;
  wire       [2:0]    m6_port_y_1;
  wire       [2:0]    m6_port_y_2;
  wire       [2:0]    m6_port_y_3;
  wire       [2:0]    m7_port_y_0;
  wire       [2:0]    m7_port_y_1;
  wire       [2:0]    m7_port_y_2;
  wire       [2:0]    m7_port_y_3;
  wire       [2:0]    m9_port_y_0;
  wire       [2:0]    m9_port_y_1;
  wire       [2:0]    m9_port_y_2;
  wire       [2:0]    m9_port_y_3;
  wire       [2:0]    m11_port_y_0;
  wire       [2:0]    m11_port_y_1;
  wire       [2:0]    m11_port_y_2;
  wire       [2:0]    m11_port_y_3;
  wire       [2:0]    m12_port_y_0;
  wire       [2:0]    m12_port_y_1;
  wire       [2:0]    m12_port_y_2;
  wire       [2:0]    m12_port_y_3;
  wire       [2:0]    m14_port_y_0;
  wire       [2:0]    m14_port_y_1;
  wire       [2:0]    m14_port_y_2;
  wire       [2:0]    m14_port_y_3;
  wire       [2:0]    m3_xor_port_y_0;
  wire       [2:0]    m3_xor_port_y_1;
  wire       [2:0]    m3_xor_port_y_2;
  wire       [2:0]    m3_xor_port_y_3;
  wire       [2:0]    m5_xor_port_y_0;
  wire       [2:0]    m5_xor_port_y_1;
  wire       [2:0]    m5_xor_port_y_2;
  wire       [2:0]    m5_xor_port_y_3;
  wire       [2:0]    m8_xor_port_y_0;
  wire       [2:0]    m8_xor_port_y_1;
  wire       [2:0]    m8_xor_port_y_2;
  wire       [2:0]    m8_xor_port_y_3;
  wire       [2:0]    m10_xor_port_y_0;
  wire       [2:0]    m10_xor_port_y_1;
  wire       [2:0]    m10_xor_port_y_2;
  wire       [2:0]    m10_xor_port_y_3;
  wire       [2:0]    m13_xor_port_y_0;
  wire       [2:0]    m13_xor_port_y_1;
  wire       [2:0]    m13_xor_port_y_2;
  wire       [2:0]    m13_xor_port_y_3;
  wire       [2:0]    m15_xor_port_y_0;
  wire       [2:0]    m15_xor_port_y_1;
  wire       [2:0]    m15_xor_port_y_2;
  wire       [2:0]    m15_xor_port_y_3;
  wire       [2:0]    m16_xor_port_y_0;
  wire       [2:0]    m16_xor_port_y_1;
  wire       [2:0]    m16_xor_port_y_2;
  wire       [2:0]    m16_xor_port_y_3;
  wire       [2:0]    m17_xor_port_y_0;
  wire       [2:0]    m17_xor_port_y_1;
  wire       [2:0]    m17_xor_port_y_2;
  wire       [2:0]    m17_xor_port_y_3;
  wire       [2:0]    m18_xor_port_y_0;
  wire       [2:0]    m18_xor_port_y_1;
  wire       [2:0]    m18_xor_port_y_2;
  wire       [2:0]    m18_xor_port_y_3;
  wire       [2:0]    m19_xor_port_y_0;
  wire       [2:0]    m19_xor_port_y_1;
  wire       [2:0]    m19_xor_port_y_2;
  wire       [2:0]    m19_xor_port_y_3;
  wire       [2:0]    m20_xor_port_y_0;
  wire       [2:0]    m20_xor_port_y_1;
  wire       [2:0]    m20_xor_port_y_2;
  wire       [2:0]    m20_xor_port_y_3;
  wire       [2:0]    m21_xor_port_y_0;
  wire       [2:0]    m21_xor_port_y_1;
  wire       [2:0]    m21_xor_port_y_2;
  wire       [2:0]    m21_xor_port_y_3;
  wire       [2:0]    m22_xor_port_y_0;
  wire       [2:0]    m22_xor_port_y_1;
  wire       [2:0]    m22_xor_port_y_2;
  wire       [2:0]    m22_xor_port_y_3;
  wire       [2:0]    m23_xor_port_y_0;
  wire       [2:0]    m23_xor_port_y_1;
  wire       [2:0]    m23_xor_port_y_2;
  wire       [2:0]    m23_xor_port_y_3;
  wire       [2:0]    m24_xor_port_y_0;
  wire       [2:0]    m24_xor_port_y_1;
  wire       [2:0]    m24_xor_port_y_2;
  wire       [2:0]    m24_xor_port_y_3;
  wire       [2:0]    m25_port_y_0;
  wire       [2:0]    m25_port_y_1;
  wire       [2:0]    m25_port_y_2;
  wire       [2:0]    m25_port_y_3;
  wire       [2:0]    m27_xor_port_y_0;
  wire       [2:0]    m27_xor_port_y_1;
  wire       [2:0]    m27_xor_port_y_2;
  wire       [2:0]    m27_xor_port_y_3;
  wire       [2:0]    m31_port_y_0;
  wire       [2:0]    m31_port_y_1;
  wire       [2:0]    m31_port_y_2;
  wire       [2:0]    m31_port_y_3;
  wire       [2:0]    m34_port_y_0;
  wire       [2:0]    m34_port_y_1;
  wire       [2:0]    m34_port_y_2;
  wire       [2:0]    m34_port_y_3;
  wire       [2:0]    m26_xor_port_y_0;
  wire       [2:0]    m26_xor_port_y_1;
  wire       [2:0]    m26_xor_port_y_2;
  wire       [2:0]    m26_xor_port_y_3;
  wire       [2:0]    m28_xor_port_y_0;
  wire       [2:0]    m28_xor_port_y_1;
  wire       [2:0]    m28_xor_port_y_2;
  wire       [2:0]    m28_xor_port_y_3;
  wire       [2:0]    m29_port_y_0;
  wire       [2:0]    m29_port_y_1;
  wire       [2:0]    m29_port_y_2;
  wire       [2:0]    m29_port_y_3;
  wire       [2:0]    m30_port_y_0;
  wire       [2:0]    m30_port_y_1;
  wire       [2:0]    m30_port_y_2;
  wire       [2:0]    m30_port_y_3;
  wire       [2:0]    m32_port_y_0;
  wire       [2:0]    m32_port_y_1;
  wire       [2:0]    m32_port_y_2;
  wire       [2:0]    m32_port_y_3;
  wire       [2:0]    m33_xor_port_y_0;
  wire       [2:0]    m33_xor_port_y_1;
  wire       [2:0]    m33_xor_port_y_2;
  wire       [2:0]    m33_xor_port_y_3;
  wire       [2:0]    m35_port_y_0;
  wire       [2:0]    m35_port_y_1;
  wire       [2:0]    m35_port_y_2;
  wire       [2:0]    m35_port_y_3;
  wire       [2:0]    m36_xor_port_y_0;
  wire       [2:0]    m36_xor_port_y_1;
  wire       [2:0]    m36_xor_port_y_2;
  wire       [2:0]    m36_xor_port_y_3;
  wire       [2:0]    m37_xor_port_y_0;
  wire       [2:0]    m37_xor_port_y_1;
  wire       [2:0]    m37_xor_port_y_2;
  wire       [2:0]    m37_xor_port_y_3;
  wire       [2:0]    m38_xor_port_y_0;
  wire       [2:0]    m38_xor_port_y_1;
  wire       [2:0]    m38_xor_port_y_2;
  wire       [2:0]    m38_xor_port_y_3;
  wire       [2:0]    m39_xor_port_y_0;
  wire       [2:0]    m39_xor_port_y_1;
  wire       [2:0]    m39_xor_port_y_2;
  wire       [2:0]    m39_xor_port_y_3;
  wire       [2:0]    m40_xor_port_y_0;
  wire       [2:0]    m40_xor_port_y_1;
  wire       [2:0]    m40_xor_port_y_2;
  wire       [2:0]    m40_xor_port_y_3;
  wire       [2:0]    m41_xor_port_y_0;
  wire       [2:0]    m41_xor_port_y_1;
  wire       [2:0]    m41_xor_port_y_2;
  wire       [2:0]    m41_xor_port_y_3;
  wire       [2:0]    m42_xor_port_y_0;
  wire       [2:0]    m42_xor_port_y_1;
  wire       [2:0]    m42_xor_port_y_2;
  wire       [2:0]    m42_xor_port_y_3;
  wire       [2:0]    m43_xor_port_y_0;
  wire       [2:0]    m43_xor_port_y_1;
  wire       [2:0]    m43_xor_port_y_2;
  wire       [2:0]    m43_xor_port_y_3;
  wire       [2:0]    m44_xor_port_y_0;
  wire       [2:0]    m44_xor_port_y_1;
  wire       [2:0]    m44_xor_port_y_2;
  wire       [2:0]    m44_xor_port_y_3;
  wire       [2:0]    m45_xor_port_y_0;
  wire       [2:0]    m45_xor_port_y_1;
  wire       [2:0]    m45_xor_port_y_2;
  wire       [2:0]    m45_xor_port_y_3;
  wire       [2:0]    m46_mul_port_y_0;
  wire       [2:0]    m46_mul_port_y_1;
  wire       [2:0]    m46_mul_port_y_2;
  wire       [2:0]    m46_mul_port_y_3;
  wire       [2:0]    m47_mul_port_y_0;
  wire       [2:0]    m47_mul_port_y_1;
  wire       [2:0]    m47_mul_port_y_2;
  wire       [2:0]    m47_mul_port_y_3;
  wire       [2:0]    m48_mul_port_y_0;
  wire       [2:0]    m48_mul_port_y_1;
  wire       [2:0]    m48_mul_port_y_2;
  wire       [2:0]    m48_mul_port_y_3;
  wire       [2:0]    m49_mul_port_y_0;
  wire       [2:0]    m49_mul_port_y_1;
  wire       [2:0]    m49_mul_port_y_2;
  wire       [2:0]    m49_mul_port_y_3;
  wire       [2:0]    m50_mul_port_y_0;
  wire       [2:0]    m50_mul_port_y_1;
  wire       [2:0]    m50_mul_port_y_2;
  wire       [2:0]    m50_mul_port_y_3;
  wire       [2:0]    m51_mul_port_y_0;
  wire       [2:0]    m51_mul_port_y_1;
  wire       [2:0]    m51_mul_port_y_2;
  wire       [2:0]    m51_mul_port_y_3;
  wire       [2:0]    m52_mul_port_y_0;
  wire       [2:0]    m52_mul_port_y_1;
  wire       [2:0]    m52_mul_port_y_2;
  wire       [2:0]    m52_mul_port_y_3;
  wire       [2:0]    m53_mul_port_y_0;
  wire       [2:0]    m53_mul_port_y_1;
  wire       [2:0]    m53_mul_port_y_2;
  wire       [2:0]    m53_mul_port_y_3;
  wire       [2:0]    m54_mul_port_y_0;
  wire       [2:0]    m54_mul_port_y_1;
  wire       [2:0]    m54_mul_port_y_2;
  wire       [2:0]    m54_mul_port_y_3;
  wire       [2:0]    m55_mul_port_y_0;
  wire       [2:0]    m55_mul_port_y_1;
  wire       [2:0]    m55_mul_port_y_2;
  wire       [2:0]    m55_mul_port_y_3;
  wire       [2:0]    m56_mul_port_y_0;
  wire       [2:0]    m56_mul_port_y_1;
  wire       [2:0]    m56_mul_port_y_2;
  wire       [2:0]    m56_mul_port_y_3;
  wire       [2:0]    m57_mul_port_y_0;
  wire       [2:0]    m57_mul_port_y_1;
  wire       [2:0]    m57_mul_port_y_2;
  wire       [2:0]    m57_mul_port_y_3;
  wire       [2:0]    m58_mul_port_y_0;
  wire       [2:0]    m58_mul_port_y_1;
  wire       [2:0]    m58_mul_port_y_2;
  wire       [2:0]    m58_mul_port_y_3;
  wire       [2:0]    m59_mul_port_y_0;
  wire       [2:0]    m59_mul_port_y_1;
  wire       [2:0]    m59_mul_port_y_2;
  wire       [2:0]    m59_mul_port_y_3;
  wire       [2:0]    m60_mul_port_y_0;
  wire       [2:0]    m60_mul_port_y_1;
  wire       [2:0]    m60_mul_port_y_2;
  wire       [2:0]    m60_mul_port_y_3;
  wire       [2:0]    m61_mul_port_y_0;
  wire       [2:0]    m61_mul_port_y_1;
  wire       [2:0]    m61_mul_port_y_2;
  wire       [2:0]    m61_mul_port_y_3;
  wire       [2:0]    m62_mul_port_y_0;
  wire       [2:0]    m62_mul_port_y_1;
  wire       [2:0]    m62_mul_port_y_2;
  wire       [2:0]    m62_mul_port_y_3;
  wire       [2:0]    m63_mul_port_y_0;
  wire       [2:0]    m63_mul_port_y_1;
  wire       [2:0]    m63_mul_port_y_2;
  wire       [2:0]    m63_mul_port_y_3;
  wire       [2:0]    l0_xor_port_y_0;
  wire       [2:0]    l0_xor_port_y_1;
  wire       [2:0]    l0_xor_port_y_2;
  wire       [2:0]    l0_xor_port_y_3;
  wire       [2:0]    l1_xor_port_y_0;
  wire       [2:0]    l1_xor_port_y_1;
  wire       [2:0]    l1_xor_port_y_2;
  wire       [2:0]    l1_xor_port_y_3;
  wire       [2:0]    l2_xor_port_y_0;
  wire       [2:0]    l2_xor_port_y_1;
  wire       [2:0]    l2_xor_port_y_2;
  wire       [2:0]    l2_xor_port_y_3;
  wire       [2:0]    l3_xor_port_y_0;
  wire       [2:0]    l3_xor_port_y_1;
  wire       [2:0]    l3_xor_port_y_2;
  wire       [2:0]    l3_xor_port_y_3;
  wire       [2:0]    l4_xor_port_y_0;
  wire       [2:0]    l4_xor_port_y_1;
  wire       [2:0]    l4_xor_port_y_2;
  wire       [2:0]    l4_xor_port_y_3;
  wire       [2:0]    l5_xor_port_y_0;
  wire       [2:0]    l5_xor_port_y_1;
  wire       [2:0]    l5_xor_port_y_2;
  wire       [2:0]    l5_xor_port_y_3;
  wire       [2:0]    l6_xor_port_y_0;
  wire       [2:0]    l6_xor_port_y_1;
  wire       [2:0]    l6_xor_port_y_2;
  wire       [2:0]    l6_xor_port_y_3;
  wire       [2:0]    l7_xor_port_y_0;
  wire       [2:0]    l7_xor_port_y_1;
  wire       [2:0]    l7_xor_port_y_2;
  wire       [2:0]    l7_xor_port_y_3;
  wire       [2:0]    l8_xor_port_y_0;
  wire       [2:0]    l8_xor_port_y_1;
  wire       [2:0]    l8_xor_port_y_2;
  wire       [2:0]    l8_xor_port_y_3;
  wire       [2:0]    l9_xor_port_y_0;
  wire       [2:0]    l9_xor_port_y_1;
  wire       [2:0]    l9_xor_port_y_2;
  wire       [2:0]    l9_xor_port_y_3;
  wire       [2:0]    l10_xor_port_y_0;
  wire       [2:0]    l10_xor_port_y_1;
  wire       [2:0]    l10_xor_port_y_2;
  wire       [2:0]    l10_xor_port_y_3;
  wire       [2:0]    l11_xor_port_y_0;
  wire       [2:0]    l11_xor_port_y_1;
  wire       [2:0]    l11_xor_port_y_2;
  wire       [2:0]    l11_xor_port_y_3;
  wire       [2:0]    l12_xor_port_y_0;
  wire       [2:0]    l12_xor_port_y_1;
  wire       [2:0]    l12_xor_port_y_2;
  wire       [2:0]    l12_xor_port_y_3;
  wire       [2:0]    l13_xor_port_y_0;
  wire       [2:0]    l13_xor_port_y_1;
  wire       [2:0]    l13_xor_port_y_2;
  wire       [2:0]    l13_xor_port_y_3;
  wire       [2:0]    l14_xor_port_y_0;
  wire       [2:0]    l14_xor_port_y_1;
  wire       [2:0]    l14_xor_port_y_2;
  wire       [2:0]    l14_xor_port_y_3;
  wire       [2:0]    l15_xor_port_y_0;
  wire       [2:0]    l15_xor_port_y_1;
  wire       [2:0]    l15_xor_port_y_2;
  wire       [2:0]    l15_xor_port_y_3;
  wire       [2:0]    l16_xor_port_y_0;
  wire       [2:0]    l16_xor_port_y_1;
  wire       [2:0]    l16_xor_port_y_2;
  wire       [2:0]    l16_xor_port_y_3;
  wire       [2:0]    l17_xor_port_y_0;
  wire       [2:0]    l17_xor_port_y_1;
  wire       [2:0]    l17_xor_port_y_2;
  wire       [2:0]    l17_xor_port_y_3;
  wire       [2:0]    l18_xor_port_y_0;
  wire       [2:0]    l18_xor_port_y_1;
  wire       [2:0]    l18_xor_port_y_2;
  wire       [2:0]    l18_xor_port_y_3;
  wire       [2:0]    l19_xor_port_y_0;
  wire       [2:0]    l19_xor_port_y_1;
  wire       [2:0]    l19_xor_port_y_2;
  wire       [2:0]    l19_xor_port_y_3;
  wire       [2:0]    l20_xor_port_y_0;
  wire       [2:0]    l20_xor_port_y_1;
  wire       [2:0]    l20_xor_port_y_2;
  wire       [2:0]    l20_xor_port_y_3;
  wire       [2:0]    l21_xor_port_y_0;
  wire       [2:0]    l21_xor_port_y_1;
  wire       [2:0]    l21_xor_port_y_2;
  wire       [2:0]    l21_xor_port_y_3;
  wire       [2:0]    l22_xor_port_y_0;
  wire       [2:0]    l22_xor_port_y_1;
  wire       [2:0]    l22_xor_port_y_2;
  wire       [2:0]    l22_xor_port_y_3;
  wire       [2:0]    l23_xor_port_y_0;
  wire       [2:0]    l23_xor_port_y_1;
  wire       [2:0]    l23_xor_port_y_2;
  wire       [2:0]    l23_xor_port_y_3;
  wire       [2:0]    l24_xor_port_y_0;
  wire       [2:0]    l24_xor_port_y_1;
  wire       [2:0]    l24_xor_port_y_2;
  wire       [2:0]    l24_xor_port_y_3;
  wire       [2:0]    l25_xor_port_y_0;
  wire       [2:0]    l25_xor_port_y_1;
  wire       [2:0]    l25_xor_port_y_2;
  wire       [2:0]    l25_xor_port_y_3;
  wire       [2:0]    l26_xor_port_y_0;
  wire       [2:0]    l26_xor_port_y_1;
  wire       [2:0]    l26_xor_port_y_2;
  wire       [2:0]    l26_xor_port_y_3;
  wire       [2:0]    l27_xor_port_y_0;
  wire       [2:0]    l27_xor_port_y_1;
  wire       [2:0]    l27_xor_port_y_2;
  wire       [2:0]    l27_xor_port_y_3;
  wire       [2:0]    l28_xor_port_y_0;
  wire       [2:0]    l28_xor_port_y_1;
  wire       [2:0]    l28_xor_port_y_2;
  wire       [2:0]    l28_xor_port_y_3;
  wire       [2:0]    l29_xor_port_y_0;
  wire       [2:0]    l29_xor_port_y_1;
  wire       [2:0]    l29_xor_port_y_2;
  wire       [2:0]    l29_xor_port_y_3;
  wire       [2:0]    s0_port_y_0;
  wire       [2:0]    s0_port_y_1;
  wire       [2:0]    s0_port_y_2;
  wire       [2:0]    s0_port_y_3;
  wire       [2:0]    s1_port_y_0;
  wire       [2:0]    s1_port_y_1;
  wire       [2:0]    s1_port_y_2;
  wire       [2:0]    s1_port_y_3;
  wire       [2:0]    s2_port_y_0;
  wire       [2:0]    s2_port_y_1;
  wire       [2:0]    s2_port_y_2;
  wire       [2:0]    s2_port_y_3;
  wire       [2:0]    s3_port_y_0;
  wire       [2:0]    s3_port_y_1;
  wire       [2:0]    s3_port_y_2;
  wire       [2:0]    s3_port_y_3;
  wire       [2:0]    s4_port_y_0;
  wire       [2:0]    s4_port_y_1;
  wire       [2:0]    s4_port_y_2;
  wire       [2:0]    s4_port_y_3;
  wire       [2:0]    s5_port_y_0;
  wire       [2:0]    s5_port_y_1;
  wire       [2:0]    s5_port_y_2;
  wire       [2:0]    s5_port_y_3;
  wire       [2:0]    s6_port_y_0;
  wire       [2:0]    s6_port_y_1;
  wire       [2:0]    s6_port_y_2;
  wire       [2:0]    s6_port_y_3;
  wire       [2:0]    s7_port_y_0;
  wire       [2:0]    s7_port_y_1;
  wire       [2:0]    s7_port_y_2;
  wire       [2:0]    s7_port_y_3;
  wire       [2:0]    in_x0_0;
  wire       [2:0]    in_x0_1;
  wire       [2:0]    in_x0_2;
  wire       [2:0]    in_x0_3;
  wire       [2:0]    in_x1_0;
  wire       [2:0]    in_x1_1;
  wire       [2:0]    in_x1_2;
  wire       [2:0]    in_x1_3;
  wire       [2:0]    in_x2_0;
  wire       [2:0]    in_x2_1;
  wire       [2:0]    in_x2_2;
  wire       [2:0]    in_x2_3;
  wire       [2:0]    in_x3_0;
  wire       [2:0]    in_x3_1;
  wire       [2:0]    in_x3_2;
  wire       [2:0]    in_x3_3;
  wire       [2:0]    in_x4_0;
  wire       [2:0]    in_x4_1;
  wire       [2:0]    in_x4_2;
  wire       [2:0]    in_x4_3;
  wire       [2:0]    in_x5_0;
  wire       [2:0]    in_x5_1;
  wire       [2:0]    in_x5_2;
  wire       [2:0]    in_x5_3;
  wire       [2:0]    in_x6_0;
  wire       [2:0]    in_x6_1;
  wire       [2:0]    in_x6_2;
  wire       [2:0]    in_x6_3;
  wire       [2:0]    in_x7_0;
  wire       [2:0]    in_x7_1;
  wire       [2:0]    in_x7_2;
  wire       [2:0]    in_x7_3;
  wire       [2:0]    out_y0_0;
  wire       [2:0]    out_y0_1;
  wire       [2:0]    out_y0_2;
  wire       [2:0]    out_y0_3;
  wire       [2:0]    out_y1_0;
  wire       [2:0]    out_y1_1;
  wire       [2:0]    out_y1_2;
  wire       [2:0]    out_y1_3;
  wire       [2:0]    out_y2_0;
  wire       [2:0]    out_y2_1;
  wire       [2:0]    out_y2_2;
  wire       [2:0]    out_y2_3;
  wire       [2:0]    out_y3_0;
  wire       [2:0]    out_y3_1;
  wire       [2:0]    out_y3_2;
  wire       [2:0]    out_y3_3;
  wire       [2:0]    out_y4_0;
  wire       [2:0]    out_y4_1;
  wire       [2:0]    out_y4_2;
  wire       [2:0]    out_y4_3;
  wire       [2:0]    out_y5_0;
  wire       [2:0]    out_y5_1;
  wire       [2:0]    out_y5_2;
  wire       [2:0]    out_y5_3;
  wire       [2:0]    out_y6_0;
  wire       [2:0]    out_y6_1;
  wire       [2:0]    out_y6_2;
  wire       [2:0]    out_y6_3;
  wire       [2:0]    out_y7_0;
  wire       [2:0]    out_y7_1;
  wire       [2:0]    out_y7_2;
  wire       [2:0]    out_y7_3;
  reg        [2:0]    x7_0;
  reg        [2:0]    x7_1;
  reg        [2:0]    x7_2;
  reg        [2:0]    x7_3;
  reg        [2:0]    t1_0;
  reg        [2:0]    t1_1;
  reg        [2:0]    t1_2;
  reg        [2:0]    t1_3;
  reg        [2:0]    t2_0;
  reg        [2:0]    t2_1;
  reg        [2:0]    t2_2;
  reg        [2:0]    t2_3;
  reg        [2:0]    t3_0;
  reg        [2:0]    t3_1;
  reg        [2:0]    t3_2;
  reg        [2:0]    t3_3;
  reg        [2:0]    t4_0;
  reg        [2:0]    t4_1;
  reg        [2:0]    t4_2;
  reg        [2:0]    t4_3;
  reg        [2:0]    t6_0;
  reg        [2:0]    t6_1;
  reg        [2:0]    t6_2;
  reg        [2:0]    t6_3;
  reg        [2:0]    t7_0;
  reg        [2:0]    t7_1;
  reg        [2:0]    t7_2;
  reg        [2:0]    t7_3;
  reg        [2:0]    t8_0;
  reg        [2:0]    t8_1;
  reg        [2:0]    t8_2;
  reg        [2:0]    t8_3;
  reg        [2:0]    t9_0;
  reg        [2:0]    t9_1;
  reg        [2:0]    t9_2;
  reg        [2:0]    t9_3;
  reg        [2:0]    t10_0;
  reg        [2:0]    t10_1;
  reg        [2:0]    t10_2;
  reg        [2:0]    t10_3;
  reg        [2:0]    t13_0;
  reg        [2:0]    t13_1;
  reg        [2:0]    t13_2;
  reg        [2:0]    t13_3;
  reg        [2:0]    t14_0;
  reg        [2:0]    t14_1;
  reg        [2:0]    t14_2;
  reg        [2:0]    t14_3;
  reg        [2:0]    t15_0;
  reg        [2:0]    t15_1;
  reg        [2:0]    t15_2;
  reg        [2:0]    t15_3;
  reg        [2:0]    t16_0;
  reg        [2:0]    t16_1;
  reg        [2:0]    t16_2;
  reg        [2:0]    t16_3;
  reg        [2:0]    t17_0;
  reg        [2:0]    t17_1;
  reg        [2:0]    t17_2;
  reg        [2:0]    t17_3;
  reg        [2:0]    t19_0;
  reg        [2:0]    t19_1;
  reg        [2:0]    t19_2;
  reg        [2:0]    t19_3;
  reg        [2:0]    t20_0;
  reg        [2:0]    t20_1;
  reg        [2:0]    t20_2;
  reg        [2:0]    t20_3;
  reg        [2:0]    t22_0;
  reg        [2:0]    t22_1;
  reg        [2:0]    t22_2;
  reg        [2:0]    t22_3;
  reg        [2:0]    t23_0;
  reg        [2:0]    t23_1;
  reg        [2:0]    t23_2;
  reg        [2:0]    t23_3;
  reg        [2:0]    t24_0;
  reg        [2:0]    t24_1;
  reg        [2:0]    t24_2;
  reg        [2:0]    t24_3;
  reg        [2:0]    t25_0;
  reg        [2:0]    t25_1;
  reg        [2:0]    t25_2;
  reg        [2:0]    t25_3;
  reg        [2:0]    t26_0;
  reg        [2:0]    t26_1;
  reg        [2:0]    t26_2;
  reg        [2:0]    t26_3;
  reg        [2:0]    t27_0;
  reg        [2:0]    t27_1;
  reg        [2:0]    t27_2;
  reg        [2:0]    t27_3;
  reg        [2:0]    x7_1_0;
  reg        [2:0]    x7_1_1;
  reg        [2:0]    x7_1_2;
  reg        [2:0]    x7_1_3;
  reg        [2:0]    t1_1_0;
  reg        [2:0]    t1_1_1;
  reg        [2:0]    t1_1_2;
  reg        [2:0]    t1_1_3;
  reg        [2:0]    t2_1_0;
  reg        [2:0]    t2_1_1;
  reg        [2:0]    t2_1_2;
  reg        [2:0]    t2_1_3;
  reg        [2:0]    t3_1_0;
  reg        [2:0]    t3_1_1;
  reg        [2:0]    t3_1_2;
  reg        [2:0]    t3_1_3;
  reg        [2:0]    t4_1_0;
  reg        [2:0]    t4_1_1;
  reg        [2:0]    t4_1_2;
  reg        [2:0]    t4_1_3;
  reg        [2:0]    t6_1_0;
  reg        [2:0]    t6_1_1;
  reg        [2:0]    t6_1_2;
  reg        [2:0]    t6_1_3;
  reg        [2:0]    t8_1_0;
  reg        [2:0]    t8_1_1;
  reg        [2:0]    t8_1_2;
  reg        [2:0]    t8_1_3;
  reg        [2:0]    t9_1_0;
  reg        [2:0]    t9_1_1;
  reg        [2:0]    t9_1_2;
  reg        [2:0]    t9_1_3;
  reg        [2:0]    t10_1_0;
  reg        [2:0]    t10_1_1;
  reg        [2:0]    t10_1_2;
  reg        [2:0]    t10_1_3;
  reg        [2:0]    t13_1_0;
  reg        [2:0]    t13_1_1;
  reg        [2:0]    t13_1_2;
  reg        [2:0]    t13_1_3;
  reg        [2:0]    t15_1_0;
  reg        [2:0]    t15_1_1;
  reg        [2:0]    t15_1_2;
  reg        [2:0]    t15_1_3;
  reg        [2:0]    t16_1_0;
  reg        [2:0]    t16_1_1;
  reg        [2:0]    t16_1_2;
  reg        [2:0]    t16_1_3;
  reg        [2:0]    t17_1_0;
  reg        [2:0]    t17_1_1;
  reg        [2:0]    t17_1_2;
  reg        [2:0]    t17_1_3;
  reg        [2:0]    t19_1_0;
  reg        [2:0]    t19_1_1;
  reg        [2:0]    t19_1_2;
  reg        [2:0]    t19_1_3;
  reg        [2:0]    t20_1_0;
  reg        [2:0]    t20_1_1;
  reg        [2:0]    t20_1_2;
  reg        [2:0]    t20_1_3;
  reg        [2:0]    t22_1_0;
  reg        [2:0]    t22_1_1;
  reg        [2:0]    t22_1_2;
  reg        [2:0]    t22_1_3;
  reg        [2:0]    t23_1_0;
  reg        [2:0]    t23_1_1;
  reg        [2:0]    t23_1_2;
  reg        [2:0]    t23_1_3;
  reg        [2:0]    t27_1_0;
  reg        [2:0]    t27_1_1;
  reg        [2:0]    t27_1_2;
  reg        [2:0]    t27_1_3;
  reg        [2:0]    m21_0;
  reg        [2:0]    m21_1;
  reg        [2:0]    m21_2;
  reg        [2:0]    m21_3;
  reg        [2:0]    m23_0;
  reg        [2:0]    m23_1;
  reg        [2:0]    m23_2;
  reg        [2:0]    m23_3;
  reg        [2:0]    m24_0;
  reg        [2:0]    m24_1;
  reg        [2:0]    m24_2;
  reg        [2:0]    m24_3;
  reg        [2:0]    m27_0;
  reg        [2:0]    m27_1;
  reg        [2:0]    m27_2;
  reg        [2:0]    m27_3;
  reg        [2:0]    x7_2_0;
  reg        [2:0]    x7_2_1;
  reg        [2:0]    x7_2_2;
  reg        [2:0]    x7_2_3;
  reg        [2:0]    t1_2_0;
  reg        [2:0]    t1_2_1;
  reg        [2:0]    t1_2_2;
  reg        [2:0]    t1_2_3;
  reg        [2:0]    t2_2_0;
  reg        [2:0]    t2_2_1;
  reg        [2:0]    t2_2_2;
  reg        [2:0]    t2_2_3;
  reg        [2:0]    t3_2_0;
  reg        [2:0]    t3_2_1;
  reg        [2:0]    t3_2_2;
  reg        [2:0]    t3_2_3;
  reg        [2:0]    t4_2_0;
  reg        [2:0]    t4_2_1;
  reg        [2:0]    t4_2_2;
  reg        [2:0]    t4_2_3;
  reg        [2:0]    t6_2_0;
  reg        [2:0]    t6_2_1;
  reg        [2:0]    t6_2_2;
  reg        [2:0]    t6_2_3;
  reg        [2:0]    t8_2_0;
  reg        [2:0]    t8_2_1;
  reg        [2:0]    t8_2_2;
  reg        [2:0]    t8_2_3;
  reg        [2:0]    t9_2_0;
  reg        [2:0]    t9_2_1;
  reg        [2:0]    t9_2_2;
  reg        [2:0]    t9_2_3;
  reg        [2:0]    t10_2_0;
  reg        [2:0]    t10_2_1;
  reg        [2:0]    t10_2_2;
  reg        [2:0]    t10_2_3;
  reg        [2:0]    t13_2_0;
  reg        [2:0]    t13_2_1;
  reg        [2:0]    t13_2_2;
  reg        [2:0]    t13_2_3;
  reg        [2:0]    t15_2_0;
  reg        [2:0]    t15_2_1;
  reg        [2:0]    t15_2_2;
  reg        [2:0]    t15_2_3;
  reg        [2:0]    t16_2_0;
  reg        [2:0]    t16_2_1;
  reg        [2:0]    t16_2_2;
  reg        [2:0]    t16_2_3;
  reg        [2:0]    t17_2_0;
  reg        [2:0]    t17_2_1;
  reg        [2:0]    t17_2_2;
  reg        [2:0]    t17_2_3;
  reg        [2:0]    t19_2_0;
  reg        [2:0]    t19_2_1;
  reg        [2:0]    t19_2_2;
  reg        [2:0]    t19_2_3;
  reg        [2:0]    t20_2_0;
  reg        [2:0]    t20_2_1;
  reg        [2:0]    t20_2_2;
  reg        [2:0]    t20_2_3;
  reg        [2:0]    t22_2_0;
  reg        [2:0]    t22_2_1;
  reg        [2:0]    t22_2_2;
  reg        [2:0]    t22_2_3;
  reg        [2:0]    t23_2_0;
  reg        [2:0]    t23_2_1;
  reg        [2:0]    t23_2_2;
  reg        [2:0]    t23_2_3;
  reg        [2:0]    t27_2_0;
  reg        [2:0]    t27_2_1;
  reg        [2:0]    t27_2_2;
  reg        [2:0]    t27_2_3;
  reg        [2:0]    m21_1_0;
  reg        [2:0]    m21_1_1;
  reg        [2:0]    m21_1_2;
  reg        [2:0]    m21_1_3;
  reg        [2:0]    m23_1_0;
  reg        [2:0]    m23_1_1;
  reg        [2:0]    m23_1_2;
  reg        [2:0]    m23_1_3;
  reg        [2:0]    m33_0;
  reg        [2:0]    m33_1;
  reg        [2:0]    m33_2;
  reg        [2:0]    m33_3;
  reg        [2:0]    m36_0;
  reg        [2:0]    m36_1;
  reg        [2:0]    m36_2;
  reg        [2:0]    m36_3;

  Addition_TI t1_xor (
    .port_x0_0 (in_x0_0[2:0]        ), //i
    .port_x0_1 (in_x0_1[2:0]        ), //i
    .port_x0_2 (in_x0_2[2:0]        ), //i
    .port_x0_3 (in_x0_3[2:0]        ), //i
    .port_x1_0 (in_x3_0[2:0]        ), //i
    .port_x1_1 (in_x3_1[2:0]        ), //i
    .port_x1_2 (in_x3_2[2:0]        ), //i
    .port_x1_3 (in_x3_3[2:0]        ), //i
    .port_y_0  (t1_xor_port_y_0[2:0]), //o
    .port_y_1  (t1_xor_port_y_1[2:0]), //o
    .port_y_2  (t1_xor_port_y_2[2:0]), //o
    .port_y_3  (t1_xor_port_y_3[2:0])  //o
  );
  Addition_TI t2_xor (
    .port_x0_0 (in_x0_0[2:0]        ), //i
    .port_x0_1 (in_x0_1[2:0]        ), //i
    .port_x0_2 (in_x0_2[2:0]        ), //i
    .port_x0_3 (in_x0_3[2:0]        ), //i
    .port_x1_0 (in_x5_0[2:0]        ), //i
    .port_x1_1 (in_x5_1[2:0]        ), //i
    .port_x1_2 (in_x5_2[2:0]        ), //i
    .port_x1_3 (in_x5_3[2:0]        ), //i
    .port_y_0  (t2_xor_port_y_0[2:0]), //o
    .port_y_1  (t2_xor_port_y_1[2:0]), //o
    .port_y_2  (t2_xor_port_y_2[2:0]), //o
    .port_y_3  (t2_xor_port_y_3[2:0])  //o
  );
  Addition_TI t3_xor (
    .port_x0_0 (in_x0_0[2:0]        ), //i
    .port_x0_1 (in_x0_1[2:0]        ), //i
    .port_x0_2 (in_x0_2[2:0]        ), //i
    .port_x0_3 (in_x0_3[2:0]        ), //i
    .port_x1_0 (in_x6_0[2:0]        ), //i
    .port_x1_1 (in_x6_1[2:0]        ), //i
    .port_x1_2 (in_x6_2[2:0]        ), //i
    .port_x1_3 (in_x6_3[2:0]        ), //i
    .port_y_0  (t3_xor_port_y_0[2:0]), //o
    .port_y_1  (t3_xor_port_y_1[2:0]), //o
    .port_y_2  (t3_xor_port_y_2[2:0]), //o
    .port_y_3  (t3_xor_port_y_3[2:0])  //o
  );
  Addition_TI t4_xor (
    .port_x0_0 (in_x3_0[2:0]        ), //i
    .port_x0_1 (in_x3_1[2:0]        ), //i
    .port_x0_2 (in_x3_2[2:0]        ), //i
    .port_x0_3 (in_x3_3[2:0]        ), //i
    .port_x1_0 (in_x5_0[2:0]        ), //i
    .port_x1_1 (in_x5_1[2:0]        ), //i
    .port_x1_2 (in_x5_2[2:0]        ), //i
    .port_x1_3 (in_x5_3[2:0]        ), //i
    .port_y_0  (t4_xor_port_y_0[2:0]), //o
    .port_y_1  (t4_xor_port_y_1[2:0]), //o
    .port_y_2  (t4_xor_port_y_2[2:0]), //o
    .port_y_3  (t4_xor_port_y_3[2:0])  //o
  );
  Addition_TI t5_xor (
    .port_x0_0 (in_x4_0[2:0]        ), //i
    .port_x0_1 (in_x4_1[2:0]        ), //i
    .port_x0_2 (in_x4_2[2:0]        ), //i
    .port_x0_3 (in_x4_3[2:0]        ), //i
    .port_x1_0 (in_x6_0[2:0]        ), //i
    .port_x1_1 (in_x6_1[2:0]        ), //i
    .port_x1_2 (in_x6_2[2:0]        ), //i
    .port_x1_3 (in_x6_3[2:0]        ), //i
    .port_y_0  (t5_xor_port_y_0[2:0]), //o
    .port_y_1  (t5_xor_port_y_1[2:0]), //o
    .port_y_2  (t5_xor_port_y_2[2:0]), //o
    .port_y_3  (t5_xor_port_y_3[2:0])  //o
  );
  Addition_TI t6_xor (
    .port_x0_0 (t1_xor_port_y_0[2:0]), //i
    .port_x0_1 (t1_xor_port_y_1[2:0]), //i
    .port_x0_2 (t1_xor_port_y_2[2:0]), //i
    .port_x0_3 (t1_xor_port_y_3[2:0]), //i
    .port_x1_0 (t5_xor_port_y_0[2:0]), //i
    .port_x1_1 (t5_xor_port_y_1[2:0]), //i
    .port_x1_2 (t5_xor_port_y_2[2:0]), //i
    .port_x1_3 (t5_xor_port_y_3[2:0]), //i
    .port_y_0  (t6_xor_port_y_0[2:0]), //o
    .port_y_1  (t6_xor_port_y_1[2:0]), //o
    .port_y_2  (t6_xor_port_y_2[2:0]), //o
    .port_y_3  (t6_xor_port_y_3[2:0])  //o
  );
  Addition_TI t7_xor (
    .port_x0_0 (in_x1_0[2:0]        ), //i
    .port_x0_1 (in_x1_1[2:0]        ), //i
    .port_x0_2 (in_x1_2[2:0]        ), //i
    .port_x0_3 (in_x1_3[2:0]        ), //i
    .port_x1_0 (in_x2_0[2:0]        ), //i
    .port_x1_1 (in_x2_1[2:0]        ), //i
    .port_x1_2 (in_x2_2[2:0]        ), //i
    .port_x1_3 (in_x2_3[2:0]        ), //i
    .port_y_0  (t7_xor_port_y_0[2:0]), //o
    .port_y_1  (t7_xor_port_y_1[2:0]), //o
    .port_y_2  (t7_xor_port_y_2[2:0]), //o
    .port_y_3  (t7_xor_port_y_3[2:0])  //o
  );
  Addition_TI t8_xor (
    .port_x0_0 (in_x7_0[2:0]        ), //i
    .port_x0_1 (in_x7_1[2:0]        ), //i
    .port_x0_2 (in_x7_2[2:0]        ), //i
    .port_x0_3 (in_x7_3[2:0]        ), //i
    .port_x1_0 (t6_xor_port_y_0[2:0]), //i
    .port_x1_1 (t6_xor_port_y_1[2:0]), //i
    .port_x1_2 (t6_xor_port_y_2[2:0]), //i
    .port_x1_3 (t6_xor_port_y_3[2:0]), //i
    .port_y_0  (t8_xor_port_y_0[2:0]), //o
    .port_y_1  (t8_xor_port_y_1[2:0]), //o
    .port_y_2  (t8_xor_port_y_2[2:0]), //o
    .port_y_3  (t8_xor_port_y_3[2:0])  //o
  );
  Addition_TI t9_xor (
    .port_x0_0 (in_x7_0[2:0]        ), //i
    .port_x0_1 (in_x7_1[2:0]        ), //i
    .port_x0_2 (in_x7_2[2:0]        ), //i
    .port_x0_3 (in_x7_3[2:0]        ), //i
    .port_x1_0 (t7_xor_port_y_0[2:0]), //i
    .port_x1_1 (t7_xor_port_y_1[2:0]), //i
    .port_x1_2 (t7_xor_port_y_2[2:0]), //i
    .port_x1_3 (t7_xor_port_y_3[2:0]), //i
    .port_y_0  (t9_xor_port_y_0[2:0]), //o
    .port_y_1  (t9_xor_port_y_1[2:0]), //o
    .port_y_2  (t9_xor_port_y_2[2:0]), //o
    .port_y_3  (t9_xor_port_y_3[2:0])  //o
  );
  Addition_TI t10_xor (
    .port_x0_0 (t6_xor_port_y_0[2:0] ), //i
    .port_x0_1 (t6_xor_port_y_1[2:0] ), //i
    .port_x0_2 (t6_xor_port_y_2[2:0] ), //i
    .port_x0_3 (t6_xor_port_y_3[2:0] ), //i
    .port_x1_0 (t7_xor_port_y_0[2:0] ), //i
    .port_x1_1 (t7_xor_port_y_1[2:0] ), //i
    .port_x1_2 (t7_xor_port_y_2[2:0] ), //i
    .port_x1_3 (t7_xor_port_y_3[2:0] ), //i
    .port_y_0  (t10_xor_port_y_0[2:0]), //o
    .port_y_1  (t10_xor_port_y_1[2:0]), //o
    .port_y_2  (t10_xor_port_y_2[2:0]), //o
    .port_y_3  (t10_xor_port_y_3[2:0])  //o
  );
  Addition_TI t11_xor (
    .port_x0_0 (in_x1_0[2:0]         ), //i
    .port_x0_1 (in_x1_1[2:0]         ), //i
    .port_x0_2 (in_x1_2[2:0]         ), //i
    .port_x0_3 (in_x1_3[2:0]         ), //i
    .port_x1_0 (in_x5_0[2:0]         ), //i
    .port_x1_1 (in_x5_1[2:0]         ), //i
    .port_x1_2 (in_x5_2[2:0]         ), //i
    .port_x1_3 (in_x5_3[2:0]         ), //i
    .port_y_0  (t11_xor_port_y_0[2:0]), //o
    .port_y_1  (t11_xor_port_y_1[2:0]), //o
    .port_y_2  (t11_xor_port_y_2[2:0]), //o
    .port_y_3  (t11_xor_port_y_3[2:0])  //o
  );
  Addition_TI t12_xor (
    .port_x0_0 (in_x2_0[2:0]         ), //i
    .port_x0_1 (in_x2_1[2:0]         ), //i
    .port_x0_2 (in_x2_2[2:0]         ), //i
    .port_x0_3 (in_x2_3[2:0]         ), //i
    .port_x1_0 (in_x5_0[2:0]         ), //i
    .port_x1_1 (in_x5_1[2:0]         ), //i
    .port_x1_2 (in_x5_2[2:0]         ), //i
    .port_x1_3 (in_x5_3[2:0]         ), //i
    .port_y_0  (t12_xor_port_y_0[2:0]), //o
    .port_y_1  (t12_xor_port_y_1[2:0]), //o
    .port_y_2  (t12_xor_port_y_2[2:0]), //o
    .port_y_3  (t12_xor_port_y_3[2:0])  //o
  );
  Addition_TI t13_xor (
    .port_x0_0 (t3_xor_port_y_0[2:0] ), //i
    .port_x0_1 (t3_xor_port_y_1[2:0] ), //i
    .port_x0_2 (t3_xor_port_y_2[2:0] ), //i
    .port_x0_3 (t3_xor_port_y_3[2:0] ), //i
    .port_x1_0 (t4_xor_port_y_0[2:0] ), //i
    .port_x1_1 (t4_xor_port_y_1[2:0] ), //i
    .port_x1_2 (t4_xor_port_y_2[2:0] ), //i
    .port_x1_3 (t4_xor_port_y_3[2:0] ), //i
    .port_y_0  (t13_xor_port_y_0[2:0]), //o
    .port_y_1  (t13_xor_port_y_1[2:0]), //o
    .port_y_2  (t13_xor_port_y_2[2:0]), //o
    .port_y_3  (t13_xor_port_y_3[2:0])  //o
  );
  Addition_TI t14_xor (
    .port_x0_0 (t6_xor_port_y_0[2:0] ), //i
    .port_x0_1 (t6_xor_port_y_1[2:0] ), //i
    .port_x0_2 (t6_xor_port_y_2[2:0] ), //i
    .port_x0_3 (t6_xor_port_y_3[2:0] ), //i
    .port_x1_0 (t11_xor_port_y_0[2:0]), //i
    .port_x1_1 (t11_xor_port_y_1[2:0]), //i
    .port_x1_2 (t11_xor_port_y_2[2:0]), //i
    .port_x1_3 (t11_xor_port_y_3[2:0]), //i
    .port_y_0  (t14_xor_port_y_0[2:0]), //o
    .port_y_1  (t14_xor_port_y_1[2:0]), //o
    .port_y_2  (t14_xor_port_y_2[2:0]), //o
    .port_y_3  (t14_xor_port_y_3[2:0])  //o
  );
  Addition_TI t15_xor (
    .port_x0_0 (t5_xor_port_y_0[2:0] ), //i
    .port_x0_1 (t5_xor_port_y_1[2:0] ), //i
    .port_x0_2 (t5_xor_port_y_2[2:0] ), //i
    .port_x0_3 (t5_xor_port_y_3[2:0] ), //i
    .port_x1_0 (t11_xor_port_y_0[2:0]), //i
    .port_x1_1 (t11_xor_port_y_1[2:0]), //i
    .port_x1_2 (t11_xor_port_y_2[2:0]), //i
    .port_x1_3 (t11_xor_port_y_3[2:0]), //i
    .port_y_0  (t15_xor_port_y_0[2:0]), //o
    .port_y_1  (t15_xor_port_y_1[2:0]), //o
    .port_y_2  (t15_xor_port_y_2[2:0]), //o
    .port_y_3  (t15_xor_port_y_3[2:0])  //o
  );
  Addition_TI t16_xor (
    .port_x0_0 (t5_xor_port_y_0[2:0] ), //i
    .port_x0_1 (t5_xor_port_y_1[2:0] ), //i
    .port_x0_2 (t5_xor_port_y_2[2:0] ), //i
    .port_x0_3 (t5_xor_port_y_3[2:0] ), //i
    .port_x1_0 (t12_xor_port_y_0[2:0]), //i
    .port_x1_1 (t12_xor_port_y_1[2:0]), //i
    .port_x1_2 (t12_xor_port_y_2[2:0]), //i
    .port_x1_3 (t12_xor_port_y_3[2:0]), //i
    .port_y_0  (t16_xor_port_y_0[2:0]), //o
    .port_y_1  (t16_xor_port_y_1[2:0]), //o
    .port_y_2  (t16_xor_port_y_2[2:0]), //o
    .port_y_3  (t16_xor_port_y_3[2:0])  //o
  );
  Addition_TI t17_xor (
    .port_x0_0 (t9_xor_port_y_0[2:0] ), //i
    .port_x0_1 (t9_xor_port_y_1[2:0] ), //i
    .port_x0_2 (t9_xor_port_y_2[2:0] ), //i
    .port_x0_3 (t9_xor_port_y_3[2:0] ), //i
    .port_x1_0 (t16_xor_port_y_0[2:0]), //i
    .port_x1_1 (t16_xor_port_y_1[2:0]), //i
    .port_x1_2 (t16_xor_port_y_2[2:0]), //i
    .port_x1_3 (t16_xor_port_y_3[2:0]), //i
    .port_y_0  (t17_xor_port_y_0[2:0]), //o
    .port_y_1  (t17_xor_port_y_1[2:0]), //o
    .port_y_2  (t17_xor_port_y_2[2:0]), //o
    .port_y_3  (t17_xor_port_y_3[2:0])  //o
  );
  Addition_TI t18_xor (
    .port_x0_0 (in_x3_0[2:0]         ), //i
    .port_x0_1 (in_x3_1[2:0]         ), //i
    .port_x0_2 (in_x3_2[2:0]         ), //i
    .port_x0_3 (in_x3_3[2:0]         ), //i
    .port_x1_0 (in_x7_0[2:0]         ), //i
    .port_x1_1 (in_x7_1[2:0]         ), //i
    .port_x1_2 (in_x7_2[2:0]         ), //i
    .port_x1_3 (in_x7_3[2:0]         ), //i
    .port_y_0  (t18_xor_port_y_0[2:0]), //o
    .port_y_1  (t18_xor_port_y_1[2:0]), //o
    .port_y_2  (t18_xor_port_y_2[2:0]), //o
    .port_y_3  (t18_xor_port_y_3[2:0])  //o
  );
  Addition_TI t19_xor (
    .port_x0_0 (t7_xor_port_y_0[2:0] ), //i
    .port_x0_1 (t7_xor_port_y_1[2:0] ), //i
    .port_x0_2 (t7_xor_port_y_2[2:0] ), //i
    .port_x0_3 (t7_xor_port_y_3[2:0] ), //i
    .port_x1_0 (t18_xor_port_y_0[2:0]), //i
    .port_x1_1 (t18_xor_port_y_1[2:0]), //i
    .port_x1_2 (t18_xor_port_y_2[2:0]), //i
    .port_x1_3 (t18_xor_port_y_3[2:0]), //i
    .port_y_0  (t19_xor_port_y_0[2:0]), //o
    .port_y_1  (t19_xor_port_y_1[2:0]), //o
    .port_y_2  (t19_xor_port_y_2[2:0]), //o
    .port_y_3  (t19_xor_port_y_3[2:0])  //o
  );
  Addition_TI t20_xor (
    .port_x0_0 (t1_xor_port_y_0[2:0] ), //i
    .port_x0_1 (t1_xor_port_y_1[2:0] ), //i
    .port_x0_2 (t1_xor_port_y_2[2:0] ), //i
    .port_x0_3 (t1_xor_port_y_3[2:0] ), //i
    .port_x1_0 (t19_xor_port_y_0[2:0]), //i
    .port_x1_1 (t19_xor_port_y_1[2:0]), //i
    .port_x1_2 (t19_xor_port_y_2[2:0]), //i
    .port_x1_3 (t19_xor_port_y_3[2:0]), //i
    .port_y_0  (t20_xor_port_y_0[2:0]), //o
    .port_y_1  (t20_xor_port_y_1[2:0]), //o
    .port_y_2  (t20_xor_port_y_2[2:0]), //o
    .port_y_3  (t20_xor_port_y_3[2:0])  //o
  );
  Addition_TI t21_xor (
    .port_x0_0 (in_x6_0[2:0]         ), //i
    .port_x0_1 (in_x6_1[2:0]         ), //i
    .port_x0_2 (in_x6_2[2:0]         ), //i
    .port_x0_3 (in_x6_3[2:0]         ), //i
    .port_x1_0 (in_x7_0[2:0]         ), //i
    .port_x1_1 (in_x7_1[2:0]         ), //i
    .port_x1_2 (in_x7_2[2:0]         ), //i
    .port_x1_3 (in_x7_3[2:0]         ), //i
    .port_y_0  (t21_xor_port_y_0[2:0]), //o
    .port_y_1  (t21_xor_port_y_1[2:0]), //o
    .port_y_2  (t21_xor_port_y_2[2:0]), //o
    .port_y_3  (t21_xor_port_y_3[2:0])  //o
  );
  Addition_TI t22_xor (
    .port_x0_0 (t7_xor_port_y_0[2:0] ), //i
    .port_x0_1 (t7_xor_port_y_1[2:0] ), //i
    .port_x0_2 (t7_xor_port_y_2[2:0] ), //i
    .port_x0_3 (t7_xor_port_y_3[2:0] ), //i
    .port_x1_0 (t21_xor_port_y_0[2:0]), //i
    .port_x1_1 (t21_xor_port_y_1[2:0]), //i
    .port_x1_2 (t21_xor_port_y_2[2:0]), //i
    .port_x1_3 (t21_xor_port_y_3[2:0]), //i
    .port_y_0  (t22_xor_port_y_0[2:0]), //o
    .port_y_1  (t22_xor_port_y_1[2:0]), //o
    .port_y_2  (t22_xor_port_y_2[2:0]), //o
    .port_y_3  (t22_xor_port_y_3[2:0])  //o
  );
  Addition_TI t23_xor (
    .port_x0_0 (t2_xor_port_y_0[2:0] ), //i
    .port_x0_1 (t2_xor_port_y_1[2:0] ), //i
    .port_x0_2 (t2_xor_port_y_2[2:0] ), //i
    .port_x0_3 (t2_xor_port_y_3[2:0] ), //i
    .port_x1_0 (t22_xor_port_y_0[2:0]), //i
    .port_x1_1 (t22_xor_port_y_1[2:0]), //i
    .port_x1_2 (t22_xor_port_y_2[2:0]), //i
    .port_x1_3 (t22_xor_port_y_3[2:0]), //i
    .port_y_0  (t23_xor_port_y_0[2:0]), //o
    .port_y_1  (t23_xor_port_y_1[2:0]), //o
    .port_y_2  (t23_xor_port_y_2[2:0]), //o
    .port_y_3  (t23_xor_port_y_3[2:0])  //o
  );
  Addition_TI t24_xor (
    .port_x0_0 (t2_xor_port_y_0[2:0] ), //i
    .port_x0_1 (t2_xor_port_y_1[2:0] ), //i
    .port_x0_2 (t2_xor_port_y_2[2:0] ), //i
    .port_x0_3 (t2_xor_port_y_3[2:0] ), //i
    .port_x1_0 (t10_xor_port_y_0[2:0]), //i
    .port_x1_1 (t10_xor_port_y_1[2:0]), //i
    .port_x1_2 (t10_xor_port_y_2[2:0]), //i
    .port_x1_3 (t10_xor_port_y_3[2:0]), //i
    .port_y_0  (t24_xor_port_y_0[2:0]), //o
    .port_y_1  (t24_xor_port_y_1[2:0]), //o
    .port_y_2  (t24_xor_port_y_2[2:0]), //o
    .port_y_3  (t24_xor_port_y_3[2:0])  //o
  );
  Addition_TI t25_xor (
    .port_x0_0 (t20_xor_port_y_0[2:0]), //i
    .port_x0_1 (t20_xor_port_y_1[2:0]), //i
    .port_x0_2 (t20_xor_port_y_2[2:0]), //i
    .port_x0_3 (t20_xor_port_y_3[2:0]), //i
    .port_x1_0 (t17_xor_port_y_0[2:0]), //i
    .port_x1_1 (t17_xor_port_y_1[2:0]), //i
    .port_x1_2 (t17_xor_port_y_2[2:0]), //i
    .port_x1_3 (t17_xor_port_y_3[2:0]), //i
    .port_y_0  (t25_xor_port_y_0[2:0]), //o
    .port_y_1  (t25_xor_port_y_1[2:0]), //o
    .port_y_2  (t25_xor_port_y_2[2:0]), //o
    .port_y_3  (t25_xor_port_y_3[2:0])  //o
  );
  Addition_TI t26_xor (
    .port_x0_0 (t3_xor_port_y_0[2:0] ), //i
    .port_x0_1 (t3_xor_port_y_1[2:0] ), //i
    .port_x0_2 (t3_xor_port_y_2[2:0] ), //i
    .port_x0_3 (t3_xor_port_y_3[2:0] ), //i
    .port_x1_0 (t16_xor_port_y_0[2:0]), //i
    .port_x1_1 (t16_xor_port_y_1[2:0]), //i
    .port_x1_2 (t16_xor_port_y_2[2:0]), //i
    .port_x1_3 (t16_xor_port_y_3[2:0]), //i
    .port_y_0  (t26_xor_port_y_0[2:0]), //o
    .port_y_1  (t26_xor_port_y_1[2:0]), //o
    .port_y_2  (t26_xor_port_y_2[2:0]), //o
    .port_y_3  (t26_xor_port_y_3[2:0])  //o
  );
  Addition_TI t27_xor (
    .port_x0_0 (t1_xor_port_y_0[2:0] ), //i
    .port_x0_1 (t1_xor_port_y_1[2:0] ), //i
    .port_x0_2 (t1_xor_port_y_2[2:0] ), //i
    .port_x0_3 (t1_xor_port_y_3[2:0] ), //i
    .port_x1_0 (t12_xor_port_y_0[2:0]), //i
    .port_x1_1 (t12_xor_port_y_1[2:0]), //i
    .port_x1_2 (t12_xor_port_y_2[2:0]), //i
    .port_x1_3 (t12_xor_port_y_3[2:0]), //i
    .port_y_0  (t27_xor_port_y_0[2:0]), //o
    .port_y_1  (t27_xor_port_y_1[2:0]), //o
    .port_y_2  (t27_xor_port_y_2[2:0]), //o
    .port_y_3  (t27_xor_port_y_3[2:0])  //o
  );
  Multiplication_TI m1 (
    .port_x0_0 (t13_xor_port_y_0[2:0]), //i
    .port_x0_1 (t13_xor_port_y_1[2:0]), //i
    .port_x0_2 (t13_xor_port_y_2[2:0]), //i
    .port_x0_3 (t13_xor_port_y_3[2:0]), //i
    .port_x1_0 (t6_xor_port_y_0[2:0] ), //i
    .port_x1_1 (t6_xor_port_y_1[2:0] ), //i
    .port_x1_2 (t6_xor_port_y_2[2:0] ), //i
    .port_x1_3 (t6_xor_port_y_3[2:0] ), //i
    .port_y_0  (m1_port_y_0[2:0]     ), //o
    .port_y_1  (m1_port_y_1[2:0]     ), //o
    .port_y_2  (m1_port_y_2[2:0]     ), //o
    .port_y_3  (m1_port_y_3[2:0]     ), //o
    .clk       (clk                  ), //i
    .reset     (reset                )  //i
  );
  Multiplication_TI m2 (
    .port_x0_0 (t23_xor_port_y_0[2:0]), //i
    .port_x0_1 (t23_xor_port_y_1[2:0]), //i
    .port_x0_2 (t23_xor_port_y_2[2:0]), //i
    .port_x0_3 (t23_xor_port_y_3[2:0]), //i
    .port_x1_0 (t8_xor_port_y_0[2:0] ), //i
    .port_x1_1 (t8_xor_port_y_1[2:0] ), //i
    .port_x1_2 (t8_xor_port_y_2[2:0] ), //i
    .port_x1_3 (t8_xor_port_y_3[2:0] ), //i
    .port_y_0  (m2_port_y_0[2:0]     ), //o
    .port_y_1  (m2_port_y_1[2:0]     ), //o
    .port_y_2  (m2_port_y_2[2:0]     ), //o
    .port_y_3  (m2_port_y_3[2:0]     ), //o
    .clk       (clk                  ), //i
    .reset     (reset                )  //i
  );
  Multiplication_TI m4 (
    .port_x0_0 (t19_xor_port_y_0[2:0]), //i
    .port_x0_1 (t19_xor_port_y_1[2:0]), //i
    .port_x0_2 (t19_xor_port_y_2[2:0]), //i
    .port_x0_3 (t19_xor_port_y_3[2:0]), //i
    .port_x1_0 (in_x7_0[2:0]         ), //i
    .port_x1_1 (in_x7_1[2:0]         ), //i
    .port_x1_2 (in_x7_2[2:0]         ), //i
    .port_x1_3 (in_x7_3[2:0]         ), //i
    .port_y_0  (m4_port_y_0[2:0]     ), //o
    .port_y_1  (m4_port_y_1[2:0]     ), //o
    .port_y_2  (m4_port_y_2[2:0]     ), //o
    .port_y_3  (m4_port_y_3[2:0]     ), //o
    .clk       (clk                  ), //i
    .reset     (reset                )  //i
  );
  Multiplication_TI m6 (
    .port_x0_0 (t3_xor_port_y_0[2:0] ), //i
    .port_x0_1 (t3_xor_port_y_1[2:0] ), //i
    .port_x0_2 (t3_xor_port_y_2[2:0] ), //i
    .port_x0_3 (t3_xor_port_y_3[2:0] ), //i
    .port_x1_0 (t16_xor_port_y_0[2:0]), //i
    .port_x1_1 (t16_xor_port_y_1[2:0]), //i
    .port_x1_2 (t16_xor_port_y_2[2:0]), //i
    .port_x1_3 (t16_xor_port_y_3[2:0]), //i
    .port_y_0  (m6_port_y_0[2:0]     ), //o
    .port_y_1  (m6_port_y_1[2:0]     ), //o
    .port_y_2  (m6_port_y_2[2:0]     ), //o
    .port_y_3  (m6_port_y_3[2:0]     ), //o
    .clk       (clk                  ), //i
    .reset     (reset                )  //i
  );
  Multiplication_TI m7 (
    .port_x0_0 (t22_xor_port_y_0[2:0]), //i
    .port_x0_1 (t22_xor_port_y_1[2:0]), //i
    .port_x0_2 (t22_xor_port_y_2[2:0]), //i
    .port_x0_3 (t22_xor_port_y_3[2:0]), //i
    .port_x1_0 (t9_xor_port_y_0[2:0] ), //i
    .port_x1_1 (t9_xor_port_y_1[2:0] ), //i
    .port_x1_2 (t9_xor_port_y_2[2:0] ), //i
    .port_x1_3 (t9_xor_port_y_3[2:0] ), //i
    .port_y_0  (m7_port_y_0[2:0]     ), //o
    .port_y_1  (m7_port_y_1[2:0]     ), //o
    .port_y_2  (m7_port_y_2[2:0]     ), //o
    .port_y_3  (m7_port_y_3[2:0]     ), //o
    .clk       (clk                  ), //i
    .reset     (reset                )  //i
  );
  Multiplication_TI m9 (
    .port_x0_0 (t20_xor_port_y_0[2:0]), //i
    .port_x0_1 (t20_xor_port_y_1[2:0]), //i
    .port_x0_2 (t20_xor_port_y_2[2:0]), //i
    .port_x0_3 (t20_xor_port_y_3[2:0]), //i
    .port_x1_0 (t17_xor_port_y_0[2:0]), //i
    .port_x1_1 (t17_xor_port_y_1[2:0]), //i
    .port_x1_2 (t17_xor_port_y_2[2:0]), //i
    .port_x1_3 (t17_xor_port_y_3[2:0]), //i
    .port_y_0  (m9_port_y_0[2:0]     ), //o
    .port_y_1  (m9_port_y_1[2:0]     ), //o
    .port_y_2  (m9_port_y_2[2:0]     ), //o
    .port_y_3  (m9_port_y_3[2:0]     ), //o
    .clk       (clk                  ), //i
    .reset     (reset                )  //i
  );
  Multiplication_TI m11 (
    .port_x0_0 (t1_xor_port_y_0[2:0] ), //i
    .port_x0_1 (t1_xor_port_y_1[2:0] ), //i
    .port_x0_2 (t1_xor_port_y_2[2:0] ), //i
    .port_x0_3 (t1_xor_port_y_3[2:0] ), //i
    .port_x1_0 (t15_xor_port_y_0[2:0]), //i
    .port_x1_1 (t15_xor_port_y_1[2:0]), //i
    .port_x1_2 (t15_xor_port_y_2[2:0]), //i
    .port_x1_3 (t15_xor_port_y_3[2:0]), //i
    .port_y_0  (m11_port_y_0[2:0]    ), //o
    .port_y_1  (m11_port_y_1[2:0]    ), //o
    .port_y_2  (m11_port_y_2[2:0]    ), //o
    .port_y_3  (m11_port_y_3[2:0]    ), //o
    .clk       (clk                  ), //i
    .reset     (reset                )  //i
  );
  Multiplication_TI m12 (
    .port_x0_0 (t4_xor_port_y_0[2:0] ), //i
    .port_x0_1 (t4_xor_port_y_1[2:0] ), //i
    .port_x0_2 (t4_xor_port_y_2[2:0] ), //i
    .port_x0_3 (t4_xor_port_y_3[2:0] ), //i
    .port_x1_0 (t27_xor_port_y_0[2:0]), //i
    .port_x1_1 (t27_xor_port_y_1[2:0]), //i
    .port_x1_2 (t27_xor_port_y_2[2:0]), //i
    .port_x1_3 (t27_xor_port_y_3[2:0]), //i
    .port_y_0  (m12_port_y_0[2:0]    ), //o
    .port_y_1  (m12_port_y_1[2:0]    ), //o
    .port_y_2  (m12_port_y_2[2:0]    ), //o
    .port_y_3  (m12_port_y_3[2:0]    ), //o
    .clk       (clk                  ), //i
    .reset     (reset                )  //i
  );
  Multiplication_TI m14 (
    .port_x0_0 (t2_xor_port_y_0[2:0] ), //i
    .port_x0_1 (t2_xor_port_y_1[2:0] ), //i
    .port_x0_2 (t2_xor_port_y_2[2:0] ), //i
    .port_x0_3 (t2_xor_port_y_3[2:0] ), //i
    .port_x1_0 (t10_xor_port_y_0[2:0]), //i
    .port_x1_1 (t10_xor_port_y_1[2:0]), //i
    .port_x1_2 (t10_xor_port_y_2[2:0]), //i
    .port_x1_3 (t10_xor_port_y_3[2:0]), //i
    .port_y_0  (m14_port_y_0[2:0]    ), //o
    .port_y_1  (m14_port_y_1[2:0]    ), //o
    .port_y_2  (m14_port_y_2[2:0]    ), //o
    .port_y_3  (m14_port_y_3[2:0]    ), //o
    .clk       (clk                  ), //i
    .reset     (reset                )  //i
  );
  Addition_TI m3_xor (
    .port_x0_0 (t14_0[2:0]          ), //i
    .port_x0_1 (t14_1[2:0]          ), //i
    .port_x0_2 (t14_2[2:0]          ), //i
    .port_x0_3 (t14_3[2:0]          ), //i
    .port_x1_0 (m1_port_y_0[2:0]    ), //i
    .port_x1_1 (m1_port_y_1[2:0]    ), //i
    .port_x1_2 (m1_port_y_2[2:0]    ), //i
    .port_x1_3 (m1_port_y_3[2:0]    ), //i
    .port_y_0  (m3_xor_port_y_0[2:0]), //o
    .port_y_1  (m3_xor_port_y_1[2:0]), //o
    .port_y_2  (m3_xor_port_y_2[2:0]), //o
    .port_y_3  (m3_xor_port_y_3[2:0])  //o
  );
  Addition_TI m5_xor (
    .port_x0_0 (m4_port_y_0[2:0]    ), //i
    .port_x0_1 (m4_port_y_1[2:0]    ), //i
    .port_x0_2 (m4_port_y_2[2:0]    ), //i
    .port_x0_3 (m4_port_y_3[2:0]    ), //i
    .port_x1_0 (m1_port_y_0[2:0]    ), //i
    .port_x1_1 (m1_port_y_1[2:0]    ), //i
    .port_x1_2 (m1_port_y_2[2:0]    ), //i
    .port_x1_3 (m1_port_y_3[2:0]    ), //i
    .port_y_0  (m5_xor_port_y_0[2:0]), //o
    .port_y_1  (m5_xor_port_y_1[2:0]), //o
    .port_y_2  (m5_xor_port_y_2[2:0]), //o
    .port_y_3  (m5_xor_port_y_3[2:0])  //o
  );
  Addition_TI m8_xor (
    .port_x0_0 (t26_0[2:0]          ), //i
    .port_x0_1 (t26_1[2:0]          ), //i
    .port_x0_2 (t26_2[2:0]          ), //i
    .port_x0_3 (t26_3[2:0]          ), //i
    .port_x1_0 (m6_port_y_0[2:0]    ), //i
    .port_x1_1 (m6_port_y_1[2:0]    ), //i
    .port_x1_2 (m6_port_y_2[2:0]    ), //i
    .port_x1_3 (m6_port_y_3[2:0]    ), //i
    .port_y_0  (m8_xor_port_y_0[2:0]), //o
    .port_y_1  (m8_xor_port_y_1[2:0]), //o
    .port_y_2  (m8_xor_port_y_2[2:0]), //o
    .port_y_3  (m8_xor_port_y_3[2:0])  //o
  );
  Addition_TI m10_xor (
    .port_x0_0 (m9_port_y_0[2:0]     ), //i
    .port_x0_1 (m9_port_y_1[2:0]     ), //i
    .port_x0_2 (m9_port_y_2[2:0]     ), //i
    .port_x0_3 (m9_port_y_3[2:0]     ), //i
    .port_x1_0 (m6_port_y_0[2:0]     ), //i
    .port_x1_1 (m6_port_y_1[2:0]     ), //i
    .port_x1_2 (m6_port_y_2[2:0]     ), //i
    .port_x1_3 (m6_port_y_3[2:0]     ), //i
    .port_y_0  (m10_xor_port_y_0[2:0]), //o
    .port_y_1  (m10_xor_port_y_1[2:0]), //o
    .port_y_2  (m10_xor_port_y_2[2:0]), //o
    .port_y_3  (m10_xor_port_y_3[2:0])  //o
  );
  Addition_TI m13_xor (
    .port_x0_0 (m12_port_y_0[2:0]    ), //i
    .port_x0_1 (m12_port_y_1[2:0]    ), //i
    .port_x0_2 (m12_port_y_2[2:0]    ), //i
    .port_x0_3 (m12_port_y_3[2:0]    ), //i
    .port_x1_0 (m11_port_y_0[2:0]    ), //i
    .port_x1_1 (m11_port_y_1[2:0]    ), //i
    .port_x1_2 (m11_port_y_2[2:0]    ), //i
    .port_x1_3 (m11_port_y_3[2:0]    ), //i
    .port_y_0  (m13_xor_port_y_0[2:0]), //o
    .port_y_1  (m13_xor_port_y_1[2:0]), //o
    .port_y_2  (m13_xor_port_y_2[2:0]), //o
    .port_y_3  (m13_xor_port_y_3[2:0])  //o
  );
  Addition_TI m15_xor (
    .port_x0_0 (m14_port_y_0[2:0]    ), //i
    .port_x0_1 (m14_port_y_1[2:0]    ), //i
    .port_x0_2 (m14_port_y_2[2:0]    ), //i
    .port_x0_3 (m14_port_y_3[2:0]    ), //i
    .port_x1_0 (m11_port_y_0[2:0]    ), //i
    .port_x1_1 (m11_port_y_1[2:0]    ), //i
    .port_x1_2 (m11_port_y_2[2:0]    ), //i
    .port_x1_3 (m11_port_y_3[2:0]    ), //i
    .port_y_0  (m15_xor_port_y_0[2:0]), //o
    .port_y_1  (m15_xor_port_y_1[2:0]), //o
    .port_y_2  (m15_xor_port_y_2[2:0]), //o
    .port_y_3  (m15_xor_port_y_3[2:0])  //o
  );
  Addition_TI m16_xor (
    .port_x0_0 (m3_xor_port_y_0[2:0] ), //i
    .port_x0_1 (m3_xor_port_y_1[2:0] ), //i
    .port_x0_2 (m3_xor_port_y_2[2:0] ), //i
    .port_x0_3 (m3_xor_port_y_3[2:0] ), //i
    .port_x1_0 (m2_port_y_0[2:0]     ), //i
    .port_x1_1 (m2_port_y_1[2:0]     ), //i
    .port_x1_2 (m2_port_y_2[2:0]     ), //i
    .port_x1_3 (m2_port_y_3[2:0]     ), //i
    .port_y_0  (m16_xor_port_y_0[2:0]), //o
    .port_y_1  (m16_xor_port_y_1[2:0]), //o
    .port_y_2  (m16_xor_port_y_2[2:0]), //o
    .port_y_3  (m16_xor_port_y_3[2:0])  //o
  );
  Addition_TI m17_xor (
    .port_x0_0 (m5_xor_port_y_0[2:0] ), //i
    .port_x0_1 (m5_xor_port_y_1[2:0] ), //i
    .port_x0_2 (m5_xor_port_y_2[2:0] ), //i
    .port_x0_3 (m5_xor_port_y_3[2:0] ), //i
    .port_x1_0 (t24_0[2:0]           ), //i
    .port_x1_1 (t24_1[2:0]           ), //i
    .port_x1_2 (t24_2[2:0]           ), //i
    .port_x1_3 (t24_3[2:0]           ), //i
    .port_y_0  (m17_xor_port_y_0[2:0]), //o
    .port_y_1  (m17_xor_port_y_1[2:0]), //o
    .port_y_2  (m17_xor_port_y_2[2:0]), //o
    .port_y_3  (m17_xor_port_y_3[2:0])  //o
  );
  Addition_TI m18_xor (
    .port_x0_0 (m8_xor_port_y_0[2:0] ), //i
    .port_x0_1 (m8_xor_port_y_1[2:0] ), //i
    .port_x0_2 (m8_xor_port_y_2[2:0] ), //i
    .port_x0_3 (m8_xor_port_y_3[2:0] ), //i
    .port_x1_0 (m7_port_y_0[2:0]     ), //i
    .port_x1_1 (m7_port_y_1[2:0]     ), //i
    .port_x1_2 (m7_port_y_2[2:0]     ), //i
    .port_x1_3 (m7_port_y_3[2:0]     ), //i
    .port_y_0  (m18_xor_port_y_0[2:0]), //o
    .port_y_1  (m18_xor_port_y_1[2:0]), //o
    .port_y_2  (m18_xor_port_y_2[2:0]), //o
    .port_y_3  (m18_xor_port_y_3[2:0])  //o
  );
  Addition_TI m19_xor (
    .port_x0_0 (m10_xor_port_y_0[2:0]), //i
    .port_x0_1 (m10_xor_port_y_1[2:0]), //i
    .port_x0_2 (m10_xor_port_y_2[2:0]), //i
    .port_x0_3 (m10_xor_port_y_3[2:0]), //i
    .port_x1_0 (m15_xor_port_y_0[2:0]), //i
    .port_x1_1 (m15_xor_port_y_1[2:0]), //i
    .port_x1_2 (m15_xor_port_y_2[2:0]), //i
    .port_x1_3 (m15_xor_port_y_3[2:0]), //i
    .port_y_0  (m19_xor_port_y_0[2:0]), //o
    .port_y_1  (m19_xor_port_y_1[2:0]), //o
    .port_y_2  (m19_xor_port_y_2[2:0]), //o
    .port_y_3  (m19_xor_port_y_3[2:0])  //o
  );
  Addition_TI m20_xor (
    .port_x0_0 (m16_xor_port_y_0[2:0]), //i
    .port_x0_1 (m16_xor_port_y_1[2:0]), //i
    .port_x0_2 (m16_xor_port_y_2[2:0]), //i
    .port_x0_3 (m16_xor_port_y_3[2:0]), //i
    .port_x1_0 (m13_xor_port_y_0[2:0]), //i
    .port_x1_1 (m13_xor_port_y_1[2:0]), //i
    .port_x1_2 (m13_xor_port_y_2[2:0]), //i
    .port_x1_3 (m13_xor_port_y_3[2:0]), //i
    .port_y_0  (m20_xor_port_y_0[2:0]), //o
    .port_y_1  (m20_xor_port_y_1[2:0]), //o
    .port_y_2  (m20_xor_port_y_2[2:0]), //o
    .port_y_3  (m20_xor_port_y_3[2:0])  //o
  );
  Addition_TI m21_xor (
    .port_x0_0 (m17_xor_port_y_0[2:0]), //i
    .port_x0_1 (m17_xor_port_y_1[2:0]), //i
    .port_x0_2 (m17_xor_port_y_2[2:0]), //i
    .port_x0_3 (m17_xor_port_y_3[2:0]), //i
    .port_x1_0 (m15_xor_port_y_0[2:0]), //i
    .port_x1_1 (m15_xor_port_y_1[2:0]), //i
    .port_x1_2 (m15_xor_port_y_2[2:0]), //i
    .port_x1_3 (m15_xor_port_y_3[2:0]), //i
    .port_y_0  (m21_xor_port_y_0[2:0]), //o
    .port_y_1  (m21_xor_port_y_1[2:0]), //o
    .port_y_2  (m21_xor_port_y_2[2:0]), //o
    .port_y_3  (m21_xor_port_y_3[2:0])  //o
  );
  Addition_TI m22_xor (
    .port_x0_0 (m18_xor_port_y_0[2:0]), //i
    .port_x0_1 (m18_xor_port_y_1[2:0]), //i
    .port_x0_2 (m18_xor_port_y_2[2:0]), //i
    .port_x0_3 (m18_xor_port_y_3[2:0]), //i
    .port_x1_0 (m13_xor_port_y_0[2:0]), //i
    .port_x1_1 (m13_xor_port_y_1[2:0]), //i
    .port_x1_2 (m13_xor_port_y_2[2:0]), //i
    .port_x1_3 (m13_xor_port_y_3[2:0]), //i
    .port_y_0  (m22_xor_port_y_0[2:0]), //o
    .port_y_1  (m22_xor_port_y_1[2:0]), //o
    .port_y_2  (m22_xor_port_y_2[2:0]), //o
    .port_y_3  (m22_xor_port_y_3[2:0])  //o
  );
  Addition_TI m23_xor (
    .port_x0_0 (m19_xor_port_y_0[2:0]), //i
    .port_x0_1 (m19_xor_port_y_1[2:0]), //i
    .port_x0_2 (m19_xor_port_y_2[2:0]), //i
    .port_x0_3 (m19_xor_port_y_3[2:0]), //i
    .port_x1_0 (t25_0[2:0]           ), //i
    .port_x1_1 (t25_1[2:0]           ), //i
    .port_x1_2 (t25_2[2:0]           ), //i
    .port_x1_3 (t25_3[2:0]           ), //i
    .port_y_0  (m23_xor_port_y_0[2:0]), //o
    .port_y_1  (m23_xor_port_y_1[2:0]), //o
    .port_y_2  (m23_xor_port_y_2[2:0]), //o
    .port_y_3  (m23_xor_port_y_3[2:0])  //o
  );
  Addition_TI m24_xor (
    .port_x0_0 (m22_xor_port_y_0[2:0]), //i
    .port_x0_1 (m22_xor_port_y_1[2:0]), //i
    .port_x0_2 (m22_xor_port_y_2[2:0]), //i
    .port_x0_3 (m22_xor_port_y_3[2:0]), //i
    .port_x1_0 (m23_xor_port_y_0[2:0]), //i
    .port_x1_1 (m23_xor_port_y_1[2:0]), //i
    .port_x1_2 (m23_xor_port_y_2[2:0]), //i
    .port_x1_3 (m23_xor_port_y_3[2:0]), //i
    .port_y_0  (m24_xor_port_y_0[2:0]), //o
    .port_y_1  (m24_xor_port_y_1[2:0]), //o
    .port_y_2  (m24_xor_port_y_2[2:0]), //o
    .port_y_3  (m24_xor_port_y_3[2:0])  //o
  );
  Multiplication_TI m25 (
    .port_x0_0 (m22_xor_port_y_0[2:0]), //i
    .port_x0_1 (m22_xor_port_y_1[2:0]), //i
    .port_x0_2 (m22_xor_port_y_2[2:0]), //i
    .port_x0_3 (m22_xor_port_y_3[2:0]), //i
    .port_x1_0 (m20_xor_port_y_0[2:0]), //i
    .port_x1_1 (m20_xor_port_y_1[2:0]), //i
    .port_x1_2 (m20_xor_port_y_2[2:0]), //i
    .port_x1_3 (m20_xor_port_y_3[2:0]), //i
    .port_y_0  (m25_port_y_0[2:0]    ), //o
    .port_y_1  (m25_port_y_1[2:0]    ), //o
    .port_y_2  (m25_port_y_2[2:0]    ), //o
    .port_y_3  (m25_port_y_3[2:0]    ), //o
    .clk       (clk                  ), //i
    .reset     (reset                )  //i
  );
  Addition_TI m27_xor (
    .port_x0_0 (m20_xor_port_y_0[2:0]), //i
    .port_x0_1 (m20_xor_port_y_1[2:0]), //i
    .port_x0_2 (m20_xor_port_y_2[2:0]), //i
    .port_x0_3 (m20_xor_port_y_3[2:0]), //i
    .port_x1_0 (m21_xor_port_y_0[2:0]), //i
    .port_x1_1 (m21_xor_port_y_1[2:0]), //i
    .port_x1_2 (m21_xor_port_y_2[2:0]), //i
    .port_x1_3 (m21_xor_port_y_3[2:0]), //i
    .port_y_0  (m27_xor_port_y_0[2:0]), //o
    .port_y_1  (m27_xor_port_y_1[2:0]), //o
    .port_y_2  (m27_xor_port_y_2[2:0]), //o
    .port_y_3  (m27_xor_port_y_3[2:0])  //o
  );
  Multiplication_TI m31 (
    .port_x0_0 (m20_xor_port_y_0[2:0]), //i
    .port_x0_1 (m20_xor_port_y_1[2:0]), //i
    .port_x0_2 (m20_xor_port_y_2[2:0]), //i
    .port_x0_3 (m20_xor_port_y_3[2:0]), //i
    .port_x1_0 (m23_xor_port_y_0[2:0]), //i
    .port_x1_1 (m23_xor_port_y_1[2:0]), //i
    .port_x1_2 (m23_xor_port_y_2[2:0]), //i
    .port_x1_3 (m23_xor_port_y_3[2:0]), //i
    .port_y_0  (m31_port_y_0[2:0]    ), //o
    .port_y_1  (m31_port_y_1[2:0]    ), //o
    .port_y_2  (m31_port_y_2[2:0]    ), //o
    .port_y_3  (m31_port_y_3[2:0]    ), //o
    .clk       (clk                  ), //i
    .reset     (reset                )  //i
  );
  Multiplication_TI m34 (
    .port_x0_0 (m21_xor_port_y_0[2:0]), //i
    .port_x0_1 (m21_xor_port_y_1[2:0]), //i
    .port_x0_2 (m21_xor_port_y_2[2:0]), //i
    .port_x0_3 (m21_xor_port_y_3[2:0]), //i
    .port_x1_0 (m22_xor_port_y_0[2:0]), //i
    .port_x1_1 (m22_xor_port_y_1[2:0]), //i
    .port_x1_2 (m22_xor_port_y_2[2:0]), //i
    .port_x1_3 (m22_xor_port_y_3[2:0]), //i
    .port_y_0  (m34_port_y_0[2:0]    ), //o
    .port_y_1  (m34_port_y_1[2:0]    ), //o
    .port_y_2  (m34_port_y_2[2:0]    ), //o
    .port_y_3  (m34_port_y_3[2:0]    ), //o
    .clk       (clk                  ), //i
    .reset     (reset                )  //i
  );
  Addition_TI m26_xor (
    .port_x0_0 (m21_0[2:0]           ), //i
    .port_x0_1 (m21_1[2:0]           ), //i
    .port_x0_2 (m21_2[2:0]           ), //i
    .port_x0_3 (m21_3[2:0]           ), //i
    .port_x1_0 (m25_port_y_0[2:0]    ), //i
    .port_x1_1 (m25_port_y_1[2:0]    ), //i
    .port_x1_2 (m25_port_y_2[2:0]    ), //i
    .port_x1_3 (m25_port_y_3[2:0]    ), //i
    .port_y_0  (m26_xor_port_y_0[2:0]), //o
    .port_y_1  (m26_xor_port_y_1[2:0]), //o
    .port_y_2  (m26_xor_port_y_2[2:0]), //o
    .port_y_3  (m26_xor_port_y_3[2:0])  //o
  );
  Addition_TI m28_xor (
    .port_x0_0 (m23_0[2:0]           ), //i
    .port_x0_1 (m23_1[2:0]           ), //i
    .port_x0_2 (m23_2[2:0]           ), //i
    .port_x0_3 (m23_3[2:0]           ), //i
    .port_x1_0 (m25_port_y_0[2:0]    ), //i
    .port_x1_1 (m25_port_y_1[2:0]    ), //i
    .port_x1_2 (m25_port_y_2[2:0]    ), //i
    .port_x1_3 (m25_port_y_3[2:0]    ), //i
    .port_y_0  (m28_xor_port_y_0[2:0]), //o
    .port_y_1  (m28_xor_port_y_1[2:0]), //o
    .port_y_2  (m28_xor_port_y_2[2:0]), //o
    .port_y_3  (m28_xor_port_y_3[2:0])  //o
  );
  Multiplication_TI m29 (
    .port_x0_0 (m28_xor_port_y_0[2:0]), //i
    .port_x0_1 (m28_xor_port_y_1[2:0]), //i
    .port_x0_2 (m28_xor_port_y_2[2:0]), //i
    .port_x0_3 (m28_xor_port_y_3[2:0]), //i
    .port_x1_0 (m27_0[2:0]           ), //i
    .port_x1_1 (m27_1[2:0]           ), //i
    .port_x1_2 (m27_2[2:0]           ), //i
    .port_x1_3 (m27_3[2:0]           ), //i
    .port_y_0  (m29_port_y_0[2:0]    ), //o
    .port_y_1  (m29_port_y_1[2:0]    ), //o
    .port_y_2  (m29_port_y_2[2:0]    ), //o
    .port_y_3  (m29_port_y_3[2:0]    ), //o
    .clk       (clk                  ), //i
    .reset     (reset                )  //i
  );
  Multiplication_TI m30 (
    .port_x0_0 (m26_xor_port_y_0[2:0]), //i
    .port_x0_1 (m26_xor_port_y_1[2:0]), //i
    .port_x0_2 (m26_xor_port_y_2[2:0]), //i
    .port_x0_3 (m26_xor_port_y_3[2:0]), //i
    .port_x1_0 (m24_0[2:0]           ), //i
    .port_x1_1 (m24_1[2:0]           ), //i
    .port_x1_2 (m24_2[2:0]           ), //i
    .port_x1_3 (m24_3[2:0]           ), //i
    .port_y_0  (m30_port_y_0[2:0]    ), //o
    .port_y_1  (m30_port_y_1[2:0]    ), //o
    .port_y_2  (m30_port_y_2[2:0]    ), //o
    .port_y_3  (m30_port_y_3[2:0]    ), //o
    .clk       (clk                  ), //i
    .reset     (reset                )  //i
  );
  Multiplication_TI m32 (
    .port_x0_0 (m27_0[2:0]       ), //i
    .port_x0_1 (m27_1[2:0]       ), //i
    .port_x0_2 (m27_2[2:0]       ), //i
    .port_x0_3 (m27_3[2:0]       ), //i
    .port_x1_0 (m31_port_y_0[2:0]), //i
    .port_x1_1 (m31_port_y_1[2:0]), //i
    .port_x1_2 (m31_port_y_2[2:0]), //i
    .port_x1_3 (m31_port_y_3[2:0]), //i
    .port_y_0  (m32_port_y_0[2:0]), //o
    .port_y_1  (m32_port_y_1[2:0]), //o
    .port_y_2  (m32_port_y_2[2:0]), //o
    .port_y_3  (m32_port_y_3[2:0]), //o
    .clk       (clk              ), //i
    .reset     (reset            )  //i
  );
  Addition_TI m33_xor (
    .port_x0_0 (m27_0[2:0]           ), //i
    .port_x0_1 (m27_1[2:0]           ), //i
    .port_x0_2 (m27_2[2:0]           ), //i
    .port_x0_3 (m27_3[2:0]           ), //i
    .port_x1_0 (m25_port_y_0[2:0]    ), //i
    .port_x1_1 (m25_port_y_1[2:0]    ), //i
    .port_x1_2 (m25_port_y_2[2:0]    ), //i
    .port_x1_3 (m25_port_y_3[2:0]    ), //i
    .port_y_0  (m33_xor_port_y_0[2:0]), //o
    .port_y_1  (m33_xor_port_y_1[2:0]), //o
    .port_y_2  (m33_xor_port_y_2[2:0]), //o
    .port_y_3  (m33_xor_port_y_3[2:0])  //o
  );
  Multiplication_TI m35 (
    .port_x0_0 (m24_0[2:0]       ), //i
    .port_x0_1 (m24_1[2:0]       ), //i
    .port_x0_2 (m24_2[2:0]       ), //i
    .port_x0_3 (m24_3[2:0]       ), //i
    .port_x1_0 (m34_port_y_0[2:0]), //i
    .port_x1_1 (m34_port_y_1[2:0]), //i
    .port_x1_2 (m34_port_y_2[2:0]), //i
    .port_x1_3 (m34_port_y_3[2:0]), //i
    .port_y_0  (m35_port_y_0[2:0]), //o
    .port_y_1  (m35_port_y_1[2:0]), //o
    .port_y_2  (m35_port_y_2[2:0]), //o
    .port_y_3  (m35_port_y_3[2:0]), //o
    .clk       (clk              ), //i
    .reset     (reset            )  //i
  );
  Addition_TI m36_xor (
    .port_x0_0 (m24_0[2:0]           ), //i
    .port_x0_1 (m24_1[2:0]           ), //i
    .port_x0_2 (m24_2[2:0]           ), //i
    .port_x0_3 (m24_3[2:0]           ), //i
    .port_x1_0 (m25_port_y_0[2:0]    ), //i
    .port_x1_1 (m25_port_y_1[2:0]    ), //i
    .port_x1_2 (m25_port_y_2[2:0]    ), //i
    .port_x1_3 (m25_port_y_3[2:0]    ), //i
    .port_y_0  (m36_xor_port_y_0[2:0]), //o
    .port_y_1  (m36_xor_port_y_1[2:0]), //o
    .port_y_2  (m36_xor_port_y_2[2:0]), //o
    .port_y_3  (m36_xor_port_y_3[2:0])  //o
  );
  Addition_TI m37_xor (
    .port_x0_0 (m21_1_0[2:0]         ), //i
    .port_x0_1 (m21_1_1[2:0]         ), //i
    .port_x0_2 (m21_1_2[2:0]         ), //i
    .port_x0_3 (m21_1_3[2:0]         ), //i
    .port_x1_0 (m29_port_y_0[2:0]    ), //i
    .port_x1_1 (m29_port_y_1[2:0]    ), //i
    .port_x1_2 (m29_port_y_2[2:0]    ), //i
    .port_x1_3 (m29_port_y_3[2:0]    ), //i
    .port_y_0  (m37_xor_port_y_0[2:0]), //o
    .port_y_1  (m37_xor_port_y_1[2:0]), //o
    .port_y_2  (m37_xor_port_y_2[2:0]), //o
    .port_y_3  (m37_xor_port_y_3[2:0])  //o
  );
  Addition_TI m38_xor (
    .port_x0_0 (m32_port_y_0[2:0]    ), //i
    .port_x0_1 (m32_port_y_1[2:0]    ), //i
    .port_x0_2 (m32_port_y_2[2:0]    ), //i
    .port_x0_3 (m32_port_y_3[2:0]    ), //i
    .port_x1_0 (m33_0[2:0]           ), //i
    .port_x1_1 (m33_1[2:0]           ), //i
    .port_x1_2 (m33_2[2:0]           ), //i
    .port_x1_3 (m33_3[2:0]           ), //i
    .port_y_0  (m38_xor_port_y_0[2:0]), //o
    .port_y_1  (m38_xor_port_y_1[2:0]), //o
    .port_y_2  (m38_xor_port_y_2[2:0]), //o
    .port_y_3  (m38_xor_port_y_3[2:0])  //o
  );
  Addition_TI m39_xor (
    .port_x0_0 (m23_1_0[2:0]         ), //i
    .port_x0_1 (m23_1_1[2:0]         ), //i
    .port_x0_2 (m23_1_2[2:0]         ), //i
    .port_x0_3 (m23_1_3[2:0]         ), //i
    .port_x1_0 (m30_port_y_0[2:0]    ), //i
    .port_x1_1 (m30_port_y_1[2:0]    ), //i
    .port_x1_2 (m30_port_y_2[2:0]    ), //i
    .port_x1_3 (m30_port_y_3[2:0]    ), //i
    .port_y_0  (m39_xor_port_y_0[2:0]), //o
    .port_y_1  (m39_xor_port_y_1[2:0]), //o
    .port_y_2  (m39_xor_port_y_2[2:0]), //o
    .port_y_3  (m39_xor_port_y_3[2:0])  //o
  );
  Addition_TI m40_xor (
    .port_x0_0 (m35_port_y_0[2:0]    ), //i
    .port_x0_1 (m35_port_y_1[2:0]    ), //i
    .port_x0_2 (m35_port_y_2[2:0]    ), //i
    .port_x0_3 (m35_port_y_3[2:0]    ), //i
    .port_x1_0 (m36_0[2:0]           ), //i
    .port_x1_1 (m36_1[2:0]           ), //i
    .port_x1_2 (m36_2[2:0]           ), //i
    .port_x1_3 (m36_3[2:0]           ), //i
    .port_y_0  (m40_xor_port_y_0[2:0]), //o
    .port_y_1  (m40_xor_port_y_1[2:0]), //o
    .port_y_2  (m40_xor_port_y_2[2:0]), //o
    .port_y_3  (m40_xor_port_y_3[2:0])  //o
  );
  Addition_TI m41_xor (
    .port_x0_0 (m38_xor_port_y_0[2:0]), //i
    .port_x0_1 (m38_xor_port_y_1[2:0]), //i
    .port_x0_2 (m38_xor_port_y_2[2:0]), //i
    .port_x0_3 (m38_xor_port_y_3[2:0]), //i
    .port_x1_0 (m40_xor_port_y_0[2:0]), //i
    .port_x1_1 (m40_xor_port_y_1[2:0]), //i
    .port_x1_2 (m40_xor_port_y_2[2:0]), //i
    .port_x1_3 (m40_xor_port_y_3[2:0]), //i
    .port_y_0  (m41_xor_port_y_0[2:0]), //o
    .port_y_1  (m41_xor_port_y_1[2:0]), //o
    .port_y_2  (m41_xor_port_y_2[2:0]), //o
    .port_y_3  (m41_xor_port_y_3[2:0])  //o
  );
  Addition_TI m42_xor (
    .port_x0_0 (m37_xor_port_y_0[2:0]), //i
    .port_x0_1 (m37_xor_port_y_1[2:0]), //i
    .port_x0_2 (m37_xor_port_y_2[2:0]), //i
    .port_x0_3 (m37_xor_port_y_3[2:0]), //i
    .port_x1_0 (m39_xor_port_y_0[2:0]), //i
    .port_x1_1 (m39_xor_port_y_1[2:0]), //i
    .port_x1_2 (m39_xor_port_y_2[2:0]), //i
    .port_x1_3 (m39_xor_port_y_3[2:0]), //i
    .port_y_0  (m42_xor_port_y_0[2:0]), //o
    .port_y_1  (m42_xor_port_y_1[2:0]), //o
    .port_y_2  (m42_xor_port_y_2[2:0]), //o
    .port_y_3  (m42_xor_port_y_3[2:0])  //o
  );
  Addition_TI m43_xor (
    .port_x0_0 (m37_xor_port_y_0[2:0]), //i
    .port_x0_1 (m37_xor_port_y_1[2:0]), //i
    .port_x0_2 (m37_xor_port_y_2[2:0]), //i
    .port_x0_3 (m37_xor_port_y_3[2:0]), //i
    .port_x1_0 (m38_xor_port_y_0[2:0]), //i
    .port_x1_1 (m38_xor_port_y_1[2:0]), //i
    .port_x1_2 (m38_xor_port_y_2[2:0]), //i
    .port_x1_3 (m38_xor_port_y_3[2:0]), //i
    .port_y_0  (m43_xor_port_y_0[2:0]), //o
    .port_y_1  (m43_xor_port_y_1[2:0]), //o
    .port_y_2  (m43_xor_port_y_2[2:0]), //o
    .port_y_3  (m43_xor_port_y_3[2:0])  //o
  );
  Addition_TI m44_xor (
    .port_x0_0 (m39_xor_port_y_0[2:0]), //i
    .port_x0_1 (m39_xor_port_y_1[2:0]), //i
    .port_x0_2 (m39_xor_port_y_2[2:0]), //i
    .port_x0_3 (m39_xor_port_y_3[2:0]), //i
    .port_x1_0 (m40_xor_port_y_0[2:0]), //i
    .port_x1_1 (m40_xor_port_y_1[2:0]), //i
    .port_x1_2 (m40_xor_port_y_2[2:0]), //i
    .port_x1_3 (m40_xor_port_y_3[2:0]), //i
    .port_y_0  (m44_xor_port_y_0[2:0]), //o
    .port_y_1  (m44_xor_port_y_1[2:0]), //o
    .port_y_2  (m44_xor_port_y_2[2:0]), //o
    .port_y_3  (m44_xor_port_y_3[2:0])  //o
  );
  Addition_TI m45_xor (
    .port_x0_0 (m42_xor_port_y_0[2:0]), //i
    .port_x0_1 (m42_xor_port_y_1[2:0]), //i
    .port_x0_2 (m42_xor_port_y_2[2:0]), //i
    .port_x0_3 (m42_xor_port_y_3[2:0]), //i
    .port_x1_0 (m41_xor_port_y_0[2:0]), //i
    .port_x1_1 (m41_xor_port_y_1[2:0]), //i
    .port_x1_2 (m41_xor_port_y_2[2:0]), //i
    .port_x1_3 (m41_xor_port_y_3[2:0]), //i
    .port_y_0  (m45_xor_port_y_0[2:0]), //o
    .port_y_1  (m45_xor_port_y_1[2:0]), //o
    .port_y_2  (m45_xor_port_y_2[2:0]), //o
    .port_y_3  (m45_xor_port_y_3[2:0])  //o
  );
  Multiplication_TI_noReg m46_mul (
    .port_x0_0 (m44_xor_port_y_0[2:0]), //i
    .port_x0_1 (m44_xor_port_y_1[2:0]), //i
    .port_x0_2 (m44_xor_port_y_2[2:0]), //i
    .port_x0_3 (m44_xor_port_y_3[2:0]), //i
    .port_x1_0 (t6_2_0[2:0]          ), //i
    .port_x1_1 (t6_2_1[2:0]          ), //i
    .port_x1_2 (t6_2_2[2:0]          ), //i
    .port_x1_3 (t6_2_3[2:0]          ), //i
    .port_y_0  (m46_mul_port_y_0[2:0]), //o
    .port_y_1  (m46_mul_port_y_1[2:0]), //o
    .port_y_2  (m46_mul_port_y_2[2:0]), //o
    .port_y_3  (m46_mul_port_y_3[2:0])  //o
  );
  Multiplication_TI_noReg m47_mul (
    .port_x0_0 (m40_xor_port_y_0[2:0]), //i
    .port_x0_1 (m40_xor_port_y_1[2:0]), //i
    .port_x0_2 (m40_xor_port_y_2[2:0]), //i
    .port_x0_3 (m40_xor_port_y_3[2:0]), //i
    .port_x1_0 (t8_2_0[2:0]          ), //i
    .port_x1_1 (t8_2_1[2:0]          ), //i
    .port_x1_2 (t8_2_2[2:0]          ), //i
    .port_x1_3 (t8_2_3[2:0]          ), //i
    .port_y_0  (m47_mul_port_y_0[2:0]), //o
    .port_y_1  (m47_mul_port_y_1[2:0]), //o
    .port_y_2  (m47_mul_port_y_2[2:0]), //o
    .port_y_3  (m47_mul_port_y_3[2:0])  //o
  );
  Multiplication_TI_noReg m48_mul (
    .port_x0_0 (m39_xor_port_y_0[2:0]), //i
    .port_x0_1 (m39_xor_port_y_1[2:0]), //i
    .port_x0_2 (m39_xor_port_y_2[2:0]), //i
    .port_x0_3 (m39_xor_port_y_3[2:0]), //i
    .port_x1_0 (x7_2_0[2:0]          ), //i
    .port_x1_1 (x7_2_1[2:0]          ), //i
    .port_x1_2 (x7_2_2[2:0]          ), //i
    .port_x1_3 (x7_2_3[2:0]          ), //i
    .port_y_0  (m48_mul_port_y_0[2:0]), //o
    .port_y_1  (m48_mul_port_y_1[2:0]), //o
    .port_y_2  (m48_mul_port_y_2[2:0]), //o
    .port_y_3  (m48_mul_port_y_3[2:0])  //o
  );
  Multiplication_TI_noReg m49_mul (
    .port_x0_0 (m43_xor_port_y_0[2:0]), //i
    .port_x0_1 (m43_xor_port_y_1[2:0]), //i
    .port_x0_2 (m43_xor_port_y_2[2:0]), //i
    .port_x0_3 (m43_xor_port_y_3[2:0]), //i
    .port_x1_0 (t16_1_0[2:0]         ), //i
    .port_x1_1 (t16_1_1[2:0]         ), //i
    .port_x1_2 (t16_1_2[2:0]         ), //i
    .port_x1_3 (t16_1_3[2:0]         ), //i
    .port_y_0  (m49_mul_port_y_0[2:0]), //o
    .port_y_1  (m49_mul_port_y_1[2:0]), //o
    .port_y_2  (m49_mul_port_y_2[2:0]), //o
    .port_y_3  (m49_mul_port_y_3[2:0])  //o
  );
  Multiplication_TI_noReg m50_mul (
    .port_x0_0 (m38_xor_port_y_0[2:0]), //i
    .port_x0_1 (m38_xor_port_y_1[2:0]), //i
    .port_x0_2 (m38_xor_port_y_2[2:0]), //i
    .port_x0_3 (m38_xor_port_y_3[2:0]), //i
    .port_x1_0 (t9_2_0[2:0]          ), //i
    .port_x1_1 (t9_2_1[2:0]          ), //i
    .port_x1_2 (t9_2_2[2:0]          ), //i
    .port_x1_3 (t9_2_3[2:0]          ), //i
    .port_y_0  (m50_mul_port_y_0[2:0]), //o
    .port_y_1  (m50_mul_port_y_1[2:0]), //o
    .port_y_2  (m50_mul_port_y_2[2:0]), //o
    .port_y_3  (m50_mul_port_y_3[2:0])  //o
  );
  Multiplication_TI_noReg m51_mul (
    .port_x0_0 (m37_xor_port_y_0[2:0]), //i
    .port_x0_1 (m37_xor_port_y_1[2:0]), //i
    .port_x0_2 (m37_xor_port_y_2[2:0]), //i
    .port_x0_3 (m37_xor_port_y_3[2:0]), //i
    .port_x1_0 (t17_2_0[2:0]         ), //i
    .port_x1_1 (t17_2_1[2:0]         ), //i
    .port_x1_2 (t17_2_2[2:0]         ), //i
    .port_x1_3 (t17_2_3[2:0]         ), //i
    .port_y_0  (m51_mul_port_y_0[2:0]), //o
    .port_y_1  (m51_mul_port_y_1[2:0]), //o
    .port_y_2  (m51_mul_port_y_2[2:0]), //o
    .port_y_3  (m51_mul_port_y_3[2:0])  //o
  );
  Multiplication_TI_noReg m52_mul (
    .port_x0_0 (m42_xor_port_y_0[2:0]), //i
    .port_x0_1 (m42_xor_port_y_1[2:0]), //i
    .port_x0_2 (m42_xor_port_y_2[2:0]), //i
    .port_x0_3 (m42_xor_port_y_3[2:0]), //i
    .port_x1_0 (t15_2_0[2:0]         ), //i
    .port_x1_1 (t15_2_1[2:0]         ), //i
    .port_x1_2 (t15_2_2[2:0]         ), //i
    .port_x1_3 (t15_2_3[2:0]         ), //i
    .port_y_0  (m52_mul_port_y_0[2:0]), //o
    .port_y_1  (m52_mul_port_y_1[2:0]), //o
    .port_y_2  (m52_mul_port_y_2[2:0]), //o
    .port_y_3  (m52_mul_port_y_3[2:0])  //o
  );
  Multiplication_TI_noReg m53_mul (
    .port_x0_0 (m45_xor_port_y_0[2:0]), //i
    .port_x0_1 (m45_xor_port_y_1[2:0]), //i
    .port_x0_2 (m45_xor_port_y_2[2:0]), //i
    .port_x0_3 (m45_xor_port_y_3[2:0]), //i
    .port_x1_0 (t27_2_0[2:0]         ), //i
    .port_x1_1 (t27_2_1[2:0]         ), //i
    .port_x1_2 (t27_2_2[2:0]         ), //i
    .port_x1_3 (t27_2_3[2:0]         ), //i
    .port_y_0  (m53_mul_port_y_0[2:0]), //o
    .port_y_1  (m53_mul_port_y_1[2:0]), //o
    .port_y_2  (m53_mul_port_y_2[2:0]), //o
    .port_y_3  (m53_mul_port_y_3[2:0])  //o
  );
  Multiplication_TI_noReg m54_mul (
    .port_x0_0 (m41_xor_port_y_0[2:0]), //i
    .port_x0_1 (m41_xor_port_y_1[2:0]), //i
    .port_x0_2 (m41_xor_port_y_2[2:0]), //i
    .port_x0_3 (m41_xor_port_y_3[2:0]), //i
    .port_x1_0 (t10_2_0[2:0]         ), //i
    .port_x1_1 (t10_2_1[2:0]         ), //i
    .port_x1_2 (t10_2_2[2:0]         ), //i
    .port_x1_3 (t10_2_3[2:0]         ), //i
    .port_y_0  (m54_mul_port_y_0[2:0]), //o
    .port_y_1  (m54_mul_port_y_1[2:0]), //o
    .port_y_2  (m54_mul_port_y_2[2:0]), //o
    .port_y_3  (m54_mul_port_y_3[2:0])  //o
  );
  Multiplication_TI_noReg m55_mul (
    .port_x0_0 (m44_xor_port_y_0[2:0]), //i
    .port_x0_1 (m44_xor_port_y_1[2:0]), //i
    .port_x0_2 (m44_xor_port_y_2[2:0]), //i
    .port_x0_3 (m44_xor_port_y_3[2:0]), //i
    .port_x1_0 (t13_2_0[2:0]         ), //i
    .port_x1_1 (t13_2_1[2:0]         ), //i
    .port_x1_2 (t13_2_2[2:0]         ), //i
    .port_x1_3 (t13_2_3[2:0]         ), //i
    .port_y_0  (m55_mul_port_y_0[2:0]), //o
    .port_y_1  (m55_mul_port_y_1[2:0]), //o
    .port_y_2  (m55_mul_port_y_2[2:0]), //o
    .port_y_3  (m55_mul_port_y_3[2:0])  //o
  );
  Multiplication_TI_noReg m56_mul (
    .port_x0_0 (m40_xor_port_y_0[2:0]), //i
    .port_x0_1 (m40_xor_port_y_1[2:0]), //i
    .port_x0_2 (m40_xor_port_y_2[2:0]), //i
    .port_x0_3 (m40_xor_port_y_3[2:0]), //i
    .port_x1_0 (t23_2_0[2:0]         ), //i
    .port_x1_1 (t23_2_1[2:0]         ), //i
    .port_x1_2 (t23_2_2[2:0]         ), //i
    .port_x1_3 (t23_2_3[2:0]         ), //i
    .port_y_0  (m56_mul_port_y_0[2:0]), //o
    .port_y_1  (m56_mul_port_y_1[2:0]), //o
    .port_y_2  (m56_mul_port_y_2[2:0]), //o
    .port_y_3  (m56_mul_port_y_3[2:0])  //o
  );
  Multiplication_TI_noReg m57_mul (
    .port_x0_0 (m39_xor_port_y_0[2:0]), //i
    .port_x0_1 (m39_xor_port_y_1[2:0]), //i
    .port_x0_2 (m39_xor_port_y_2[2:0]), //i
    .port_x0_3 (m39_xor_port_y_3[2:0]), //i
    .port_x1_0 (t19_2_0[2:0]         ), //i
    .port_x1_1 (t19_2_1[2:0]         ), //i
    .port_x1_2 (t19_2_2[2:0]         ), //i
    .port_x1_3 (t19_2_3[2:0]         ), //i
    .port_y_0  (m57_mul_port_y_0[2:0]), //o
    .port_y_1  (m57_mul_port_y_1[2:0]), //o
    .port_y_2  (m57_mul_port_y_2[2:0]), //o
    .port_y_3  (m57_mul_port_y_3[2:0])  //o
  );
  Multiplication_TI_noReg m58_mul (
    .port_x0_0 (m43_xor_port_y_0[2:0]), //i
    .port_x0_1 (m43_xor_port_y_1[2:0]), //i
    .port_x0_2 (m43_xor_port_y_2[2:0]), //i
    .port_x0_3 (m43_xor_port_y_3[2:0]), //i
    .port_x1_0 (t3_2_0[2:0]          ), //i
    .port_x1_1 (t3_2_1[2:0]          ), //i
    .port_x1_2 (t3_2_2[2:0]          ), //i
    .port_x1_3 (t3_2_3[2:0]          ), //i
    .port_y_0  (m58_mul_port_y_0[2:0]), //o
    .port_y_1  (m58_mul_port_y_1[2:0]), //o
    .port_y_2  (m58_mul_port_y_2[2:0]), //o
    .port_y_3  (m58_mul_port_y_3[2:0])  //o
  );
  Multiplication_TI_noReg m59_mul (
    .port_x0_0 (m38_xor_port_y_0[2:0]), //i
    .port_x0_1 (m38_xor_port_y_1[2:0]), //i
    .port_x0_2 (m38_xor_port_y_2[2:0]), //i
    .port_x0_3 (m38_xor_port_y_3[2:0]), //i
    .port_x1_0 (t22_2_0[2:0]         ), //i
    .port_x1_1 (t22_2_1[2:0]         ), //i
    .port_x1_2 (t22_2_2[2:0]         ), //i
    .port_x1_3 (t22_2_3[2:0]         ), //i
    .port_y_0  (m59_mul_port_y_0[2:0]), //o
    .port_y_1  (m59_mul_port_y_1[2:0]), //o
    .port_y_2  (m59_mul_port_y_2[2:0]), //o
    .port_y_3  (m59_mul_port_y_3[2:0])  //o
  );
  Multiplication_TI_noReg m60_mul (
    .port_x0_0 (m37_xor_port_y_0[2:0]), //i
    .port_x0_1 (m37_xor_port_y_1[2:0]), //i
    .port_x0_2 (m37_xor_port_y_2[2:0]), //i
    .port_x0_3 (m37_xor_port_y_3[2:0]), //i
    .port_x1_0 (t20_2_0[2:0]         ), //i
    .port_x1_1 (t20_2_1[2:0]         ), //i
    .port_x1_2 (t20_2_2[2:0]         ), //i
    .port_x1_3 (t20_2_3[2:0]         ), //i
    .port_y_0  (m60_mul_port_y_0[2:0]), //o
    .port_y_1  (m60_mul_port_y_1[2:0]), //o
    .port_y_2  (m60_mul_port_y_2[2:0]), //o
    .port_y_3  (m60_mul_port_y_3[2:0])  //o
  );
  Multiplication_TI_noReg m61_mul (
    .port_x0_0 (m42_xor_port_y_0[2:0]), //i
    .port_x0_1 (m42_xor_port_y_1[2:0]), //i
    .port_x0_2 (m42_xor_port_y_2[2:0]), //i
    .port_x0_3 (m42_xor_port_y_3[2:0]), //i
    .port_x1_0 (t1_2_0[2:0]          ), //i
    .port_x1_1 (t1_2_1[2:0]          ), //i
    .port_x1_2 (t1_2_2[2:0]          ), //i
    .port_x1_3 (t1_2_3[2:0]          ), //i
    .port_y_0  (m61_mul_port_y_0[2:0]), //o
    .port_y_1  (m61_mul_port_y_1[2:0]), //o
    .port_y_2  (m61_mul_port_y_2[2:0]), //o
    .port_y_3  (m61_mul_port_y_3[2:0])  //o
  );
  Multiplication_TI_noReg m62_mul (
    .port_x0_0 (m45_xor_port_y_0[2:0]), //i
    .port_x0_1 (m45_xor_port_y_1[2:0]), //i
    .port_x0_2 (m45_xor_port_y_2[2:0]), //i
    .port_x0_3 (m45_xor_port_y_3[2:0]), //i
    .port_x1_0 (t4_2_0[2:0]          ), //i
    .port_x1_1 (t4_2_1[2:0]          ), //i
    .port_x1_2 (t4_2_2[2:0]          ), //i
    .port_x1_3 (t4_2_3[2:0]          ), //i
    .port_y_0  (m62_mul_port_y_0[2:0]), //o
    .port_y_1  (m62_mul_port_y_1[2:0]), //o
    .port_y_2  (m62_mul_port_y_2[2:0]), //o
    .port_y_3  (m62_mul_port_y_3[2:0])  //o
  );
  Multiplication_TI_noReg m63_mul (
    .port_x0_0 (m41_xor_port_y_0[2:0]), //i
    .port_x0_1 (m41_xor_port_y_1[2:0]), //i
    .port_x0_2 (m41_xor_port_y_2[2:0]), //i
    .port_x0_3 (m41_xor_port_y_3[2:0]), //i
    .port_x1_0 (t2_2_0[2:0]          ), //i
    .port_x1_1 (t2_2_1[2:0]          ), //i
    .port_x1_2 (t2_2_2[2:0]          ), //i
    .port_x1_3 (t2_2_3[2:0]          ), //i
    .port_y_0  (m63_mul_port_y_0[2:0]), //o
    .port_y_1  (m63_mul_port_y_1[2:0]), //o
    .port_y_2  (m63_mul_port_y_2[2:0]), //o
    .port_y_3  (m63_mul_port_y_3[2:0])  //o
  );
  Addition_TI l0_xor (
    .port_x0_0 (m61_mul_port_y_0[2:0]), //i
    .port_x0_1 (m61_mul_port_y_1[2:0]), //i
    .port_x0_2 (m61_mul_port_y_2[2:0]), //i
    .port_x0_3 (m61_mul_port_y_3[2:0]), //i
    .port_x1_0 (m62_mul_port_y_0[2:0]), //i
    .port_x1_1 (m62_mul_port_y_1[2:0]), //i
    .port_x1_2 (m62_mul_port_y_2[2:0]), //i
    .port_x1_3 (m62_mul_port_y_3[2:0]), //i
    .port_y_0  (l0_xor_port_y_0[2:0] ), //o
    .port_y_1  (l0_xor_port_y_1[2:0] ), //o
    .port_y_2  (l0_xor_port_y_2[2:0] ), //o
    .port_y_3  (l0_xor_port_y_3[2:0] )  //o
  );
  Addition_TI l1_xor (
    .port_x0_0 (m50_mul_port_y_0[2:0]), //i
    .port_x0_1 (m50_mul_port_y_1[2:0]), //i
    .port_x0_2 (m50_mul_port_y_2[2:0]), //i
    .port_x0_3 (m50_mul_port_y_3[2:0]), //i
    .port_x1_0 (m56_mul_port_y_0[2:0]), //i
    .port_x1_1 (m56_mul_port_y_1[2:0]), //i
    .port_x1_2 (m56_mul_port_y_2[2:0]), //i
    .port_x1_3 (m56_mul_port_y_3[2:0]), //i
    .port_y_0  (l1_xor_port_y_0[2:0] ), //o
    .port_y_1  (l1_xor_port_y_1[2:0] ), //o
    .port_y_2  (l1_xor_port_y_2[2:0] ), //o
    .port_y_3  (l1_xor_port_y_3[2:0] )  //o
  );
  Addition_TI l2_xor (
    .port_x0_0 (m46_mul_port_y_0[2:0]), //i
    .port_x0_1 (m46_mul_port_y_1[2:0]), //i
    .port_x0_2 (m46_mul_port_y_2[2:0]), //i
    .port_x0_3 (m46_mul_port_y_3[2:0]), //i
    .port_x1_0 (m48_mul_port_y_0[2:0]), //i
    .port_x1_1 (m48_mul_port_y_1[2:0]), //i
    .port_x1_2 (m48_mul_port_y_2[2:0]), //i
    .port_x1_3 (m48_mul_port_y_3[2:0]), //i
    .port_y_0  (l2_xor_port_y_0[2:0] ), //o
    .port_y_1  (l2_xor_port_y_1[2:0] ), //o
    .port_y_2  (l2_xor_port_y_2[2:0] ), //o
    .port_y_3  (l2_xor_port_y_3[2:0] )  //o
  );
  Addition_TI l3_xor (
    .port_x0_0 (m47_mul_port_y_0[2:0]), //i
    .port_x0_1 (m47_mul_port_y_1[2:0]), //i
    .port_x0_2 (m47_mul_port_y_2[2:0]), //i
    .port_x0_3 (m47_mul_port_y_3[2:0]), //i
    .port_x1_0 (m55_mul_port_y_0[2:0]), //i
    .port_x1_1 (m55_mul_port_y_1[2:0]), //i
    .port_x1_2 (m55_mul_port_y_2[2:0]), //i
    .port_x1_3 (m55_mul_port_y_3[2:0]), //i
    .port_y_0  (l3_xor_port_y_0[2:0] ), //o
    .port_y_1  (l3_xor_port_y_1[2:0] ), //o
    .port_y_2  (l3_xor_port_y_2[2:0] ), //o
    .port_y_3  (l3_xor_port_y_3[2:0] )  //o
  );
  Addition_TI l4_xor (
    .port_x0_0 (m54_mul_port_y_0[2:0]), //i
    .port_x0_1 (m54_mul_port_y_1[2:0]), //i
    .port_x0_2 (m54_mul_port_y_2[2:0]), //i
    .port_x0_3 (m54_mul_port_y_3[2:0]), //i
    .port_x1_0 (m58_mul_port_y_0[2:0]), //i
    .port_x1_1 (m58_mul_port_y_1[2:0]), //i
    .port_x1_2 (m58_mul_port_y_2[2:0]), //i
    .port_x1_3 (m58_mul_port_y_3[2:0]), //i
    .port_y_0  (l4_xor_port_y_0[2:0] ), //o
    .port_y_1  (l4_xor_port_y_1[2:0] ), //o
    .port_y_2  (l4_xor_port_y_2[2:0] ), //o
    .port_y_3  (l4_xor_port_y_3[2:0] )  //o
  );
  Addition_TI l5_xor (
    .port_x0_0 (m49_mul_port_y_0[2:0]), //i
    .port_x0_1 (m49_mul_port_y_1[2:0]), //i
    .port_x0_2 (m49_mul_port_y_2[2:0]), //i
    .port_x0_3 (m49_mul_port_y_3[2:0]), //i
    .port_x1_0 (m61_mul_port_y_0[2:0]), //i
    .port_x1_1 (m61_mul_port_y_1[2:0]), //i
    .port_x1_2 (m61_mul_port_y_2[2:0]), //i
    .port_x1_3 (m61_mul_port_y_3[2:0]), //i
    .port_y_0  (l5_xor_port_y_0[2:0] ), //o
    .port_y_1  (l5_xor_port_y_1[2:0] ), //o
    .port_y_2  (l5_xor_port_y_2[2:0] ), //o
    .port_y_3  (l5_xor_port_y_3[2:0] )  //o
  );
  Addition_TI l6_xor (
    .port_x0_0 (m62_mul_port_y_0[2:0]), //i
    .port_x0_1 (m62_mul_port_y_1[2:0]), //i
    .port_x0_2 (m62_mul_port_y_2[2:0]), //i
    .port_x0_3 (m62_mul_port_y_3[2:0]), //i
    .port_x1_0 (l5_xor_port_y_0[2:0] ), //i
    .port_x1_1 (l5_xor_port_y_1[2:0] ), //i
    .port_x1_2 (l5_xor_port_y_2[2:0] ), //i
    .port_x1_3 (l5_xor_port_y_3[2:0] ), //i
    .port_y_0  (l6_xor_port_y_0[2:0] ), //o
    .port_y_1  (l6_xor_port_y_1[2:0] ), //o
    .port_y_2  (l6_xor_port_y_2[2:0] ), //o
    .port_y_3  (l6_xor_port_y_3[2:0] )  //o
  );
  Addition_TI l7_xor (
    .port_x0_0 (m46_mul_port_y_0[2:0]), //i
    .port_x0_1 (m46_mul_port_y_1[2:0]), //i
    .port_x0_2 (m46_mul_port_y_2[2:0]), //i
    .port_x0_3 (m46_mul_port_y_3[2:0]), //i
    .port_x1_0 (l3_xor_port_y_0[2:0] ), //i
    .port_x1_1 (l3_xor_port_y_1[2:0] ), //i
    .port_x1_2 (l3_xor_port_y_2[2:0] ), //i
    .port_x1_3 (l3_xor_port_y_3[2:0] ), //i
    .port_y_0  (l7_xor_port_y_0[2:0] ), //o
    .port_y_1  (l7_xor_port_y_1[2:0] ), //o
    .port_y_2  (l7_xor_port_y_2[2:0] ), //o
    .port_y_3  (l7_xor_port_y_3[2:0] )  //o
  );
  Addition_TI l8_xor (
    .port_x0_0 (m51_mul_port_y_0[2:0]), //i
    .port_x0_1 (m51_mul_port_y_1[2:0]), //i
    .port_x0_2 (m51_mul_port_y_2[2:0]), //i
    .port_x0_3 (m51_mul_port_y_3[2:0]), //i
    .port_x1_0 (m59_mul_port_y_0[2:0]), //i
    .port_x1_1 (m59_mul_port_y_1[2:0]), //i
    .port_x1_2 (m59_mul_port_y_2[2:0]), //i
    .port_x1_3 (m59_mul_port_y_3[2:0]), //i
    .port_y_0  (l8_xor_port_y_0[2:0] ), //o
    .port_y_1  (l8_xor_port_y_1[2:0] ), //o
    .port_y_2  (l8_xor_port_y_2[2:0] ), //o
    .port_y_3  (l8_xor_port_y_3[2:0] )  //o
  );
  Addition_TI l9_xor (
    .port_x0_0 (m52_mul_port_y_0[2:0]), //i
    .port_x0_1 (m52_mul_port_y_1[2:0]), //i
    .port_x0_2 (m52_mul_port_y_2[2:0]), //i
    .port_x0_3 (m52_mul_port_y_3[2:0]), //i
    .port_x1_0 (m53_mul_port_y_0[2:0]), //i
    .port_x1_1 (m53_mul_port_y_1[2:0]), //i
    .port_x1_2 (m53_mul_port_y_2[2:0]), //i
    .port_x1_3 (m53_mul_port_y_3[2:0]), //i
    .port_y_0  (l9_xor_port_y_0[2:0] ), //o
    .port_y_1  (l9_xor_port_y_1[2:0] ), //o
    .port_y_2  (l9_xor_port_y_2[2:0] ), //o
    .port_y_3  (l9_xor_port_y_3[2:0] )  //o
  );
  Addition_TI l10_xor (
    .port_x0_0 (m53_mul_port_y_0[2:0]), //i
    .port_x0_1 (m53_mul_port_y_1[2:0]), //i
    .port_x0_2 (m53_mul_port_y_2[2:0]), //i
    .port_x0_3 (m53_mul_port_y_3[2:0]), //i
    .port_x1_0 (l4_xor_port_y_0[2:0] ), //i
    .port_x1_1 (l4_xor_port_y_1[2:0] ), //i
    .port_x1_2 (l4_xor_port_y_2[2:0] ), //i
    .port_x1_3 (l4_xor_port_y_3[2:0] ), //i
    .port_y_0  (l10_xor_port_y_0[2:0]), //o
    .port_y_1  (l10_xor_port_y_1[2:0]), //o
    .port_y_2  (l10_xor_port_y_2[2:0]), //o
    .port_y_3  (l10_xor_port_y_3[2:0])  //o
  );
  Addition_TI l11_xor (
    .port_x0_0 (m60_mul_port_y_0[2:0]), //i
    .port_x0_1 (m60_mul_port_y_1[2:0]), //i
    .port_x0_2 (m60_mul_port_y_2[2:0]), //i
    .port_x0_3 (m60_mul_port_y_3[2:0]), //i
    .port_x1_0 (l2_xor_port_y_0[2:0] ), //i
    .port_x1_1 (l2_xor_port_y_1[2:0] ), //i
    .port_x1_2 (l2_xor_port_y_2[2:0] ), //i
    .port_x1_3 (l2_xor_port_y_3[2:0] ), //i
    .port_y_0  (l11_xor_port_y_0[2:0]), //o
    .port_y_1  (l11_xor_port_y_1[2:0]), //o
    .port_y_2  (l11_xor_port_y_2[2:0]), //o
    .port_y_3  (l11_xor_port_y_3[2:0])  //o
  );
  Addition_TI l12_xor (
    .port_x0_0 (m48_mul_port_y_0[2:0]), //i
    .port_x0_1 (m48_mul_port_y_1[2:0]), //i
    .port_x0_2 (m48_mul_port_y_2[2:0]), //i
    .port_x0_3 (m48_mul_port_y_3[2:0]), //i
    .port_x1_0 (m51_mul_port_y_0[2:0]), //i
    .port_x1_1 (m51_mul_port_y_1[2:0]), //i
    .port_x1_2 (m51_mul_port_y_2[2:0]), //i
    .port_x1_3 (m51_mul_port_y_3[2:0]), //i
    .port_y_0  (l12_xor_port_y_0[2:0]), //o
    .port_y_1  (l12_xor_port_y_1[2:0]), //o
    .port_y_2  (l12_xor_port_y_2[2:0]), //o
    .port_y_3  (l12_xor_port_y_3[2:0])  //o
  );
  Addition_TI l13_xor (
    .port_x0_0 (m50_mul_port_y_0[2:0]), //i
    .port_x0_1 (m50_mul_port_y_1[2:0]), //i
    .port_x0_2 (m50_mul_port_y_2[2:0]), //i
    .port_x0_3 (m50_mul_port_y_3[2:0]), //i
    .port_x1_0 (l0_xor_port_y_0[2:0] ), //i
    .port_x1_1 (l0_xor_port_y_1[2:0] ), //i
    .port_x1_2 (l0_xor_port_y_2[2:0] ), //i
    .port_x1_3 (l0_xor_port_y_3[2:0] ), //i
    .port_y_0  (l13_xor_port_y_0[2:0]), //o
    .port_y_1  (l13_xor_port_y_1[2:0]), //o
    .port_y_2  (l13_xor_port_y_2[2:0]), //o
    .port_y_3  (l13_xor_port_y_3[2:0])  //o
  );
  Addition_TI l14_xor (
    .port_x0_0 (m52_mul_port_y_0[2:0]), //i
    .port_x0_1 (m52_mul_port_y_1[2:0]), //i
    .port_x0_2 (m52_mul_port_y_2[2:0]), //i
    .port_x0_3 (m52_mul_port_y_3[2:0]), //i
    .port_x1_0 (m61_mul_port_y_0[2:0]), //i
    .port_x1_1 (m61_mul_port_y_1[2:0]), //i
    .port_x1_2 (m61_mul_port_y_2[2:0]), //i
    .port_x1_3 (m61_mul_port_y_3[2:0]), //i
    .port_y_0  (l14_xor_port_y_0[2:0]), //o
    .port_y_1  (l14_xor_port_y_1[2:0]), //o
    .port_y_2  (l14_xor_port_y_2[2:0]), //o
    .port_y_3  (l14_xor_port_y_3[2:0])  //o
  );
  Addition_TI l15_xor (
    .port_x0_0 (m55_mul_port_y_0[2:0]), //i
    .port_x0_1 (m55_mul_port_y_1[2:0]), //i
    .port_x0_2 (m55_mul_port_y_2[2:0]), //i
    .port_x0_3 (m55_mul_port_y_3[2:0]), //i
    .port_x1_0 (l1_xor_port_y_0[2:0] ), //i
    .port_x1_1 (l1_xor_port_y_1[2:0] ), //i
    .port_x1_2 (l1_xor_port_y_2[2:0] ), //i
    .port_x1_3 (l1_xor_port_y_3[2:0] ), //i
    .port_y_0  (l15_xor_port_y_0[2:0]), //o
    .port_y_1  (l15_xor_port_y_1[2:0]), //o
    .port_y_2  (l15_xor_port_y_2[2:0]), //o
    .port_y_3  (l15_xor_port_y_3[2:0])  //o
  );
  Addition_TI l16_xor (
    .port_x0_0 (m56_mul_port_y_0[2:0]), //i
    .port_x0_1 (m56_mul_port_y_1[2:0]), //i
    .port_x0_2 (m56_mul_port_y_2[2:0]), //i
    .port_x0_3 (m56_mul_port_y_3[2:0]), //i
    .port_x1_0 (l0_xor_port_y_0[2:0] ), //i
    .port_x1_1 (l0_xor_port_y_1[2:0] ), //i
    .port_x1_2 (l0_xor_port_y_2[2:0] ), //i
    .port_x1_3 (l0_xor_port_y_3[2:0] ), //i
    .port_y_0  (l16_xor_port_y_0[2:0]), //o
    .port_y_1  (l16_xor_port_y_1[2:0]), //o
    .port_y_2  (l16_xor_port_y_2[2:0]), //o
    .port_y_3  (l16_xor_port_y_3[2:0])  //o
  );
  Addition_TI l17_xor (
    .port_x0_0 (m57_mul_port_y_0[2:0]), //i
    .port_x0_1 (m57_mul_port_y_1[2:0]), //i
    .port_x0_2 (m57_mul_port_y_2[2:0]), //i
    .port_x0_3 (m57_mul_port_y_3[2:0]), //i
    .port_x1_0 (l1_xor_port_y_0[2:0] ), //i
    .port_x1_1 (l1_xor_port_y_1[2:0] ), //i
    .port_x1_2 (l1_xor_port_y_2[2:0] ), //i
    .port_x1_3 (l1_xor_port_y_3[2:0] ), //i
    .port_y_0  (l17_xor_port_y_0[2:0]), //o
    .port_y_1  (l17_xor_port_y_1[2:0]), //o
    .port_y_2  (l17_xor_port_y_2[2:0]), //o
    .port_y_3  (l17_xor_port_y_3[2:0])  //o
  );
  Addition_TI l18_xor (
    .port_x0_0 (m58_mul_port_y_0[2:0]), //i
    .port_x0_1 (m58_mul_port_y_1[2:0]), //i
    .port_x0_2 (m58_mul_port_y_2[2:0]), //i
    .port_x0_3 (m58_mul_port_y_3[2:0]), //i
    .port_x1_0 (l8_xor_port_y_0[2:0] ), //i
    .port_x1_1 (l8_xor_port_y_1[2:0] ), //i
    .port_x1_2 (l8_xor_port_y_2[2:0] ), //i
    .port_x1_3 (l8_xor_port_y_3[2:0] ), //i
    .port_y_0  (l18_xor_port_y_0[2:0]), //o
    .port_y_1  (l18_xor_port_y_1[2:0]), //o
    .port_y_2  (l18_xor_port_y_2[2:0]), //o
    .port_y_3  (l18_xor_port_y_3[2:0])  //o
  );
  Addition_TI l19_xor (
    .port_x0_0 (m63_mul_port_y_0[2:0]), //i
    .port_x0_1 (m63_mul_port_y_1[2:0]), //i
    .port_x0_2 (m63_mul_port_y_2[2:0]), //i
    .port_x0_3 (m63_mul_port_y_3[2:0]), //i
    .port_x1_0 (l4_xor_port_y_0[2:0] ), //i
    .port_x1_1 (l4_xor_port_y_1[2:0] ), //i
    .port_x1_2 (l4_xor_port_y_2[2:0] ), //i
    .port_x1_3 (l4_xor_port_y_3[2:0] ), //i
    .port_y_0  (l19_xor_port_y_0[2:0]), //o
    .port_y_1  (l19_xor_port_y_1[2:0]), //o
    .port_y_2  (l19_xor_port_y_2[2:0]), //o
    .port_y_3  (l19_xor_port_y_3[2:0])  //o
  );
  Addition_TI l20_xor (
    .port_x0_0 (l0_xor_port_y_0[2:0] ), //i
    .port_x0_1 (l0_xor_port_y_1[2:0] ), //i
    .port_x0_2 (l0_xor_port_y_2[2:0] ), //i
    .port_x0_3 (l0_xor_port_y_3[2:0] ), //i
    .port_x1_0 (l1_xor_port_y_0[2:0] ), //i
    .port_x1_1 (l1_xor_port_y_1[2:0] ), //i
    .port_x1_2 (l1_xor_port_y_2[2:0] ), //i
    .port_x1_3 (l1_xor_port_y_3[2:0] ), //i
    .port_y_0  (l20_xor_port_y_0[2:0]), //o
    .port_y_1  (l20_xor_port_y_1[2:0]), //o
    .port_y_2  (l20_xor_port_y_2[2:0]), //o
    .port_y_3  (l20_xor_port_y_3[2:0])  //o
  );
  Addition_TI l21_xor (
    .port_x0_0 (l1_xor_port_y_0[2:0] ), //i
    .port_x0_1 (l1_xor_port_y_1[2:0] ), //i
    .port_x0_2 (l1_xor_port_y_2[2:0] ), //i
    .port_x0_3 (l1_xor_port_y_3[2:0] ), //i
    .port_x1_0 (l7_xor_port_y_0[2:0] ), //i
    .port_x1_1 (l7_xor_port_y_1[2:0] ), //i
    .port_x1_2 (l7_xor_port_y_2[2:0] ), //i
    .port_x1_3 (l7_xor_port_y_3[2:0] ), //i
    .port_y_0  (l21_xor_port_y_0[2:0]), //o
    .port_y_1  (l21_xor_port_y_1[2:0]), //o
    .port_y_2  (l21_xor_port_y_2[2:0]), //o
    .port_y_3  (l21_xor_port_y_3[2:0])  //o
  );
  Addition_TI l22_xor (
    .port_x0_0 (l3_xor_port_y_0[2:0] ), //i
    .port_x0_1 (l3_xor_port_y_1[2:0] ), //i
    .port_x0_2 (l3_xor_port_y_2[2:0] ), //i
    .port_x0_3 (l3_xor_port_y_3[2:0] ), //i
    .port_x1_0 (l12_xor_port_y_0[2:0]), //i
    .port_x1_1 (l12_xor_port_y_1[2:0]), //i
    .port_x1_2 (l12_xor_port_y_2[2:0]), //i
    .port_x1_3 (l12_xor_port_y_3[2:0]), //i
    .port_y_0  (l22_xor_port_y_0[2:0]), //o
    .port_y_1  (l22_xor_port_y_1[2:0]), //o
    .port_y_2  (l22_xor_port_y_2[2:0]), //o
    .port_y_3  (l22_xor_port_y_3[2:0])  //o
  );
  Addition_TI l23_xor (
    .port_x0_0 (l18_xor_port_y_0[2:0]), //i
    .port_x0_1 (l18_xor_port_y_1[2:0]), //i
    .port_x0_2 (l18_xor_port_y_2[2:0]), //i
    .port_x0_3 (l18_xor_port_y_3[2:0]), //i
    .port_x1_0 (l2_xor_port_y_0[2:0] ), //i
    .port_x1_1 (l2_xor_port_y_1[2:0] ), //i
    .port_x1_2 (l2_xor_port_y_2[2:0] ), //i
    .port_x1_3 (l2_xor_port_y_3[2:0] ), //i
    .port_y_0  (l23_xor_port_y_0[2:0]), //o
    .port_y_1  (l23_xor_port_y_1[2:0]), //o
    .port_y_2  (l23_xor_port_y_2[2:0]), //o
    .port_y_3  (l23_xor_port_y_3[2:0])  //o
  );
  Addition_TI l24_xor (
    .port_x0_0 (l15_xor_port_y_0[2:0]), //i
    .port_x0_1 (l15_xor_port_y_1[2:0]), //i
    .port_x0_2 (l15_xor_port_y_2[2:0]), //i
    .port_x0_3 (l15_xor_port_y_3[2:0]), //i
    .port_x1_0 (l9_xor_port_y_0[2:0] ), //i
    .port_x1_1 (l9_xor_port_y_1[2:0] ), //i
    .port_x1_2 (l9_xor_port_y_2[2:0] ), //i
    .port_x1_3 (l9_xor_port_y_3[2:0] ), //i
    .port_y_0  (l24_xor_port_y_0[2:0]), //o
    .port_y_1  (l24_xor_port_y_1[2:0]), //o
    .port_y_2  (l24_xor_port_y_2[2:0]), //o
    .port_y_3  (l24_xor_port_y_3[2:0])  //o
  );
  Addition_TI l25_xor (
    .port_x0_0 (l6_xor_port_y_0[2:0] ), //i
    .port_x0_1 (l6_xor_port_y_1[2:0] ), //i
    .port_x0_2 (l6_xor_port_y_2[2:0] ), //i
    .port_x0_3 (l6_xor_port_y_3[2:0] ), //i
    .port_x1_0 (l10_xor_port_y_0[2:0]), //i
    .port_x1_1 (l10_xor_port_y_1[2:0]), //i
    .port_x1_2 (l10_xor_port_y_2[2:0]), //i
    .port_x1_3 (l10_xor_port_y_3[2:0]), //i
    .port_y_0  (l25_xor_port_y_0[2:0]), //o
    .port_y_1  (l25_xor_port_y_1[2:0]), //o
    .port_y_2  (l25_xor_port_y_2[2:0]), //o
    .port_y_3  (l25_xor_port_y_3[2:0])  //o
  );
  Addition_TI l26_xor (
    .port_x0_0 (l7_xor_port_y_0[2:0] ), //i
    .port_x0_1 (l7_xor_port_y_1[2:0] ), //i
    .port_x0_2 (l7_xor_port_y_2[2:0] ), //i
    .port_x0_3 (l7_xor_port_y_3[2:0] ), //i
    .port_x1_0 (l9_xor_port_y_0[2:0] ), //i
    .port_x1_1 (l9_xor_port_y_1[2:0] ), //i
    .port_x1_2 (l9_xor_port_y_2[2:0] ), //i
    .port_x1_3 (l9_xor_port_y_3[2:0] ), //i
    .port_y_0  (l26_xor_port_y_0[2:0]), //o
    .port_y_1  (l26_xor_port_y_1[2:0]), //o
    .port_y_2  (l26_xor_port_y_2[2:0]), //o
    .port_y_3  (l26_xor_port_y_3[2:0])  //o
  );
  Addition_TI l27_xor (
    .port_x0_0 (l8_xor_port_y_0[2:0] ), //i
    .port_x0_1 (l8_xor_port_y_1[2:0] ), //i
    .port_x0_2 (l8_xor_port_y_2[2:0] ), //i
    .port_x0_3 (l8_xor_port_y_3[2:0] ), //i
    .port_x1_0 (l10_xor_port_y_0[2:0]), //i
    .port_x1_1 (l10_xor_port_y_1[2:0]), //i
    .port_x1_2 (l10_xor_port_y_2[2:0]), //i
    .port_x1_3 (l10_xor_port_y_3[2:0]), //i
    .port_y_0  (l27_xor_port_y_0[2:0]), //o
    .port_y_1  (l27_xor_port_y_1[2:0]), //o
    .port_y_2  (l27_xor_port_y_2[2:0]), //o
    .port_y_3  (l27_xor_port_y_3[2:0])  //o
  );
  Addition_TI l28_xor (
    .port_x0_0 (l11_xor_port_y_0[2:0]), //i
    .port_x0_1 (l11_xor_port_y_1[2:0]), //i
    .port_x0_2 (l11_xor_port_y_2[2:0]), //i
    .port_x0_3 (l11_xor_port_y_3[2:0]), //i
    .port_x1_0 (l14_xor_port_y_0[2:0]), //i
    .port_x1_1 (l14_xor_port_y_1[2:0]), //i
    .port_x1_2 (l14_xor_port_y_2[2:0]), //i
    .port_x1_3 (l14_xor_port_y_3[2:0]), //i
    .port_y_0  (l28_xor_port_y_0[2:0]), //o
    .port_y_1  (l28_xor_port_y_1[2:0]), //o
    .port_y_2  (l28_xor_port_y_2[2:0]), //o
    .port_y_3  (l28_xor_port_y_3[2:0])  //o
  );
  Addition_TI l29_xor (
    .port_x0_0 (l11_xor_port_y_0[2:0]), //i
    .port_x0_1 (l11_xor_port_y_1[2:0]), //i
    .port_x0_2 (l11_xor_port_y_2[2:0]), //i
    .port_x0_3 (l11_xor_port_y_3[2:0]), //i
    .port_x1_0 (l17_xor_port_y_0[2:0]), //i
    .port_x1_1 (l17_xor_port_y_1[2:0]), //i
    .port_x1_2 (l17_xor_port_y_2[2:0]), //i
    .port_x1_3 (l17_xor_port_y_3[2:0]), //i
    .port_y_0  (l29_xor_port_y_0[2:0]), //o
    .port_y_1  (l29_xor_port_y_1[2:0]), //o
    .port_y_2  (l29_xor_port_y_2[2:0]), //o
    .port_y_3  (l29_xor_port_y_3[2:0])  //o
  );
  Addition_TI s0 (
    .port_x0_0 (l6_xor_port_y_0[2:0] ), //i
    .port_x0_1 (l6_xor_port_y_1[2:0] ), //i
    .port_x0_2 (l6_xor_port_y_2[2:0] ), //i
    .port_x0_3 (l6_xor_port_y_3[2:0] ), //i
    .port_x1_0 (l24_xor_port_y_0[2:0]), //i
    .port_x1_1 (l24_xor_port_y_1[2:0]), //i
    .port_x1_2 (l24_xor_port_y_2[2:0]), //i
    .port_x1_3 (l24_xor_port_y_3[2:0]), //i
    .port_y_0  (s0_port_y_0[2:0]     ), //o
    .port_y_1  (s0_port_y_1[2:0]     ), //o
    .port_y_2  (s0_port_y_2[2:0]     ), //o
    .port_y_3  (s0_port_y_3[2:0]     )  //o
  );
  Addition_Inv_TI s1 (
    .port_x0_0 (l16_xor_port_y_0[2:0]), //i
    .port_x0_1 (l16_xor_port_y_1[2:0]), //i
    .port_x0_2 (l16_xor_port_y_2[2:0]), //i
    .port_x0_3 (l16_xor_port_y_3[2:0]), //i
    .port_x1_0 (l26_xor_port_y_0[2:0]), //i
    .port_x1_1 (l26_xor_port_y_1[2:0]), //i
    .port_x1_2 (l26_xor_port_y_2[2:0]), //i
    .port_x1_3 (l26_xor_port_y_3[2:0]), //i
    .port_y_0  (s1_port_y_0[2:0]     ), //o
    .port_y_1  (s1_port_y_1[2:0]     ), //o
    .port_y_2  (s1_port_y_2[2:0]     ), //o
    .port_y_3  (s1_port_y_3[2:0]     )  //o
  );
  Addition_Inv_TI s2 (
    .port_x0_0 (l19_xor_port_y_0[2:0]), //i
    .port_x0_1 (l19_xor_port_y_1[2:0]), //i
    .port_x0_2 (l19_xor_port_y_2[2:0]), //i
    .port_x0_3 (l19_xor_port_y_3[2:0]), //i
    .port_x1_0 (l28_xor_port_y_0[2:0]), //i
    .port_x1_1 (l28_xor_port_y_1[2:0]), //i
    .port_x1_2 (l28_xor_port_y_2[2:0]), //i
    .port_x1_3 (l28_xor_port_y_3[2:0]), //i
    .port_y_0  (s2_port_y_0[2:0]     ), //o
    .port_y_1  (s2_port_y_1[2:0]     ), //o
    .port_y_2  (s2_port_y_2[2:0]     ), //o
    .port_y_3  (s2_port_y_3[2:0]     )  //o
  );
  Addition_TI s3 (
    .port_x0_0 (l6_xor_port_y_0[2:0] ), //i
    .port_x0_1 (l6_xor_port_y_1[2:0] ), //i
    .port_x0_2 (l6_xor_port_y_2[2:0] ), //i
    .port_x0_3 (l6_xor_port_y_3[2:0] ), //i
    .port_x1_0 (l21_xor_port_y_0[2:0]), //i
    .port_x1_1 (l21_xor_port_y_1[2:0]), //i
    .port_x1_2 (l21_xor_port_y_2[2:0]), //i
    .port_x1_3 (l21_xor_port_y_3[2:0]), //i
    .port_y_0  (s3_port_y_0[2:0]     ), //o
    .port_y_1  (s3_port_y_1[2:0]     ), //o
    .port_y_2  (s3_port_y_2[2:0]     ), //o
    .port_y_3  (s3_port_y_3[2:0]     )  //o
  );
  Addition_TI s4 (
    .port_x0_0 (l20_xor_port_y_0[2:0]), //i
    .port_x0_1 (l20_xor_port_y_1[2:0]), //i
    .port_x0_2 (l20_xor_port_y_2[2:0]), //i
    .port_x0_3 (l20_xor_port_y_3[2:0]), //i
    .port_x1_0 (l22_xor_port_y_0[2:0]), //i
    .port_x1_1 (l22_xor_port_y_1[2:0]), //i
    .port_x1_2 (l22_xor_port_y_2[2:0]), //i
    .port_x1_3 (l22_xor_port_y_3[2:0]), //i
    .port_y_0  (s4_port_y_0[2:0]     ), //o
    .port_y_1  (s4_port_y_1[2:0]     ), //o
    .port_y_2  (s4_port_y_2[2:0]     ), //o
    .port_y_3  (s4_port_y_3[2:0]     )  //o
  );
  Addition_TI s5 (
    .port_x0_0 (l25_xor_port_y_0[2:0]), //i
    .port_x0_1 (l25_xor_port_y_1[2:0]), //i
    .port_x0_2 (l25_xor_port_y_2[2:0]), //i
    .port_x0_3 (l25_xor_port_y_3[2:0]), //i
    .port_x1_0 (l29_xor_port_y_0[2:0]), //i
    .port_x1_1 (l29_xor_port_y_1[2:0]), //i
    .port_x1_2 (l29_xor_port_y_2[2:0]), //i
    .port_x1_3 (l29_xor_port_y_3[2:0]), //i
    .port_y_0  (s5_port_y_0[2:0]     ), //o
    .port_y_1  (s5_port_y_1[2:0]     ), //o
    .port_y_2  (s5_port_y_2[2:0]     ), //o
    .port_y_3  (s5_port_y_3[2:0]     )  //o
  );
  Addition_Inv_TI s6 (
    .port_x0_0 (l13_xor_port_y_0[2:0]), //i
    .port_x0_1 (l13_xor_port_y_1[2:0]), //i
    .port_x0_2 (l13_xor_port_y_2[2:0]), //i
    .port_x0_3 (l13_xor_port_y_3[2:0]), //i
    .port_x1_0 (l27_xor_port_y_0[2:0]), //i
    .port_x1_1 (l27_xor_port_y_1[2:0]), //i
    .port_x1_2 (l27_xor_port_y_2[2:0]), //i
    .port_x1_3 (l27_xor_port_y_3[2:0]), //i
    .port_y_0  (s6_port_y_0[2:0]     ), //o
    .port_y_1  (s6_port_y_1[2:0]     ), //o
    .port_y_2  (s6_port_y_2[2:0]     ), //o
    .port_y_3  (s6_port_y_3[2:0]     )  //o
  );
  Addition_Inv_TI s7 (
    .port_x0_0 (l6_xor_port_y_0[2:0] ), //i
    .port_x0_1 (l6_xor_port_y_1[2:0] ), //i
    .port_x0_2 (l6_xor_port_y_2[2:0] ), //i
    .port_x0_3 (l6_xor_port_y_3[2:0] ), //i
    .port_x1_0 (l23_xor_port_y_0[2:0]), //i
    .port_x1_1 (l23_xor_port_y_1[2:0]), //i
    .port_x1_2 (l23_xor_port_y_2[2:0]), //i
    .port_x1_3 (l23_xor_port_y_3[2:0]), //i
    .port_y_0  (s7_port_y_0[2:0]     ), //o
    .port_y_1  (s7_port_y_1[2:0]     ), //o
    .port_y_2  (s7_port_y_2[2:0]     ), //o
    .port_y_3  (s7_port_y_3[2:0]     )  //o
  );
  assign in_x0_0 = port_i_0_7;
  assign in_x1_0 = port_i_0_6;
  assign in_x2_0 = port_i_0_5;
  assign in_x3_0 = port_i_0_4;
  assign in_x4_0 = port_i_0_3;
  assign in_x5_0 = port_i_0_2;
  assign in_x6_0 = port_i_0_1;
  assign in_x7_0 = port_i_0_0;
  assign in_x0_1 = port_i_1_7;
  assign in_x1_1 = port_i_1_6;
  assign in_x2_1 = port_i_1_5;
  assign in_x3_1 = port_i_1_4;
  assign in_x4_1 = port_i_1_3;
  assign in_x5_1 = port_i_1_2;
  assign in_x6_1 = port_i_1_1;
  assign in_x7_1 = port_i_1_0;
  assign in_x0_2 = port_i_2_7;
  assign in_x1_2 = port_i_2_6;
  assign in_x2_2 = port_i_2_5;
  assign in_x3_2 = port_i_2_4;
  assign in_x4_2 = port_i_2_3;
  assign in_x5_2 = port_i_2_2;
  assign in_x6_2 = port_i_2_1;
  assign in_x7_2 = port_i_2_0;
  assign in_x0_3 = port_i_3_7;
  assign in_x1_3 = port_i_3_6;
  assign in_x2_3 = port_i_3_5;
  assign in_x3_3 = port_i_3_4;
  assign in_x4_3 = port_i_3_3;
  assign in_x5_3 = port_i_3_2;
  assign in_x6_3 = port_i_3_1;
  assign in_x7_3 = port_i_3_0;
  assign out_y0_0 = s0_port_y_0;
  assign out_y0_1 = s0_port_y_1;
  assign out_y0_2 = s0_port_y_2;
  assign out_y0_3 = s0_port_y_3;
  assign out_y1_0 = s1_port_y_0;
  assign out_y1_1 = s1_port_y_1;
  assign out_y1_2 = s1_port_y_2;
  assign out_y1_3 = s1_port_y_3;
  assign out_y2_0 = s2_port_y_0;
  assign out_y2_1 = s2_port_y_1;
  assign out_y2_2 = s2_port_y_2;
  assign out_y2_3 = s2_port_y_3;
  assign out_y3_0 = s3_port_y_0;
  assign out_y3_1 = s3_port_y_1;
  assign out_y3_2 = s3_port_y_2;
  assign out_y3_3 = s3_port_y_3;
  assign out_y4_0 = s4_port_y_0;
  assign out_y4_1 = s4_port_y_1;
  assign out_y4_2 = s4_port_y_2;
  assign out_y4_3 = s4_port_y_3;
  assign out_y5_0 = s5_port_y_0;
  assign out_y5_1 = s5_port_y_1;
  assign out_y5_2 = s5_port_y_2;
  assign out_y5_3 = s5_port_y_3;
  assign out_y6_0 = s6_port_y_0;
  assign out_y6_1 = s6_port_y_1;
  assign out_y6_2 = s6_port_y_2;
  assign out_y6_3 = s6_port_y_3;
  assign out_y7_0 = s7_port_y_0;
  assign out_y7_1 = s7_port_y_1;
  assign out_y7_2 = s7_port_y_2;
  assign out_y7_3 = s7_port_y_3;
  assign port_o_0_7 = out_y0_0;
  assign port_o_0_6 = out_y1_0;
  assign port_o_0_5 = out_y2_0;
  assign port_o_0_4 = out_y3_0;
  assign port_o_0_3 = out_y4_0;
  assign port_o_0_2 = out_y5_0;
  assign port_o_0_1 = out_y6_0;
  assign port_o_0_0 = out_y7_0;
  assign port_o_1_7 = out_y0_1;
  assign port_o_1_6 = out_y1_1;
  assign port_o_1_5 = out_y2_1;
  assign port_o_1_4 = out_y3_1;
  assign port_o_1_3 = out_y4_1;
  assign port_o_1_2 = out_y5_1;
  assign port_o_1_1 = out_y6_1;
  assign port_o_1_0 = out_y7_1;
  assign port_o_2_7 = out_y0_2;
  assign port_o_2_6 = out_y1_2;
  assign port_o_2_5 = out_y2_2;
  assign port_o_2_4 = out_y3_2;
  assign port_o_2_3 = out_y4_2;
  assign port_o_2_2 = out_y5_2;
  assign port_o_2_1 = out_y6_2;
  assign port_o_2_0 = out_y7_2;
  assign port_o_3_7 = out_y0_3;
  assign port_o_3_6 = out_y1_3;
  assign port_o_3_5 = out_y2_3;
  assign port_o_3_4 = out_y3_3;
  assign port_o_3_3 = out_y4_3;
  assign port_o_3_2 = out_y5_3;
  assign port_o_3_1 = out_y6_3;
  assign port_o_3_0 = out_y7_3;
  always @(posedge clk) begin
    x7_0 <= in_x7_0;
    x7_1 <= in_x7_1;
    x7_2 <= in_x7_2;
    x7_3 <= in_x7_3;
    t1_0 <= t1_xor_port_y_0;
    t1_1 <= t1_xor_port_y_1;
    t1_2 <= t1_xor_port_y_2;
    t1_3 <= t1_xor_port_y_3;
    t2_0 <= t2_xor_port_y_0;
    t2_1 <= t2_xor_port_y_1;
    t2_2 <= t2_xor_port_y_2;
    t2_3 <= t2_xor_port_y_3;
    t3_0 <= t3_xor_port_y_0;
    t3_1 <= t3_xor_port_y_1;
    t3_2 <= t3_xor_port_y_2;
    t3_3 <= t3_xor_port_y_3;
    t4_0 <= t4_xor_port_y_0;
    t4_1 <= t4_xor_port_y_1;
    t4_2 <= t4_xor_port_y_2;
    t4_3 <= t4_xor_port_y_3;
    t6_0 <= t6_xor_port_y_0;
    t6_1 <= t6_xor_port_y_1;
    t6_2 <= t6_xor_port_y_2;
    t6_3 <= t6_xor_port_y_3;
    t7_0 <= t7_xor_port_y_0;
    t7_1 <= t7_xor_port_y_1;
    t7_2 <= t7_xor_port_y_2;
    t7_3 <= t7_xor_port_y_3;
    t8_0 <= t8_xor_port_y_0;
    t8_1 <= t8_xor_port_y_1;
    t8_2 <= t8_xor_port_y_2;
    t8_3 <= t8_xor_port_y_3;
    t9_0 <= t9_xor_port_y_0;
    t9_1 <= t9_xor_port_y_1;
    t9_2 <= t9_xor_port_y_2;
    t9_3 <= t9_xor_port_y_3;
    t10_0 <= t10_xor_port_y_0;
    t10_1 <= t10_xor_port_y_1;
    t10_2 <= t10_xor_port_y_2;
    t10_3 <= t10_xor_port_y_3;
    t13_0 <= t13_xor_port_y_0;
    t13_1 <= t13_xor_port_y_1;
    t13_2 <= t13_xor_port_y_2;
    t13_3 <= t13_xor_port_y_3;
    t14_0 <= t14_xor_port_y_0;
    t14_1 <= t14_xor_port_y_1;
    t14_2 <= t14_xor_port_y_2;
    t14_3 <= t14_xor_port_y_3;
    t15_0 <= t15_xor_port_y_0;
    t15_1 <= t15_xor_port_y_1;
    t15_2 <= t15_xor_port_y_2;
    t15_3 <= t15_xor_port_y_3;
    t16_0 <= t16_xor_port_y_0;
    t16_1 <= t16_xor_port_y_1;
    t16_2 <= t16_xor_port_y_2;
    t16_3 <= t16_xor_port_y_3;
    t17_0 <= t17_xor_port_y_0;
    t17_1 <= t17_xor_port_y_1;
    t17_2 <= t17_xor_port_y_2;
    t17_3 <= t17_xor_port_y_3;
    t19_0 <= t19_xor_port_y_0;
    t19_1 <= t19_xor_port_y_1;
    t19_2 <= t19_xor_port_y_2;
    t19_3 <= t19_xor_port_y_3;
    t20_0 <= t20_xor_port_y_0;
    t20_1 <= t20_xor_port_y_1;
    t20_2 <= t20_xor_port_y_2;
    t20_3 <= t20_xor_port_y_3;
    t22_0 <= t22_xor_port_y_0;
    t22_1 <= t22_xor_port_y_1;
    t22_2 <= t22_xor_port_y_2;
    t22_3 <= t22_xor_port_y_3;
    t23_0 <= t23_xor_port_y_0;
    t23_1 <= t23_xor_port_y_1;
    t23_2 <= t23_xor_port_y_2;
    t23_3 <= t23_xor_port_y_3;
    t24_0 <= t24_xor_port_y_0;
    t24_1 <= t24_xor_port_y_1;
    t24_2 <= t24_xor_port_y_2;
    t24_3 <= t24_xor_port_y_3;
    t25_0 <= t25_xor_port_y_0;
    t25_1 <= t25_xor_port_y_1;
    t25_2 <= t25_xor_port_y_2;
    t25_3 <= t25_xor_port_y_3;
    t26_0 <= t26_xor_port_y_0;
    t26_1 <= t26_xor_port_y_1;
    t26_2 <= t26_xor_port_y_2;
    t26_3 <= t26_xor_port_y_3;
    t27_0 <= t27_xor_port_y_0;
    t27_1 <= t27_xor_port_y_1;
    t27_2 <= t27_xor_port_y_2;
    t27_3 <= t27_xor_port_y_3;
    x7_1_0 <= x7_0;
    x7_1_1 <= x7_1;
    x7_1_2 <= x7_2;
    x7_1_3 <= x7_3;
    t1_1_0 <= t1_0;
    t1_1_1 <= t1_1;
    t1_1_2 <= t1_2;
    t1_1_3 <= t1_3;
    t2_1_0 <= t2_0;
    t2_1_1 <= t2_1;
    t2_1_2 <= t2_2;
    t2_1_3 <= t2_3;
    t3_1_0 <= t3_0;
    t3_1_1 <= t3_1;
    t3_1_2 <= t3_2;
    t3_1_3 <= t3_3;
    t4_1_0 <= t4_0;
    t4_1_1 <= t4_1;
    t4_1_2 <= t4_2;
    t4_1_3 <= t4_3;
    t6_1_0 <= t6_0;
    t6_1_1 <= t6_1;
    t6_1_2 <= t6_2;
    t6_1_3 <= t6_3;
    t8_1_0 <= t8_0;
    t8_1_1 <= t8_1;
    t8_1_2 <= t8_2;
    t8_1_3 <= t8_3;
    t9_1_0 <= t9_0;
    t9_1_1 <= t9_1;
    t9_1_2 <= t9_2;
    t9_1_3 <= t9_3;
    t10_1_0 <= t10_0;
    t10_1_1 <= t10_1;
    t10_1_2 <= t10_2;
    t10_1_3 <= t10_3;
    t13_1_0 <= t13_0;
    t13_1_1 <= t13_1;
    t13_1_2 <= t13_2;
    t13_1_3 <= t13_3;
    t15_1_0 <= t15_0;
    t15_1_1 <= t15_1;
    t15_1_2 <= t15_2;
    t15_1_3 <= t15_3;
    t16_1_0 <= t16_0;
    t16_1_1 <= t16_1;
    t16_1_2 <= t16_2;
    t16_1_3 <= t16_3;
    t17_1_0 <= t17_0;
    t17_1_1 <= t17_1;
    t17_1_2 <= t17_2;
    t17_1_3 <= t17_3;
    t19_1_0 <= t19_0;
    t19_1_1 <= t19_1;
    t19_1_2 <= t19_2;
    t19_1_3 <= t19_3;
    t20_1_0 <= t20_0;
    t20_1_1 <= t20_1;
    t20_1_2 <= t20_2;
    t20_1_3 <= t20_3;
    t22_1_0 <= t22_0;
    t22_1_1 <= t22_1;
    t22_1_2 <= t22_2;
    t22_1_3 <= t22_3;
    t23_1_0 <= t23_0;
    t23_1_1 <= t23_1;
    t23_1_2 <= t23_2;
    t23_1_3 <= t23_3;
    t27_1_0 <= t27_0;
    t27_1_1 <= t27_1;
    t27_1_2 <= t27_2;
    t27_1_3 <= t27_3;
    m21_0 <= m21_xor_port_y_0;
    m21_1 <= m21_xor_port_y_1;
    m21_2 <= m21_xor_port_y_2;
    m21_3 <= m21_xor_port_y_3;
    m23_0 <= m23_xor_port_y_0;
    m23_1 <= m23_xor_port_y_1;
    m23_2 <= m23_xor_port_y_2;
    m23_3 <= m23_xor_port_y_3;
    m24_0 <= m24_xor_port_y_0;
    m24_1 <= m24_xor_port_y_1;
    m24_2 <= m24_xor_port_y_2;
    m24_3 <= m24_xor_port_y_3;
    m27_0 <= m27_xor_port_y_0;
    m27_1 <= m27_xor_port_y_1;
    m27_2 <= m27_xor_port_y_2;
    m27_3 <= m27_xor_port_y_3;
    x7_2_0 <= x7_1_0;
    x7_2_1 <= x7_1_1;
    x7_2_2 <= x7_1_2;
    x7_2_3 <= x7_1_3;
    t1_2_0 <= t1_1_0;
    t1_2_1 <= t1_1_1;
    t1_2_2 <= t1_1_2;
    t1_2_3 <= t1_1_3;
    t2_2_0 <= t2_1_0;
    t2_2_1 <= t2_1_1;
    t2_2_2 <= t2_1_2;
    t2_2_3 <= t2_1_3;
    t3_2_0 <= t3_1_0;
    t3_2_1 <= t3_1_1;
    t3_2_2 <= t3_1_2;
    t3_2_3 <= t3_1_3;
    t4_2_0 <= t4_1_0;
    t4_2_1 <= t4_1_1;
    t4_2_2 <= t4_1_2;
    t4_2_3 <= t4_1_3;
    t6_2_0 <= t6_1_0;
    t6_2_1 <= t6_1_1;
    t6_2_2 <= t6_1_2;
    t6_2_3 <= t6_1_3;
    t8_2_0 <= t8_1_0;
    t8_2_1 <= t8_1_1;
    t8_2_2 <= t8_1_2;
    t8_2_3 <= t8_1_3;
    t9_2_0 <= t9_1_0;
    t9_2_1 <= t9_1_1;
    t9_2_2 <= t9_1_2;
    t9_2_3 <= t9_1_3;
    t10_2_0 <= t10_1_0;
    t10_2_1 <= t10_1_1;
    t10_2_2 <= t10_1_2;
    t10_2_3 <= t10_1_3;
    t13_2_0 <= t13_1_0;
    t13_2_1 <= t13_1_1;
    t13_2_2 <= t13_1_2;
    t13_2_3 <= t13_1_3;
    t15_2_0 <= t15_1_0;
    t15_2_1 <= t15_1_1;
    t15_2_2 <= t15_1_2;
    t15_2_3 <= t15_1_3;
    t16_2_0 <= t16_1_0;
    t16_2_1 <= t16_1_1;
    t16_2_2 <= t16_1_2;
    t16_2_3 <= t16_1_3;
    t17_2_0 <= t17_1_0;
    t17_2_1 <= t17_1_1;
    t17_2_2 <= t17_1_2;
    t17_2_3 <= t17_1_3;
    t19_2_0 <= t19_1_0;
    t19_2_1 <= t19_1_1;
    t19_2_2 <= t19_1_2;
    t19_2_3 <= t19_1_3;
    t20_2_0 <= t20_1_0;
    t20_2_1 <= t20_1_1;
    t20_2_2 <= t20_1_2;
    t20_2_3 <= t20_1_3;
    t22_2_0 <= t22_1_0;
    t22_2_1 <= t22_1_1;
    t22_2_2 <= t22_1_2;
    t22_2_3 <= t22_1_3;
    t23_2_0 <= t23_1_0;
    t23_2_1 <= t23_1_1;
    t23_2_2 <= t23_1_2;
    t23_2_3 <= t23_1_3;
    t27_2_0 <= t27_1_0;
    t27_2_1 <= t27_1_1;
    t27_2_2 <= t27_1_2;
    t27_2_3 <= t27_1_3;
    m21_1_0 <= m21_0;
    m21_1_1 <= m21_1;
    m21_1_2 <= m21_2;
    m21_1_3 <= m21_3;
    m23_1_0 <= m23_0;
    m23_1_1 <= m23_1;
    m23_1_2 <= m23_2;
    m23_1_3 <= m23_3;
    m33_0 <= m33_xor_port_y_0;
    m33_1 <= m33_xor_port_y_1;
    m33_2 <= m33_xor_port_y_2;
    m33_3 <= m33_xor_port_y_3;
    m36_0 <= m36_xor_port_y_0;
    m36_1 <= m36_xor_port_y_1;
    m36_2 <= m36_xor_port_y_2;
    m36_3 <= m36_xor_port_y_3;
  end


endmodule

module AES_KeyAddition (
  input      [2:0]    port_state_in_0_0_0,
  input      [2:0]    port_state_in_0_0_1,
  input      [2:0]    port_state_in_0_0_2,
  input      [2:0]    port_state_in_0_0_3,
  input      [2:0]    port_state_in_0_0_4,
  input      [2:0]    port_state_in_0_0_5,
  input      [2:0]    port_state_in_0_0_6,
  input      [2:0]    port_state_in_0_0_7,
  input      [2:0]    port_state_in_0_1_0,
  input      [2:0]    port_state_in_0_1_1,
  input      [2:0]    port_state_in_0_1_2,
  input      [2:0]    port_state_in_0_1_3,
  input      [2:0]    port_state_in_0_1_4,
  input      [2:0]    port_state_in_0_1_5,
  input      [2:0]    port_state_in_0_1_6,
  input      [2:0]    port_state_in_0_1_7,
  input      [2:0]    port_state_in_0_2_0,
  input      [2:0]    port_state_in_0_2_1,
  input      [2:0]    port_state_in_0_2_2,
  input      [2:0]    port_state_in_0_2_3,
  input      [2:0]    port_state_in_0_2_4,
  input      [2:0]    port_state_in_0_2_5,
  input      [2:0]    port_state_in_0_2_6,
  input      [2:0]    port_state_in_0_2_7,
  input      [2:0]    port_state_in_0_3_0,
  input      [2:0]    port_state_in_0_3_1,
  input      [2:0]    port_state_in_0_3_2,
  input      [2:0]    port_state_in_0_3_3,
  input      [2:0]    port_state_in_0_3_4,
  input      [2:0]    port_state_in_0_3_5,
  input      [2:0]    port_state_in_0_3_6,
  input      [2:0]    port_state_in_0_3_7,
  input      [2:0]    port_state_in_1_0_0,
  input      [2:0]    port_state_in_1_0_1,
  input      [2:0]    port_state_in_1_0_2,
  input      [2:0]    port_state_in_1_0_3,
  input      [2:0]    port_state_in_1_0_4,
  input      [2:0]    port_state_in_1_0_5,
  input      [2:0]    port_state_in_1_0_6,
  input      [2:0]    port_state_in_1_0_7,
  input      [2:0]    port_state_in_1_1_0,
  input      [2:0]    port_state_in_1_1_1,
  input      [2:0]    port_state_in_1_1_2,
  input      [2:0]    port_state_in_1_1_3,
  input      [2:0]    port_state_in_1_1_4,
  input      [2:0]    port_state_in_1_1_5,
  input      [2:0]    port_state_in_1_1_6,
  input      [2:0]    port_state_in_1_1_7,
  input      [2:0]    port_state_in_1_2_0,
  input      [2:0]    port_state_in_1_2_1,
  input      [2:0]    port_state_in_1_2_2,
  input      [2:0]    port_state_in_1_2_3,
  input      [2:0]    port_state_in_1_2_4,
  input      [2:0]    port_state_in_1_2_5,
  input      [2:0]    port_state_in_1_2_6,
  input      [2:0]    port_state_in_1_2_7,
  input      [2:0]    port_state_in_1_3_0,
  input      [2:0]    port_state_in_1_3_1,
  input      [2:0]    port_state_in_1_3_2,
  input      [2:0]    port_state_in_1_3_3,
  input      [2:0]    port_state_in_1_3_4,
  input      [2:0]    port_state_in_1_3_5,
  input      [2:0]    port_state_in_1_3_6,
  input      [2:0]    port_state_in_1_3_7,
  input      [2:0]    port_state_in_2_0_0,
  input      [2:0]    port_state_in_2_0_1,
  input      [2:0]    port_state_in_2_0_2,
  input      [2:0]    port_state_in_2_0_3,
  input      [2:0]    port_state_in_2_0_4,
  input      [2:0]    port_state_in_2_0_5,
  input      [2:0]    port_state_in_2_0_6,
  input      [2:0]    port_state_in_2_0_7,
  input      [2:0]    port_state_in_2_1_0,
  input      [2:0]    port_state_in_2_1_1,
  input      [2:0]    port_state_in_2_1_2,
  input      [2:0]    port_state_in_2_1_3,
  input      [2:0]    port_state_in_2_1_4,
  input      [2:0]    port_state_in_2_1_5,
  input      [2:0]    port_state_in_2_1_6,
  input      [2:0]    port_state_in_2_1_7,
  input      [2:0]    port_state_in_2_2_0,
  input      [2:0]    port_state_in_2_2_1,
  input      [2:0]    port_state_in_2_2_2,
  input      [2:0]    port_state_in_2_2_3,
  input      [2:0]    port_state_in_2_2_4,
  input      [2:0]    port_state_in_2_2_5,
  input      [2:0]    port_state_in_2_2_6,
  input      [2:0]    port_state_in_2_2_7,
  input      [2:0]    port_state_in_2_3_0,
  input      [2:0]    port_state_in_2_3_1,
  input      [2:0]    port_state_in_2_3_2,
  input      [2:0]    port_state_in_2_3_3,
  input      [2:0]    port_state_in_2_3_4,
  input      [2:0]    port_state_in_2_3_5,
  input      [2:0]    port_state_in_2_3_6,
  input      [2:0]    port_state_in_2_3_7,
  input      [2:0]    port_state_in_3_0_0,
  input      [2:0]    port_state_in_3_0_1,
  input      [2:0]    port_state_in_3_0_2,
  input      [2:0]    port_state_in_3_0_3,
  input      [2:0]    port_state_in_3_0_4,
  input      [2:0]    port_state_in_3_0_5,
  input      [2:0]    port_state_in_3_0_6,
  input      [2:0]    port_state_in_3_0_7,
  input      [2:0]    port_state_in_3_1_0,
  input      [2:0]    port_state_in_3_1_1,
  input      [2:0]    port_state_in_3_1_2,
  input      [2:0]    port_state_in_3_1_3,
  input      [2:0]    port_state_in_3_1_4,
  input      [2:0]    port_state_in_3_1_5,
  input      [2:0]    port_state_in_3_1_6,
  input      [2:0]    port_state_in_3_1_7,
  input      [2:0]    port_state_in_3_2_0,
  input      [2:0]    port_state_in_3_2_1,
  input      [2:0]    port_state_in_3_2_2,
  input      [2:0]    port_state_in_3_2_3,
  input      [2:0]    port_state_in_3_2_4,
  input      [2:0]    port_state_in_3_2_5,
  input      [2:0]    port_state_in_3_2_6,
  input      [2:0]    port_state_in_3_2_7,
  input      [2:0]    port_state_in_3_3_0,
  input      [2:0]    port_state_in_3_3_1,
  input      [2:0]    port_state_in_3_3_2,
  input      [2:0]    port_state_in_3_3_3,
  input      [2:0]    port_state_in_3_3_4,
  input      [2:0]    port_state_in_3_3_5,
  input      [2:0]    port_state_in_3_3_6,
  input      [2:0]    port_state_in_3_3_7,
  input      [2:0]    port_state_in_4_0_0,
  input      [2:0]    port_state_in_4_0_1,
  input      [2:0]    port_state_in_4_0_2,
  input      [2:0]    port_state_in_4_0_3,
  input      [2:0]    port_state_in_4_0_4,
  input      [2:0]    port_state_in_4_0_5,
  input      [2:0]    port_state_in_4_0_6,
  input      [2:0]    port_state_in_4_0_7,
  input      [2:0]    port_state_in_4_1_0,
  input      [2:0]    port_state_in_4_1_1,
  input      [2:0]    port_state_in_4_1_2,
  input      [2:0]    port_state_in_4_1_3,
  input      [2:0]    port_state_in_4_1_4,
  input      [2:0]    port_state_in_4_1_5,
  input      [2:0]    port_state_in_4_1_6,
  input      [2:0]    port_state_in_4_1_7,
  input      [2:0]    port_state_in_4_2_0,
  input      [2:0]    port_state_in_4_2_1,
  input      [2:0]    port_state_in_4_2_2,
  input      [2:0]    port_state_in_4_2_3,
  input      [2:0]    port_state_in_4_2_4,
  input      [2:0]    port_state_in_4_2_5,
  input      [2:0]    port_state_in_4_2_6,
  input      [2:0]    port_state_in_4_2_7,
  input      [2:0]    port_state_in_4_3_0,
  input      [2:0]    port_state_in_4_3_1,
  input      [2:0]    port_state_in_4_3_2,
  input      [2:0]    port_state_in_4_3_3,
  input      [2:0]    port_state_in_4_3_4,
  input      [2:0]    port_state_in_4_3_5,
  input      [2:0]    port_state_in_4_3_6,
  input      [2:0]    port_state_in_4_3_7,
  input      [2:0]    port_state_in_5_0_0,
  input      [2:0]    port_state_in_5_0_1,
  input      [2:0]    port_state_in_5_0_2,
  input      [2:0]    port_state_in_5_0_3,
  input      [2:0]    port_state_in_5_0_4,
  input      [2:0]    port_state_in_5_0_5,
  input      [2:0]    port_state_in_5_0_6,
  input      [2:0]    port_state_in_5_0_7,
  input      [2:0]    port_state_in_5_1_0,
  input      [2:0]    port_state_in_5_1_1,
  input      [2:0]    port_state_in_5_1_2,
  input      [2:0]    port_state_in_5_1_3,
  input      [2:0]    port_state_in_5_1_4,
  input      [2:0]    port_state_in_5_1_5,
  input      [2:0]    port_state_in_5_1_6,
  input      [2:0]    port_state_in_5_1_7,
  input      [2:0]    port_state_in_5_2_0,
  input      [2:0]    port_state_in_5_2_1,
  input      [2:0]    port_state_in_5_2_2,
  input      [2:0]    port_state_in_5_2_3,
  input      [2:0]    port_state_in_5_2_4,
  input      [2:0]    port_state_in_5_2_5,
  input      [2:0]    port_state_in_5_2_6,
  input      [2:0]    port_state_in_5_2_7,
  input      [2:0]    port_state_in_5_3_0,
  input      [2:0]    port_state_in_5_3_1,
  input      [2:0]    port_state_in_5_3_2,
  input      [2:0]    port_state_in_5_3_3,
  input      [2:0]    port_state_in_5_3_4,
  input      [2:0]    port_state_in_5_3_5,
  input      [2:0]    port_state_in_5_3_6,
  input      [2:0]    port_state_in_5_3_7,
  input      [2:0]    port_state_in_6_0_0,
  input      [2:0]    port_state_in_6_0_1,
  input      [2:0]    port_state_in_6_0_2,
  input      [2:0]    port_state_in_6_0_3,
  input      [2:0]    port_state_in_6_0_4,
  input      [2:0]    port_state_in_6_0_5,
  input      [2:0]    port_state_in_6_0_6,
  input      [2:0]    port_state_in_6_0_7,
  input      [2:0]    port_state_in_6_1_0,
  input      [2:0]    port_state_in_6_1_1,
  input      [2:0]    port_state_in_6_1_2,
  input      [2:0]    port_state_in_6_1_3,
  input      [2:0]    port_state_in_6_1_4,
  input      [2:0]    port_state_in_6_1_5,
  input      [2:0]    port_state_in_6_1_6,
  input      [2:0]    port_state_in_6_1_7,
  input      [2:0]    port_state_in_6_2_0,
  input      [2:0]    port_state_in_6_2_1,
  input      [2:0]    port_state_in_6_2_2,
  input      [2:0]    port_state_in_6_2_3,
  input      [2:0]    port_state_in_6_2_4,
  input      [2:0]    port_state_in_6_2_5,
  input      [2:0]    port_state_in_6_2_6,
  input      [2:0]    port_state_in_6_2_7,
  input      [2:0]    port_state_in_6_3_0,
  input      [2:0]    port_state_in_6_3_1,
  input      [2:0]    port_state_in_6_3_2,
  input      [2:0]    port_state_in_6_3_3,
  input      [2:0]    port_state_in_6_3_4,
  input      [2:0]    port_state_in_6_3_5,
  input      [2:0]    port_state_in_6_3_6,
  input      [2:0]    port_state_in_6_3_7,
  input      [2:0]    port_state_in_7_0_0,
  input      [2:0]    port_state_in_7_0_1,
  input      [2:0]    port_state_in_7_0_2,
  input      [2:0]    port_state_in_7_0_3,
  input      [2:0]    port_state_in_7_0_4,
  input      [2:0]    port_state_in_7_0_5,
  input      [2:0]    port_state_in_7_0_6,
  input      [2:0]    port_state_in_7_0_7,
  input      [2:0]    port_state_in_7_1_0,
  input      [2:0]    port_state_in_7_1_1,
  input      [2:0]    port_state_in_7_1_2,
  input      [2:0]    port_state_in_7_1_3,
  input      [2:0]    port_state_in_7_1_4,
  input      [2:0]    port_state_in_7_1_5,
  input      [2:0]    port_state_in_7_1_6,
  input      [2:0]    port_state_in_7_1_7,
  input      [2:0]    port_state_in_7_2_0,
  input      [2:0]    port_state_in_7_2_1,
  input      [2:0]    port_state_in_7_2_2,
  input      [2:0]    port_state_in_7_2_3,
  input      [2:0]    port_state_in_7_2_4,
  input      [2:0]    port_state_in_7_2_5,
  input      [2:0]    port_state_in_7_2_6,
  input      [2:0]    port_state_in_7_2_7,
  input      [2:0]    port_state_in_7_3_0,
  input      [2:0]    port_state_in_7_3_1,
  input      [2:0]    port_state_in_7_3_2,
  input      [2:0]    port_state_in_7_3_3,
  input      [2:0]    port_state_in_7_3_4,
  input      [2:0]    port_state_in_7_3_5,
  input      [2:0]    port_state_in_7_3_6,
  input      [2:0]    port_state_in_7_3_7,
  input      [2:0]    port_state_in_8_0_0,
  input      [2:0]    port_state_in_8_0_1,
  input      [2:0]    port_state_in_8_0_2,
  input      [2:0]    port_state_in_8_0_3,
  input      [2:0]    port_state_in_8_0_4,
  input      [2:0]    port_state_in_8_0_5,
  input      [2:0]    port_state_in_8_0_6,
  input      [2:0]    port_state_in_8_0_7,
  input      [2:0]    port_state_in_8_1_0,
  input      [2:0]    port_state_in_8_1_1,
  input      [2:0]    port_state_in_8_1_2,
  input      [2:0]    port_state_in_8_1_3,
  input      [2:0]    port_state_in_8_1_4,
  input      [2:0]    port_state_in_8_1_5,
  input      [2:0]    port_state_in_8_1_6,
  input      [2:0]    port_state_in_8_1_7,
  input      [2:0]    port_state_in_8_2_0,
  input      [2:0]    port_state_in_8_2_1,
  input      [2:0]    port_state_in_8_2_2,
  input      [2:0]    port_state_in_8_2_3,
  input      [2:0]    port_state_in_8_2_4,
  input      [2:0]    port_state_in_8_2_5,
  input      [2:0]    port_state_in_8_2_6,
  input      [2:0]    port_state_in_8_2_7,
  input      [2:0]    port_state_in_8_3_0,
  input      [2:0]    port_state_in_8_3_1,
  input      [2:0]    port_state_in_8_3_2,
  input      [2:0]    port_state_in_8_3_3,
  input      [2:0]    port_state_in_8_3_4,
  input      [2:0]    port_state_in_8_3_5,
  input      [2:0]    port_state_in_8_3_6,
  input      [2:0]    port_state_in_8_3_7,
  input      [2:0]    port_state_in_9_0_0,
  input      [2:0]    port_state_in_9_0_1,
  input      [2:0]    port_state_in_9_0_2,
  input      [2:0]    port_state_in_9_0_3,
  input      [2:0]    port_state_in_9_0_4,
  input      [2:0]    port_state_in_9_0_5,
  input      [2:0]    port_state_in_9_0_6,
  input      [2:0]    port_state_in_9_0_7,
  input      [2:0]    port_state_in_9_1_0,
  input      [2:0]    port_state_in_9_1_1,
  input      [2:0]    port_state_in_9_1_2,
  input      [2:0]    port_state_in_9_1_3,
  input      [2:0]    port_state_in_9_1_4,
  input      [2:0]    port_state_in_9_1_5,
  input      [2:0]    port_state_in_9_1_6,
  input      [2:0]    port_state_in_9_1_7,
  input      [2:0]    port_state_in_9_2_0,
  input      [2:0]    port_state_in_9_2_1,
  input      [2:0]    port_state_in_9_2_2,
  input      [2:0]    port_state_in_9_2_3,
  input      [2:0]    port_state_in_9_2_4,
  input      [2:0]    port_state_in_9_2_5,
  input      [2:0]    port_state_in_9_2_6,
  input      [2:0]    port_state_in_9_2_7,
  input      [2:0]    port_state_in_9_3_0,
  input      [2:0]    port_state_in_9_3_1,
  input      [2:0]    port_state_in_9_3_2,
  input      [2:0]    port_state_in_9_3_3,
  input      [2:0]    port_state_in_9_3_4,
  input      [2:0]    port_state_in_9_3_5,
  input      [2:0]    port_state_in_9_3_6,
  input      [2:0]    port_state_in_9_3_7,
  input      [2:0]    port_state_in_10_0_0,
  input      [2:0]    port_state_in_10_0_1,
  input      [2:0]    port_state_in_10_0_2,
  input      [2:0]    port_state_in_10_0_3,
  input      [2:0]    port_state_in_10_0_4,
  input      [2:0]    port_state_in_10_0_5,
  input      [2:0]    port_state_in_10_0_6,
  input      [2:0]    port_state_in_10_0_7,
  input      [2:0]    port_state_in_10_1_0,
  input      [2:0]    port_state_in_10_1_1,
  input      [2:0]    port_state_in_10_1_2,
  input      [2:0]    port_state_in_10_1_3,
  input      [2:0]    port_state_in_10_1_4,
  input      [2:0]    port_state_in_10_1_5,
  input      [2:0]    port_state_in_10_1_6,
  input      [2:0]    port_state_in_10_1_7,
  input      [2:0]    port_state_in_10_2_0,
  input      [2:0]    port_state_in_10_2_1,
  input      [2:0]    port_state_in_10_2_2,
  input      [2:0]    port_state_in_10_2_3,
  input      [2:0]    port_state_in_10_2_4,
  input      [2:0]    port_state_in_10_2_5,
  input      [2:0]    port_state_in_10_2_6,
  input      [2:0]    port_state_in_10_2_7,
  input      [2:0]    port_state_in_10_3_0,
  input      [2:0]    port_state_in_10_3_1,
  input      [2:0]    port_state_in_10_3_2,
  input      [2:0]    port_state_in_10_3_3,
  input      [2:0]    port_state_in_10_3_4,
  input      [2:0]    port_state_in_10_3_5,
  input      [2:0]    port_state_in_10_3_6,
  input      [2:0]    port_state_in_10_3_7,
  input      [2:0]    port_state_in_11_0_0,
  input      [2:0]    port_state_in_11_0_1,
  input      [2:0]    port_state_in_11_0_2,
  input      [2:0]    port_state_in_11_0_3,
  input      [2:0]    port_state_in_11_0_4,
  input      [2:0]    port_state_in_11_0_5,
  input      [2:0]    port_state_in_11_0_6,
  input      [2:0]    port_state_in_11_0_7,
  input      [2:0]    port_state_in_11_1_0,
  input      [2:0]    port_state_in_11_1_1,
  input      [2:0]    port_state_in_11_1_2,
  input      [2:0]    port_state_in_11_1_3,
  input      [2:0]    port_state_in_11_1_4,
  input      [2:0]    port_state_in_11_1_5,
  input      [2:0]    port_state_in_11_1_6,
  input      [2:0]    port_state_in_11_1_7,
  input      [2:0]    port_state_in_11_2_0,
  input      [2:0]    port_state_in_11_2_1,
  input      [2:0]    port_state_in_11_2_2,
  input      [2:0]    port_state_in_11_2_3,
  input      [2:0]    port_state_in_11_2_4,
  input      [2:0]    port_state_in_11_2_5,
  input      [2:0]    port_state_in_11_2_6,
  input      [2:0]    port_state_in_11_2_7,
  input      [2:0]    port_state_in_11_3_0,
  input      [2:0]    port_state_in_11_3_1,
  input      [2:0]    port_state_in_11_3_2,
  input      [2:0]    port_state_in_11_3_3,
  input      [2:0]    port_state_in_11_3_4,
  input      [2:0]    port_state_in_11_3_5,
  input      [2:0]    port_state_in_11_3_6,
  input      [2:0]    port_state_in_11_3_7,
  input      [2:0]    port_state_in_12_0_0,
  input      [2:0]    port_state_in_12_0_1,
  input      [2:0]    port_state_in_12_0_2,
  input      [2:0]    port_state_in_12_0_3,
  input      [2:0]    port_state_in_12_0_4,
  input      [2:0]    port_state_in_12_0_5,
  input      [2:0]    port_state_in_12_0_6,
  input      [2:0]    port_state_in_12_0_7,
  input      [2:0]    port_state_in_12_1_0,
  input      [2:0]    port_state_in_12_1_1,
  input      [2:0]    port_state_in_12_1_2,
  input      [2:0]    port_state_in_12_1_3,
  input      [2:0]    port_state_in_12_1_4,
  input      [2:0]    port_state_in_12_1_5,
  input      [2:0]    port_state_in_12_1_6,
  input      [2:0]    port_state_in_12_1_7,
  input      [2:0]    port_state_in_12_2_0,
  input      [2:0]    port_state_in_12_2_1,
  input      [2:0]    port_state_in_12_2_2,
  input      [2:0]    port_state_in_12_2_3,
  input      [2:0]    port_state_in_12_2_4,
  input      [2:0]    port_state_in_12_2_5,
  input      [2:0]    port_state_in_12_2_6,
  input      [2:0]    port_state_in_12_2_7,
  input      [2:0]    port_state_in_12_3_0,
  input      [2:0]    port_state_in_12_3_1,
  input      [2:0]    port_state_in_12_3_2,
  input      [2:0]    port_state_in_12_3_3,
  input      [2:0]    port_state_in_12_3_4,
  input      [2:0]    port_state_in_12_3_5,
  input      [2:0]    port_state_in_12_3_6,
  input      [2:0]    port_state_in_12_3_7,
  input      [2:0]    port_state_in_13_0_0,
  input      [2:0]    port_state_in_13_0_1,
  input      [2:0]    port_state_in_13_0_2,
  input      [2:0]    port_state_in_13_0_3,
  input      [2:0]    port_state_in_13_0_4,
  input      [2:0]    port_state_in_13_0_5,
  input      [2:0]    port_state_in_13_0_6,
  input      [2:0]    port_state_in_13_0_7,
  input      [2:0]    port_state_in_13_1_0,
  input      [2:0]    port_state_in_13_1_1,
  input      [2:0]    port_state_in_13_1_2,
  input      [2:0]    port_state_in_13_1_3,
  input      [2:0]    port_state_in_13_1_4,
  input      [2:0]    port_state_in_13_1_5,
  input      [2:0]    port_state_in_13_1_6,
  input      [2:0]    port_state_in_13_1_7,
  input      [2:0]    port_state_in_13_2_0,
  input      [2:0]    port_state_in_13_2_1,
  input      [2:0]    port_state_in_13_2_2,
  input      [2:0]    port_state_in_13_2_3,
  input      [2:0]    port_state_in_13_2_4,
  input      [2:0]    port_state_in_13_2_5,
  input      [2:0]    port_state_in_13_2_6,
  input      [2:0]    port_state_in_13_2_7,
  input      [2:0]    port_state_in_13_3_0,
  input      [2:0]    port_state_in_13_3_1,
  input      [2:0]    port_state_in_13_3_2,
  input      [2:0]    port_state_in_13_3_3,
  input      [2:0]    port_state_in_13_3_4,
  input      [2:0]    port_state_in_13_3_5,
  input      [2:0]    port_state_in_13_3_6,
  input      [2:0]    port_state_in_13_3_7,
  input      [2:0]    port_state_in_14_0_0,
  input      [2:0]    port_state_in_14_0_1,
  input      [2:0]    port_state_in_14_0_2,
  input      [2:0]    port_state_in_14_0_3,
  input      [2:0]    port_state_in_14_0_4,
  input      [2:0]    port_state_in_14_0_5,
  input      [2:0]    port_state_in_14_0_6,
  input      [2:0]    port_state_in_14_0_7,
  input      [2:0]    port_state_in_14_1_0,
  input      [2:0]    port_state_in_14_1_1,
  input      [2:0]    port_state_in_14_1_2,
  input      [2:0]    port_state_in_14_1_3,
  input      [2:0]    port_state_in_14_1_4,
  input      [2:0]    port_state_in_14_1_5,
  input      [2:0]    port_state_in_14_1_6,
  input      [2:0]    port_state_in_14_1_7,
  input      [2:0]    port_state_in_14_2_0,
  input      [2:0]    port_state_in_14_2_1,
  input      [2:0]    port_state_in_14_2_2,
  input      [2:0]    port_state_in_14_2_3,
  input      [2:0]    port_state_in_14_2_4,
  input      [2:0]    port_state_in_14_2_5,
  input      [2:0]    port_state_in_14_2_6,
  input      [2:0]    port_state_in_14_2_7,
  input      [2:0]    port_state_in_14_3_0,
  input      [2:0]    port_state_in_14_3_1,
  input      [2:0]    port_state_in_14_3_2,
  input      [2:0]    port_state_in_14_3_3,
  input      [2:0]    port_state_in_14_3_4,
  input      [2:0]    port_state_in_14_3_5,
  input      [2:0]    port_state_in_14_3_6,
  input      [2:0]    port_state_in_14_3_7,
  input      [2:0]    port_state_in_15_0_0,
  input      [2:0]    port_state_in_15_0_1,
  input      [2:0]    port_state_in_15_0_2,
  input      [2:0]    port_state_in_15_0_3,
  input      [2:0]    port_state_in_15_0_4,
  input      [2:0]    port_state_in_15_0_5,
  input      [2:0]    port_state_in_15_0_6,
  input      [2:0]    port_state_in_15_0_7,
  input      [2:0]    port_state_in_15_1_0,
  input      [2:0]    port_state_in_15_1_1,
  input      [2:0]    port_state_in_15_1_2,
  input      [2:0]    port_state_in_15_1_3,
  input      [2:0]    port_state_in_15_1_4,
  input      [2:0]    port_state_in_15_1_5,
  input      [2:0]    port_state_in_15_1_6,
  input      [2:0]    port_state_in_15_1_7,
  input      [2:0]    port_state_in_15_2_0,
  input      [2:0]    port_state_in_15_2_1,
  input      [2:0]    port_state_in_15_2_2,
  input      [2:0]    port_state_in_15_2_3,
  input      [2:0]    port_state_in_15_2_4,
  input      [2:0]    port_state_in_15_2_5,
  input      [2:0]    port_state_in_15_2_6,
  input      [2:0]    port_state_in_15_2_7,
  input      [2:0]    port_state_in_15_3_0,
  input      [2:0]    port_state_in_15_3_1,
  input      [2:0]    port_state_in_15_3_2,
  input      [2:0]    port_state_in_15_3_3,
  input      [2:0]    port_state_in_15_3_4,
  input      [2:0]    port_state_in_15_3_5,
  input      [2:0]    port_state_in_15_3_6,
  input      [2:0]    port_state_in_15_3_7,
  input      [2:0]    port_key_0_0_0,
  input      [2:0]    port_key_0_0_1,
  input      [2:0]    port_key_0_0_2,
  input      [2:0]    port_key_0_0_3,
  input      [2:0]    port_key_0_0_4,
  input      [2:0]    port_key_0_0_5,
  input      [2:0]    port_key_0_0_6,
  input      [2:0]    port_key_0_0_7,
  input      [2:0]    port_key_0_1_0,
  input      [2:0]    port_key_0_1_1,
  input      [2:0]    port_key_0_1_2,
  input      [2:0]    port_key_0_1_3,
  input      [2:0]    port_key_0_1_4,
  input      [2:0]    port_key_0_1_5,
  input      [2:0]    port_key_0_1_6,
  input      [2:0]    port_key_0_1_7,
  input      [2:0]    port_key_0_2_0,
  input      [2:0]    port_key_0_2_1,
  input      [2:0]    port_key_0_2_2,
  input      [2:0]    port_key_0_2_3,
  input      [2:0]    port_key_0_2_4,
  input      [2:0]    port_key_0_2_5,
  input      [2:0]    port_key_0_2_6,
  input      [2:0]    port_key_0_2_7,
  input      [2:0]    port_key_0_3_0,
  input      [2:0]    port_key_0_3_1,
  input      [2:0]    port_key_0_3_2,
  input      [2:0]    port_key_0_3_3,
  input      [2:0]    port_key_0_3_4,
  input      [2:0]    port_key_0_3_5,
  input      [2:0]    port_key_0_3_6,
  input      [2:0]    port_key_0_3_7,
  input      [2:0]    port_key_1_0_0,
  input      [2:0]    port_key_1_0_1,
  input      [2:0]    port_key_1_0_2,
  input      [2:0]    port_key_1_0_3,
  input      [2:0]    port_key_1_0_4,
  input      [2:0]    port_key_1_0_5,
  input      [2:0]    port_key_1_0_6,
  input      [2:0]    port_key_1_0_7,
  input      [2:0]    port_key_1_1_0,
  input      [2:0]    port_key_1_1_1,
  input      [2:0]    port_key_1_1_2,
  input      [2:0]    port_key_1_1_3,
  input      [2:0]    port_key_1_1_4,
  input      [2:0]    port_key_1_1_5,
  input      [2:0]    port_key_1_1_6,
  input      [2:0]    port_key_1_1_7,
  input      [2:0]    port_key_1_2_0,
  input      [2:0]    port_key_1_2_1,
  input      [2:0]    port_key_1_2_2,
  input      [2:0]    port_key_1_2_3,
  input      [2:0]    port_key_1_2_4,
  input      [2:0]    port_key_1_2_5,
  input      [2:0]    port_key_1_2_6,
  input      [2:0]    port_key_1_2_7,
  input      [2:0]    port_key_1_3_0,
  input      [2:0]    port_key_1_3_1,
  input      [2:0]    port_key_1_3_2,
  input      [2:0]    port_key_1_3_3,
  input      [2:0]    port_key_1_3_4,
  input      [2:0]    port_key_1_3_5,
  input      [2:0]    port_key_1_3_6,
  input      [2:0]    port_key_1_3_7,
  input      [2:0]    port_key_2_0_0,
  input      [2:0]    port_key_2_0_1,
  input      [2:0]    port_key_2_0_2,
  input      [2:0]    port_key_2_0_3,
  input      [2:0]    port_key_2_0_4,
  input      [2:0]    port_key_2_0_5,
  input      [2:0]    port_key_2_0_6,
  input      [2:0]    port_key_2_0_7,
  input      [2:0]    port_key_2_1_0,
  input      [2:0]    port_key_2_1_1,
  input      [2:0]    port_key_2_1_2,
  input      [2:0]    port_key_2_1_3,
  input      [2:0]    port_key_2_1_4,
  input      [2:0]    port_key_2_1_5,
  input      [2:0]    port_key_2_1_6,
  input      [2:0]    port_key_2_1_7,
  input      [2:0]    port_key_2_2_0,
  input      [2:0]    port_key_2_2_1,
  input      [2:0]    port_key_2_2_2,
  input      [2:0]    port_key_2_2_3,
  input      [2:0]    port_key_2_2_4,
  input      [2:0]    port_key_2_2_5,
  input      [2:0]    port_key_2_2_6,
  input      [2:0]    port_key_2_2_7,
  input      [2:0]    port_key_2_3_0,
  input      [2:0]    port_key_2_3_1,
  input      [2:0]    port_key_2_3_2,
  input      [2:0]    port_key_2_3_3,
  input      [2:0]    port_key_2_3_4,
  input      [2:0]    port_key_2_3_5,
  input      [2:0]    port_key_2_3_6,
  input      [2:0]    port_key_2_3_7,
  input      [2:0]    port_key_3_0_0,
  input      [2:0]    port_key_3_0_1,
  input      [2:0]    port_key_3_0_2,
  input      [2:0]    port_key_3_0_3,
  input      [2:0]    port_key_3_0_4,
  input      [2:0]    port_key_3_0_5,
  input      [2:0]    port_key_3_0_6,
  input      [2:0]    port_key_3_0_7,
  input      [2:0]    port_key_3_1_0,
  input      [2:0]    port_key_3_1_1,
  input      [2:0]    port_key_3_1_2,
  input      [2:0]    port_key_3_1_3,
  input      [2:0]    port_key_3_1_4,
  input      [2:0]    port_key_3_1_5,
  input      [2:0]    port_key_3_1_6,
  input      [2:0]    port_key_3_1_7,
  input      [2:0]    port_key_3_2_0,
  input      [2:0]    port_key_3_2_1,
  input      [2:0]    port_key_3_2_2,
  input      [2:0]    port_key_3_2_3,
  input      [2:0]    port_key_3_2_4,
  input      [2:0]    port_key_3_2_5,
  input      [2:0]    port_key_3_2_6,
  input      [2:0]    port_key_3_2_7,
  input      [2:0]    port_key_3_3_0,
  input      [2:0]    port_key_3_3_1,
  input      [2:0]    port_key_3_3_2,
  input      [2:0]    port_key_3_3_3,
  input      [2:0]    port_key_3_3_4,
  input      [2:0]    port_key_3_3_5,
  input      [2:0]    port_key_3_3_6,
  input      [2:0]    port_key_3_3_7,
  input      [2:0]    port_key_4_0_0,
  input      [2:0]    port_key_4_0_1,
  input      [2:0]    port_key_4_0_2,
  input      [2:0]    port_key_4_0_3,
  input      [2:0]    port_key_4_0_4,
  input      [2:0]    port_key_4_0_5,
  input      [2:0]    port_key_4_0_6,
  input      [2:0]    port_key_4_0_7,
  input      [2:0]    port_key_4_1_0,
  input      [2:0]    port_key_4_1_1,
  input      [2:0]    port_key_4_1_2,
  input      [2:0]    port_key_4_1_3,
  input      [2:0]    port_key_4_1_4,
  input      [2:0]    port_key_4_1_5,
  input      [2:0]    port_key_4_1_6,
  input      [2:0]    port_key_4_1_7,
  input      [2:0]    port_key_4_2_0,
  input      [2:0]    port_key_4_2_1,
  input      [2:0]    port_key_4_2_2,
  input      [2:0]    port_key_4_2_3,
  input      [2:0]    port_key_4_2_4,
  input      [2:0]    port_key_4_2_5,
  input      [2:0]    port_key_4_2_6,
  input      [2:0]    port_key_4_2_7,
  input      [2:0]    port_key_4_3_0,
  input      [2:0]    port_key_4_3_1,
  input      [2:0]    port_key_4_3_2,
  input      [2:0]    port_key_4_3_3,
  input      [2:0]    port_key_4_3_4,
  input      [2:0]    port_key_4_3_5,
  input      [2:0]    port_key_4_3_6,
  input      [2:0]    port_key_4_3_7,
  input      [2:0]    port_key_5_0_0,
  input      [2:0]    port_key_5_0_1,
  input      [2:0]    port_key_5_0_2,
  input      [2:0]    port_key_5_0_3,
  input      [2:0]    port_key_5_0_4,
  input      [2:0]    port_key_5_0_5,
  input      [2:0]    port_key_5_0_6,
  input      [2:0]    port_key_5_0_7,
  input      [2:0]    port_key_5_1_0,
  input      [2:0]    port_key_5_1_1,
  input      [2:0]    port_key_5_1_2,
  input      [2:0]    port_key_5_1_3,
  input      [2:0]    port_key_5_1_4,
  input      [2:0]    port_key_5_1_5,
  input      [2:0]    port_key_5_1_6,
  input      [2:0]    port_key_5_1_7,
  input      [2:0]    port_key_5_2_0,
  input      [2:0]    port_key_5_2_1,
  input      [2:0]    port_key_5_2_2,
  input      [2:0]    port_key_5_2_3,
  input      [2:0]    port_key_5_2_4,
  input      [2:0]    port_key_5_2_5,
  input      [2:0]    port_key_5_2_6,
  input      [2:0]    port_key_5_2_7,
  input      [2:0]    port_key_5_3_0,
  input      [2:0]    port_key_5_3_1,
  input      [2:0]    port_key_5_3_2,
  input      [2:0]    port_key_5_3_3,
  input      [2:0]    port_key_5_3_4,
  input      [2:0]    port_key_5_3_5,
  input      [2:0]    port_key_5_3_6,
  input      [2:0]    port_key_5_3_7,
  input      [2:0]    port_key_6_0_0,
  input      [2:0]    port_key_6_0_1,
  input      [2:0]    port_key_6_0_2,
  input      [2:0]    port_key_6_0_3,
  input      [2:0]    port_key_6_0_4,
  input      [2:0]    port_key_6_0_5,
  input      [2:0]    port_key_6_0_6,
  input      [2:0]    port_key_6_0_7,
  input      [2:0]    port_key_6_1_0,
  input      [2:0]    port_key_6_1_1,
  input      [2:0]    port_key_6_1_2,
  input      [2:0]    port_key_6_1_3,
  input      [2:0]    port_key_6_1_4,
  input      [2:0]    port_key_6_1_5,
  input      [2:0]    port_key_6_1_6,
  input      [2:0]    port_key_6_1_7,
  input      [2:0]    port_key_6_2_0,
  input      [2:0]    port_key_6_2_1,
  input      [2:0]    port_key_6_2_2,
  input      [2:0]    port_key_6_2_3,
  input      [2:0]    port_key_6_2_4,
  input      [2:0]    port_key_6_2_5,
  input      [2:0]    port_key_6_2_6,
  input      [2:0]    port_key_6_2_7,
  input      [2:0]    port_key_6_3_0,
  input      [2:0]    port_key_6_3_1,
  input      [2:0]    port_key_6_3_2,
  input      [2:0]    port_key_6_3_3,
  input      [2:0]    port_key_6_3_4,
  input      [2:0]    port_key_6_3_5,
  input      [2:0]    port_key_6_3_6,
  input      [2:0]    port_key_6_3_7,
  input      [2:0]    port_key_7_0_0,
  input      [2:0]    port_key_7_0_1,
  input      [2:0]    port_key_7_0_2,
  input      [2:0]    port_key_7_0_3,
  input      [2:0]    port_key_7_0_4,
  input      [2:0]    port_key_7_0_5,
  input      [2:0]    port_key_7_0_6,
  input      [2:0]    port_key_7_0_7,
  input      [2:0]    port_key_7_1_0,
  input      [2:0]    port_key_7_1_1,
  input      [2:0]    port_key_7_1_2,
  input      [2:0]    port_key_7_1_3,
  input      [2:0]    port_key_7_1_4,
  input      [2:0]    port_key_7_1_5,
  input      [2:0]    port_key_7_1_6,
  input      [2:0]    port_key_7_1_7,
  input      [2:0]    port_key_7_2_0,
  input      [2:0]    port_key_7_2_1,
  input      [2:0]    port_key_7_2_2,
  input      [2:0]    port_key_7_2_3,
  input      [2:0]    port_key_7_2_4,
  input      [2:0]    port_key_7_2_5,
  input      [2:0]    port_key_7_2_6,
  input      [2:0]    port_key_7_2_7,
  input      [2:0]    port_key_7_3_0,
  input      [2:0]    port_key_7_3_1,
  input      [2:0]    port_key_7_3_2,
  input      [2:0]    port_key_7_3_3,
  input      [2:0]    port_key_7_3_4,
  input      [2:0]    port_key_7_3_5,
  input      [2:0]    port_key_7_3_6,
  input      [2:0]    port_key_7_3_7,
  input      [2:0]    port_key_8_0_0,
  input      [2:0]    port_key_8_0_1,
  input      [2:0]    port_key_8_0_2,
  input      [2:0]    port_key_8_0_3,
  input      [2:0]    port_key_8_0_4,
  input      [2:0]    port_key_8_0_5,
  input      [2:0]    port_key_8_0_6,
  input      [2:0]    port_key_8_0_7,
  input      [2:0]    port_key_8_1_0,
  input      [2:0]    port_key_8_1_1,
  input      [2:0]    port_key_8_1_2,
  input      [2:0]    port_key_8_1_3,
  input      [2:0]    port_key_8_1_4,
  input      [2:0]    port_key_8_1_5,
  input      [2:0]    port_key_8_1_6,
  input      [2:0]    port_key_8_1_7,
  input      [2:0]    port_key_8_2_0,
  input      [2:0]    port_key_8_2_1,
  input      [2:0]    port_key_8_2_2,
  input      [2:0]    port_key_8_2_3,
  input      [2:0]    port_key_8_2_4,
  input      [2:0]    port_key_8_2_5,
  input      [2:0]    port_key_8_2_6,
  input      [2:0]    port_key_8_2_7,
  input      [2:0]    port_key_8_3_0,
  input      [2:0]    port_key_8_3_1,
  input      [2:0]    port_key_8_3_2,
  input      [2:0]    port_key_8_3_3,
  input      [2:0]    port_key_8_3_4,
  input      [2:0]    port_key_8_3_5,
  input      [2:0]    port_key_8_3_6,
  input      [2:0]    port_key_8_3_7,
  input      [2:0]    port_key_9_0_0,
  input      [2:0]    port_key_9_0_1,
  input      [2:0]    port_key_9_0_2,
  input      [2:0]    port_key_9_0_3,
  input      [2:0]    port_key_9_0_4,
  input      [2:0]    port_key_9_0_5,
  input      [2:0]    port_key_9_0_6,
  input      [2:0]    port_key_9_0_7,
  input      [2:0]    port_key_9_1_0,
  input      [2:0]    port_key_9_1_1,
  input      [2:0]    port_key_9_1_2,
  input      [2:0]    port_key_9_1_3,
  input      [2:0]    port_key_9_1_4,
  input      [2:0]    port_key_9_1_5,
  input      [2:0]    port_key_9_1_6,
  input      [2:0]    port_key_9_1_7,
  input      [2:0]    port_key_9_2_0,
  input      [2:0]    port_key_9_2_1,
  input      [2:0]    port_key_9_2_2,
  input      [2:0]    port_key_9_2_3,
  input      [2:0]    port_key_9_2_4,
  input      [2:0]    port_key_9_2_5,
  input      [2:0]    port_key_9_2_6,
  input      [2:0]    port_key_9_2_7,
  input      [2:0]    port_key_9_3_0,
  input      [2:0]    port_key_9_3_1,
  input      [2:0]    port_key_9_3_2,
  input      [2:0]    port_key_9_3_3,
  input      [2:0]    port_key_9_3_4,
  input      [2:0]    port_key_9_3_5,
  input      [2:0]    port_key_9_3_6,
  input      [2:0]    port_key_9_3_7,
  input      [2:0]    port_key_10_0_0,
  input      [2:0]    port_key_10_0_1,
  input      [2:0]    port_key_10_0_2,
  input      [2:0]    port_key_10_0_3,
  input      [2:0]    port_key_10_0_4,
  input      [2:0]    port_key_10_0_5,
  input      [2:0]    port_key_10_0_6,
  input      [2:0]    port_key_10_0_7,
  input      [2:0]    port_key_10_1_0,
  input      [2:0]    port_key_10_1_1,
  input      [2:0]    port_key_10_1_2,
  input      [2:0]    port_key_10_1_3,
  input      [2:0]    port_key_10_1_4,
  input      [2:0]    port_key_10_1_5,
  input      [2:0]    port_key_10_1_6,
  input      [2:0]    port_key_10_1_7,
  input      [2:0]    port_key_10_2_0,
  input      [2:0]    port_key_10_2_1,
  input      [2:0]    port_key_10_2_2,
  input      [2:0]    port_key_10_2_3,
  input      [2:0]    port_key_10_2_4,
  input      [2:0]    port_key_10_2_5,
  input      [2:0]    port_key_10_2_6,
  input      [2:0]    port_key_10_2_7,
  input      [2:0]    port_key_10_3_0,
  input      [2:0]    port_key_10_3_1,
  input      [2:0]    port_key_10_3_2,
  input      [2:0]    port_key_10_3_3,
  input      [2:0]    port_key_10_3_4,
  input      [2:0]    port_key_10_3_5,
  input      [2:0]    port_key_10_3_6,
  input      [2:0]    port_key_10_3_7,
  input      [2:0]    port_key_11_0_0,
  input      [2:0]    port_key_11_0_1,
  input      [2:0]    port_key_11_0_2,
  input      [2:0]    port_key_11_0_3,
  input      [2:0]    port_key_11_0_4,
  input      [2:0]    port_key_11_0_5,
  input      [2:0]    port_key_11_0_6,
  input      [2:0]    port_key_11_0_7,
  input      [2:0]    port_key_11_1_0,
  input      [2:0]    port_key_11_1_1,
  input      [2:0]    port_key_11_1_2,
  input      [2:0]    port_key_11_1_3,
  input      [2:0]    port_key_11_1_4,
  input      [2:0]    port_key_11_1_5,
  input      [2:0]    port_key_11_1_6,
  input      [2:0]    port_key_11_1_7,
  input      [2:0]    port_key_11_2_0,
  input      [2:0]    port_key_11_2_1,
  input      [2:0]    port_key_11_2_2,
  input      [2:0]    port_key_11_2_3,
  input      [2:0]    port_key_11_2_4,
  input      [2:0]    port_key_11_2_5,
  input      [2:0]    port_key_11_2_6,
  input      [2:0]    port_key_11_2_7,
  input      [2:0]    port_key_11_3_0,
  input      [2:0]    port_key_11_3_1,
  input      [2:0]    port_key_11_3_2,
  input      [2:0]    port_key_11_3_3,
  input      [2:0]    port_key_11_3_4,
  input      [2:0]    port_key_11_3_5,
  input      [2:0]    port_key_11_3_6,
  input      [2:0]    port_key_11_3_7,
  input      [2:0]    port_key_12_0_0,
  input      [2:0]    port_key_12_0_1,
  input      [2:0]    port_key_12_0_2,
  input      [2:0]    port_key_12_0_3,
  input      [2:0]    port_key_12_0_4,
  input      [2:0]    port_key_12_0_5,
  input      [2:0]    port_key_12_0_6,
  input      [2:0]    port_key_12_0_7,
  input      [2:0]    port_key_12_1_0,
  input      [2:0]    port_key_12_1_1,
  input      [2:0]    port_key_12_1_2,
  input      [2:0]    port_key_12_1_3,
  input      [2:0]    port_key_12_1_4,
  input      [2:0]    port_key_12_1_5,
  input      [2:0]    port_key_12_1_6,
  input      [2:0]    port_key_12_1_7,
  input      [2:0]    port_key_12_2_0,
  input      [2:0]    port_key_12_2_1,
  input      [2:0]    port_key_12_2_2,
  input      [2:0]    port_key_12_2_3,
  input      [2:0]    port_key_12_2_4,
  input      [2:0]    port_key_12_2_5,
  input      [2:0]    port_key_12_2_6,
  input      [2:0]    port_key_12_2_7,
  input      [2:0]    port_key_12_3_0,
  input      [2:0]    port_key_12_3_1,
  input      [2:0]    port_key_12_3_2,
  input      [2:0]    port_key_12_3_3,
  input      [2:0]    port_key_12_3_4,
  input      [2:0]    port_key_12_3_5,
  input      [2:0]    port_key_12_3_6,
  input      [2:0]    port_key_12_3_7,
  input      [2:0]    port_key_13_0_0,
  input      [2:0]    port_key_13_0_1,
  input      [2:0]    port_key_13_0_2,
  input      [2:0]    port_key_13_0_3,
  input      [2:0]    port_key_13_0_4,
  input      [2:0]    port_key_13_0_5,
  input      [2:0]    port_key_13_0_6,
  input      [2:0]    port_key_13_0_7,
  input      [2:0]    port_key_13_1_0,
  input      [2:0]    port_key_13_1_1,
  input      [2:0]    port_key_13_1_2,
  input      [2:0]    port_key_13_1_3,
  input      [2:0]    port_key_13_1_4,
  input      [2:0]    port_key_13_1_5,
  input      [2:0]    port_key_13_1_6,
  input      [2:0]    port_key_13_1_7,
  input      [2:0]    port_key_13_2_0,
  input      [2:0]    port_key_13_2_1,
  input      [2:0]    port_key_13_2_2,
  input      [2:0]    port_key_13_2_3,
  input      [2:0]    port_key_13_2_4,
  input      [2:0]    port_key_13_2_5,
  input      [2:0]    port_key_13_2_6,
  input      [2:0]    port_key_13_2_7,
  input      [2:0]    port_key_13_3_0,
  input      [2:0]    port_key_13_3_1,
  input      [2:0]    port_key_13_3_2,
  input      [2:0]    port_key_13_3_3,
  input      [2:0]    port_key_13_3_4,
  input      [2:0]    port_key_13_3_5,
  input      [2:0]    port_key_13_3_6,
  input      [2:0]    port_key_13_3_7,
  input      [2:0]    port_key_14_0_0,
  input      [2:0]    port_key_14_0_1,
  input      [2:0]    port_key_14_0_2,
  input      [2:0]    port_key_14_0_3,
  input      [2:0]    port_key_14_0_4,
  input      [2:0]    port_key_14_0_5,
  input      [2:0]    port_key_14_0_6,
  input      [2:0]    port_key_14_0_7,
  input      [2:0]    port_key_14_1_0,
  input      [2:0]    port_key_14_1_1,
  input      [2:0]    port_key_14_1_2,
  input      [2:0]    port_key_14_1_3,
  input      [2:0]    port_key_14_1_4,
  input      [2:0]    port_key_14_1_5,
  input      [2:0]    port_key_14_1_6,
  input      [2:0]    port_key_14_1_7,
  input      [2:0]    port_key_14_2_0,
  input      [2:0]    port_key_14_2_1,
  input      [2:0]    port_key_14_2_2,
  input      [2:0]    port_key_14_2_3,
  input      [2:0]    port_key_14_2_4,
  input      [2:0]    port_key_14_2_5,
  input      [2:0]    port_key_14_2_6,
  input      [2:0]    port_key_14_2_7,
  input      [2:0]    port_key_14_3_0,
  input      [2:0]    port_key_14_3_1,
  input      [2:0]    port_key_14_3_2,
  input      [2:0]    port_key_14_3_3,
  input      [2:0]    port_key_14_3_4,
  input      [2:0]    port_key_14_3_5,
  input      [2:0]    port_key_14_3_6,
  input      [2:0]    port_key_14_3_7,
  input      [2:0]    port_key_15_0_0,
  input      [2:0]    port_key_15_0_1,
  input      [2:0]    port_key_15_0_2,
  input      [2:0]    port_key_15_0_3,
  input      [2:0]    port_key_15_0_4,
  input      [2:0]    port_key_15_0_5,
  input      [2:0]    port_key_15_0_6,
  input      [2:0]    port_key_15_0_7,
  input      [2:0]    port_key_15_1_0,
  input      [2:0]    port_key_15_1_1,
  input      [2:0]    port_key_15_1_2,
  input      [2:0]    port_key_15_1_3,
  input      [2:0]    port_key_15_1_4,
  input      [2:0]    port_key_15_1_5,
  input      [2:0]    port_key_15_1_6,
  input      [2:0]    port_key_15_1_7,
  input      [2:0]    port_key_15_2_0,
  input      [2:0]    port_key_15_2_1,
  input      [2:0]    port_key_15_2_2,
  input      [2:0]    port_key_15_2_3,
  input      [2:0]    port_key_15_2_4,
  input      [2:0]    port_key_15_2_5,
  input      [2:0]    port_key_15_2_6,
  input      [2:0]    port_key_15_2_7,
  input      [2:0]    port_key_15_3_0,
  input      [2:0]    port_key_15_3_1,
  input      [2:0]    port_key_15_3_2,
  input      [2:0]    port_key_15_3_3,
  input      [2:0]    port_key_15_3_4,
  input      [2:0]    port_key_15_3_5,
  input      [2:0]    port_key_15_3_6,
  input      [2:0]    port_key_15_3_7,
  output     [2:0]    port_state_out_0_0_0,
  output     [2:0]    port_state_out_0_0_1,
  output     [2:0]    port_state_out_0_0_2,
  output     [2:0]    port_state_out_0_0_3,
  output     [2:0]    port_state_out_0_0_4,
  output     [2:0]    port_state_out_0_0_5,
  output     [2:0]    port_state_out_0_0_6,
  output     [2:0]    port_state_out_0_0_7,
  output     [2:0]    port_state_out_0_1_0,
  output     [2:0]    port_state_out_0_1_1,
  output     [2:0]    port_state_out_0_1_2,
  output     [2:0]    port_state_out_0_1_3,
  output     [2:0]    port_state_out_0_1_4,
  output     [2:0]    port_state_out_0_1_5,
  output     [2:0]    port_state_out_0_1_6,
  output     [2:0]    port_state_out_0_1_7,
  output     [2:0]    port_state_out_0_2_0,
  output     [2:0]    port_state_out_0_2_1,
  output     [2:0]    port_state_out_0_2_2,
  output     [2:0]    port_state_out_0_2_3,
  output     [2:0]    port_state_out_0_2_4,
  output     [2:0]    port_state_out_0_2_5,
  output     [2:0]    port_state_out_0_2_6,
  output     [2:0]    port_state_out_0_2_7,
  output     [2:0]    port_state_out_0_3_0,
  output     [2:0]    port_state_out_0_3_1,
  output     [2:0]    port_state_out_0_3_2,
  output     [2:0]    port_state_out_0_3_3,
  output     [2:0]    port_state_out_0_3_4,
  output     [2:0]    port_state_out_0_3_5,
  output     [2:0]    port_state_out_0_3_6,
  output     [2:0]    port_state_out_0_3_7,
  output     [2:0]    port_state_out_1_0_0,
  output     [2:0]    port_state_out_1_0_1,
  output     [2:0]    port_state_out_1_0_2,
  output     [2:0]    port_state_out_1_0_3,
  output     [2:0]    port_state_out_1_0_4,
  output     [2:0]    port_state_out_1_0_5,
  output     [2:0]    port_state_out_1_0_6,
  output     [2:0]    port_state_out_1_0_7,
  output     [2:0]    port_state_out_1_1_0,
  output     [2:0]    port_state_out_1_1_1,
  output     [2:0]    port_state_out_1_1_2,
  output     [2:0]    port_state_out_1_1_3,
  output     [2:0]    port_state_out_1_1_4,
  output     [2:0]    port_state_out_1_1_5,
  output     [2:0]    port_state_out_1_1_6,
  output     [2:0]    port_state_out_1_1_7,
  output     [2:0]    port_state_out_1_2_0,
  output     [2:0]    port_state_out_1_2_1,
  output     [2:0]    port_state_out_1_2_2,
  output     [2:0]    port_state_out_1_2_3,
  output     [2:0]    port_state_out_1_2_4,
  output     [2:0]    port_state_out_1_2_5,
  output     [2:0]    port_state_out_1_2_6,
  output     [2:0]    port_state_out_1_2_7,
  output     [2:0]    port_state_out_1_3_0,
  output     [2:0]    port_state_out_1_3_1,
  output     [2:0]    port_state_out_1_3_2,
  output     [2:0]    port_state_out_1_3_3,
  output     [2:0]    port_state_out_1_3_4,
  output     [2:0]    port_state_out_1_3_5,
  output     [2:0]    port_state_out_1_3_6,
  output     [2:0]    port_state_out_1_3_7,
  output     [2:0]    port_state_out_2_0_0,
  output     [2:0]    port_state_out_2_0_1,
  output     [2:0]    port_state_out_2_0_2,
  output     [2:0]    port_state_out_2_0_3,
  output     [2:0]    port_state_out_2_0_4,
  output     [2:0]    port_state_out_2_0_5,
  output     [2:0]    port_state_out_2_0_6,
  output     [2:0]    port_state_out_2_0_7,
  output     [2:0]    port_state_out_2_1_0,
  output     [2:0]    port_state_out_2_1_1,
  output     [2:0]    port_state_out_2_1_2,
  output     [2:0]    port_state_out_2_1_3,
  output     [2:0]    port_state_out_2_1_4,
  output     [2:0]    port_state_out_2_1_5,
  output     [2:0]    port_state_out_2_1_6,
  output     [2:0]    port_state_out_2_1_7,
  output     [2:0]    port_state_out_2_2_0,
  output     [2:0]    port_state_out_2_2_1,
  output     [2:0]    port_state_out_2_2_2,
  output     [2:0]    port_state_out_2_2_3,
  output     [2:0]    port_state_out_2_2_4,
  output     [2:0]    port_state_out_2_2_5,
  output     [2:0]    port_state_out_2_2_6,
  output     [2:0]    port_state_out_2_2_7,
  output     [2:0]    port_state_out_2_3_0,
  output     [2:0]    port_state_out_2_3_1,
  output     [2:0]    port_state_out_2_3_2,
  output     [2:0]    port_state_out_2_3_3,
  output     [2:0]    port_state_out_2_3_4,
  output     [2:0]    port_state_out_2_3_5,
  output     [2:0]    port_state_out_2_3_6,
  output     [2:0]    port_state_out_2_3_7,
  output     [2:0]    port_state_out_3_0_0,
  output     [2:0]    port_state_out_3_0_1,
  output     [2:0]    port_state_out_3_0_2,
  output     [2:0]    port_state_out_3_0_3,
  output     [2:0]    port_state_out_3_0_4,
  output     [2:0]    port_state_out_3_0_5,
  output     [2:0]    port_state_out_3_0_6,
  output     [2:0]    port_state_out_3_0_7,
  output     [2:0]    port_state_out_3_1_0,
  output     [2:0]    port_state_out_3_1_1,
  output     [2:0]    port_state_out_3_1_2,
  output     [2:0]    port_state_out_3_1_3,
  output     [2:0]    port_state_out_3_1_4,
  output     [2:0]    port_state_out_3_1_5,
  output     [2:0]    port_state_out_3_1_6,
  output     [2:0]    port_state_out_3_1_7,
  output     [2:0]    port_state_out_3_2_0,
  output     [2:0]    port_state_out_3_2_1,
  output     [2:0]    port_state_out_3_2_2,
  output     [2:0]    port_state_out_3_2_3,
  output     [2:0]    port_state_out_3_2_4,
  output     [2:0]    port_state_out_3_2_5,
  output     [2:0]    port_state_out_3_2_6,
  output     [2:0]    port_state_out_3_2_7,
  output     [2:0]    port_state_out_3_3_0,
  output     [2:0]    port_state_out_3_3_1,
  output     [2:0]    port_state_out_3_3_2,
  output     [2:0]    port_state_out_3_3_3,
  output     [2:0]    port_state_out_3_3_4,
  output     [2:0]    port_state_out_3_3_5,
  output     [2:0]    port_state_out_3_3_6,
  output     [2:0]    port_state_out_3_3_7,
  output     [2:0]    port_state_out_4_0_0,
  output     [2:0]    port_state_out_4_0_1,
  output     [2:0]    port_state_out_4_0_2,
  output     [2:0]    port_state_out_4_0_3,
  output     [2:0]    port_state_out_4_0_4,
  output     [2:0]    port_state_out_4_0_5,
  output     [2:0]    port_state_out_4_0_6,
  output     [2:0]    port_state_out_4_0_7,
  output     [2:0]    port_state_out_4_1_0,
  output     [2:0]    port_state_out_4_1_1,
  output     [2:0]    port_state_out_4_1_2,
  output     [2:0]    port_state_out_4_1_3,
  output     [2:0]    port_state_out_4_1_4,
  output     [2:0]    port_state_out_4_1_5,
  output     [2:0]    port_state_out_4_1_6,
  output     [2:0]    port_state_out_4_1_7,
  output     [2:0]    port_state_out_4_2_0,
  output     [2:0]    port_state_out_4_2_1,
  output     [2:0]    port_state_out_4_2_2,
  output     [2:0]    port_state_out_4_2_3,
  output     [2:0]    port_state_out_4_2_4,
  output     [2:0]    port_state_out_4_2_5,
  output     [2:0]    port_state_out_4_2_6,
  output     [2:0]    port_state_out_4_2_7,
  output     [2:0]    port_state_out_4_3_0,
  output     [2:0]    port_state_out_4_3_1,
  output     [2:0]    port_state_out_4_3_2,
  output     [2:0]    port_state_out_4_3_3,
  output     [2:0]    port_state_out_4_3_4,
  output     [2:0]    port_state_out_4_3_5,
  output     [2:0]    port_state_out_4_3_6,
  output     [2:0]    port_state_out_4_3_7,
  output     [2:0]    port_state_out_5_0_0,
  output     [2:0]    port_state_out_5_0_1,
  output     [2:0]    port_state_out_5_0_2,
  output     [2:0]    port_state_out_5_0_3,
  output     [2:0]    port_state_out_5_0_4,
  output     [2:0]    port_state_out_5_0_5,
  output     [2:0]    port_state_out_5_0_6,
  output     [2:0]    port_state_out_5_0_7,
  output     [2:0]    port_state_out_5_1_0,
  output     [2:0]    port_state_out_5_1_1,
  output     [2:0]    port_state_out_5_1_2,
  output     [2:0]    port_state_out_5_1_3,
  output     [2:0]    port_state_out_5_1_4,
  output     [2:0]    port_state_out_5_1_5,
  output     [2:0]    port_state_out_5_1_6,
  output     [2:0]    port_state_out_5_1_7,
  output     [2:0]    port_state_out_5_2_0,
  output     [2:0]    port_state_out_5_2_1,
  output     [2:0]    port_state_out_5_2_2,
  output     [2:0]    port_state_out_5_2_3,
  output     [2:0]    port_state_out_5_2_4,
  output     [2:0]    port_state_out_5_2_5,
  output     [2:0]    port_state_out_5_2_6,
  output     [2:0]    port_state_out_5_2_7,
  output     [2:0]    port_state_out_5_3_0,
  output     [2:0]    port_state_out_5_3_1,
  output     [2:0]    port_state_out_5_3_2,
  output     [2:0]    port_state_out_5_3_3,
  output     [2:0]    port_state_out_5_3_4,
  output     [2:0]    port_state_out_5_3_5,
  output     [2:0]    port_state_out_5_3_6,
  output     [2:0]    port_state_out_5_3_7,
  output     [2:0]    port_state_out_6_0_0,
  output     [2:0]    port_state_out_6_0_1,
  output     [2:0]    port_state_out_6_0_2,
  output     [2:0]    port_state_out_6_0_3,
  output     [2:0]    port_state_out_6_0_4,
  output     [2:0]    port_state_out_6_0_5,
  output     [2:0]    port_state_out_6_0_6,
  output     [2:0]    port_state_out_6_0_7,
  output     [2:0]    port_state_out_6_1_0,
  output     [2:0]    port_state_out_6_1_1,
  output     [2:0]    port_state_out_6_1_2,
  output     [2:0]    port_state_out_6_1_3,
  output     [2:0]    port_state_out_6_1_4,
  output     [2:0]    port_state_out_6_1_5,
  output     [2:0]    port_state_out_6_1_6,
  output     [2:0]    port_state_out_6_1_7,
  output     [2:0]    port_state_out_6_2_0,
  output     [2:0]    port_state_out_6_2_1,
  output     [2:0]    port_state_out_6_2_2,
  output     [2:0]    port_state_out_6_2_3,
  output     [2:0]    port_state_out_6_2_4,
  output     [2:0]    port_state_out_6_2_5,
  output     [2:0]    port_state_out_6_2_6,
  output     [2:0]    port_state_out_6_2_7,
  output     [2:0]    port_state_out_6_3_0,
  output     [2:0]    port_state_out_6_3_1,
  output     [2:0]    port_state_out_6_3_2,
  output     [2:0]    port_state_out_6_3_3,
  output     [2:0]    port_state_out_6_3_4,
  output     [2:0]    port_state_out_6_3_5,
  output     [2:0]    port_state_out_6_3_6,
  output     [2:0]    port_state_out_6_3_7,
  output     [2:0]    port_state_out_7_0_0,
  output     [2:0]    port_state_out_7_0_1,
  output     [2:0]    port_state_out_7_0_2,
  output     [2:0]    port_state_out_7_0_3,
  output     [2:0]    port_state_out_7_0_4,
  output     [2:0]    port_state_out_7_0_5,
  output     [2:0]    port_state_out_7_0_6,
  output     [2:0]    port_state_out_7_0_7,
  output     [2:0]    port_state_out_7_1_0,
  output     [2:0]    port_state_out_7_1_1,
  output     [2:0]    port_state_out_7_1_2,
  output     [2:0]    port_state_out_7_1_3,
  output     [2:0]    port_state_out_7_1_4,
  output     [2:0]    port_state_out_7_1_5,
  output     [2:0]    port_state_out_7_1_6,
  output     [2:0]    port_state_out_7_1_7,
  output     [2:0]    port_state_out_7_2_0,
  output     [2:0]    port_state_out_7_2_1,
  output     [2:0]    port_state_out_7_2_2,
  output     [2:0]    port_state_out_7_2_3,
  output     [2:0]    port_state_out_7_2_4,
  output     [2:0]    port_state_out_7_2_5,
  output     [2:0]    port_state_out_7_2_6,
  output     [2:0]    port_state_out_7_2_7,
  output     [2:0]    port_state_out_7_3_0,
  output     [2:0]    port_state_out_7_3_1,
  output     [2:0]    port_state_out_7_3_2,
  output     [2:0]    port_state_out_7_3_3,
  output     [2:0]    port_state_out_7_3_4,
  output     [2:0]    port_state_out_7_3_5,
  output     [2:0]    port_state_out_7_3_6,
  output     [2:0]    port_state_out_7_3_7,
  output     [2:0]    port_state_out_8_0_0,
  output     [2:0]    port_state_out_8_0_1,
  output     [2:0]    port_state_out_8_0_2,
  output     [2:0]    port_state_out_8_0_3,
  output     [2:0]    port_state_out_8_0_4,
  output     [2:0]    port_state_out_8_0_5,
  output     [2:0]    port_state_out_8_0_6,
  output     [2:0]    port_state_out_8_0_7,
  output     [2:0]    port_state_out_8_1_0,
  output     [2:0]    port_state_out_8_1_1,
  output     [2:0]    port_state_out_8_1_2,
  output     [2:0]    port_state_out_8_1_3,
  output     [2:0]    port_state_out_8_1_4,
  output     [2:0]    port_state_out_8_1_5,
  output     [2:0]    port_state_out_8_1_6,
  output     [2:0]    port_state_out_8_1_7,
  output     [2:0]    port_state_out_8_2_0,
  output     [2:0]    port_state_out_8_2_1,
  output     [2:0]    port_state_out_8_2_2,
  output     [2:0]    port_state_out_8_2_3,
  output     [2:0]    port_state_out_8_2_4,
  output     [2:0]    port_state_out_8_2_5,
  output     [2:0]    port_state_out_8_2_6,
  output     [2:0]    port_state_out_8_2_7,
  output     [2:0]    port_state_out_8_3_0,
  output     [2:0]    port_state_out_8_3_1,
  output     [2:0]    port_state_out_8_3_2,
  output     [2:0]    port_state_out_8_3_3,
  output     [2:0]    port_state_out_8_3_4,
  output     [2:0]    port_state_out_8_3_5,
  output     [2:0]    port_state_out_8_3_6,
  output     [2:0]    port_state_out_8_3_7,
  output     [2:0]    port_state_out_9_0_0,
  output     [2:0]    port_state_out_9_0_1,
  output     [2:0]    port_state_out_9_0_2,
  output     [2:0]    port_state_out_9_0_3,
  output     [2:0]    port_state_out_9_0_4,
  output     [2:0]    port_state_out_9_0_5,
  output     [2:0]    port_state_out_9_0_6,
  output     [2:0]    port_state_out_9_0_7,
  output     [2:0]    port_state_out_9_1_0,
  output     [2:0]    port_state_out_9_1_1,
  output     [2:0]    port_state_out_9_1_2,
  output     [2:0]    port_state_out_9_1_3,
  output     [2:0]    port_state_out_9_1_4,
  output     [2:0]    port_state_out_9_1_5,
  output     [2:0]    port_state_out_9_1_6,
  output     [2:0]    port_state_out_9_1_7,
  output     [2:0]    port_state_out_9_2_0,
  output     [2:0]    port_state_out_9_2_1,
  output     [2:0]    port_state_out_9_2_2,
  output     [2:0]    port_state_out_9_2_3,
  output     [2:0]    port_state_out_9_2_4,
  output     [2:0]    port_state_out_9_2_5,
  output     [2:0]    port_state_out_9_2_6,
  output     [2:0]    port_state_out_9_2_7,
  output     [2:0]    port_state_out_9_3_0,
  output     [2:0]    port_state_out_9_3_1,
  output     [2:0]    port_state_out_9_3_2,
  output     [2:0]    port_state_out_9_3_3,
  output     [2:0]    port_state_out_9_3_4,
  output     [2:0]    port_state_out_9_3_5,
  output     [2:0]    port_state_out_9_3_6,
  output     [2:0]    port_state_out_9_3_7,
  output     [2:0]    port_state_out_10_0_0,
  output     [2:0]    port_state_out_10_0_1,
  output     [2:0]    port_state_out_10_0_2,
  output     [2:0]    port_state_out_10_0_3,
  output     [2:0]    port_state_out_10_0_4,
  output     [2:0]    port_state_out_10_0_5,
  output     [2:0]    port_state_out_10_0_6,
  output     [2:0]    port_state_out_10_0_7,
  output     [2:0]    port_state_out_10_1_0,
  output     [2:0]    port_state_out_10_1_1,
  output     [2:0]    port_state_out_10_1_2,
  output     [2:0]    port_state_out_10_1_3,
  output     [2:0]    port_state_out_10_1_4,
  output     [2:0]    port_state_out_10_1_5,
  output     [2:0]    port_state_out_10_1_6,
  output     [2:0]    port_state_out_10_1_7,
  output     [2:0]    port_state_out_10_2_0,
  output     [2:0]    port_state_out_10_2_1,
  output     [2:0]    port_state_out_10_2_2,
  output     [2:0]    port_state_out_10_2_3,
  output     [2:0]    port_state_out_10_2_4,
  output     [2:0]    port_state_out_10_2_5,
  output     [2:0]    port_state_out_10_2_6,
  output     [2:0]    port_state_out_10_2_7,
  output     [2:0]    port_state_out_10_3_0,
  output     [2:0]    port_state_out_10_3_1,
  output     [2:0]    port_state_out_10_3_2,
  output     [2:0]    port_state_out_10_3_3,
  output     [2:0]    port_state_out_10_3_4,
  output     [2:0]    port_state_out_10_3_5,
  output     [2:0]    port_state_out_10_3_6,
  output     [2:0]    port_state_out_10_3_7,
  output     [2:0]    port_state_out_11_0_0,
  output     [2:0]    port_state_out_11_0_1,
  output     [2:0]    port_state_out_11_0_2,
  output     [2:0]    port_state_out_11_0_3,
  output     [2:0]    port_state_out_11_0_4,
  output     [2:0]    port_state_out_11_0_5,
  output     [2:0]    port_state_out_11_0_6,
  output     [2:0]    port_state_out_11_0_7,
  output     [2:0]    port_state_out_11_1_0,
  output     [2:0]    port_state_out_11_1_1,
  output     [2:0]    port_state_out_11_1_2,
  output     [2:0]    port_state_out_11_1_3,
  output     [2:0]    port_state_out_11_1_4,
  output     [2:0]    port_state_out_11_1_5,
  output     [2:0]    port_state_out_11_1_6,
  output     [2:0]    port_state_out_11_1_7,
  output     [2:0]    port_state_out_11_2_0,
  output     [2:0]    port_state_out_11_2_1,
  output     [2:0]    port_state_out_11_2_2,
  output     [2:0]    port_state_out_11_2_3,
  output     [2:0]    port_state_out_11_2_4,
  output     [2:0]    port_state_out_11_2_5,
  output     [2:0]    port_state_out_11_2_6,
  output     [2:0]    port_state_out_11_2_7,
  output     [2:0]    port_state_out_11_3_0,
  output     [2:0]    port_state_out_11_3_1,
  output     [2:0]    port_state_out_11_3_2,
  output     [2:0]    port_state_out_11_3_3,
  output     [2:0]    port_state_out_11_3_4,
  output     [2:0]    port_state_out_11_3_5,
  output     [2:0]    port_state_out_11_3_6,
  output     [2:0]    port_state_out_11_3_7,
  output     [2:0]    port_state_out_12_0_0,
  output     [2:0]    port_state_out_12_0_1,
  output     [2:0]    port_state_out_12_0_2,
  output     [2:0]    port_state_out_12_0_3,
  output     [2:0]    port_state_out_12_0_4,
  output     [2:0]    port_state_out_12_0_5,
  output     [2:0]    port_state_out_12_0_6,
  output     [2:0]    port_state_out_12_0_7,
  output     [2:0]    port_state_out_12_1_0,
  output     [2:0]    port_state_out_12_1_1,
  output     [2:0]    port_state_out_12_1_2,
  output     [2:0]    port_state_out_12_1_3,
  output     [2:0]    port_state_out_12_1_4,
  output     [2:0]    port_state_out_12_1_5,
  output     [2:0]    port_state_out_12_1_6,
  output     [2:0]    port_state_out_12_1_7,
  output     [2:0]    port_state_out_12_2_0,
  output     [2:0]    port_state_out_12_2_1,
  output     [2:0]    port_state_out_12_2_2,
  output     [2:0]    port_state_out_12_2_3,
  output     [2:0]    port_state_out_12_2_4,
  output     [2:0]    port_state_out_12_2_5,
  output     [2:0]    port_state_out_12_2_6,
  output     [2:0]    port_state_out_12_2_7,
  output     [2:0]    port_state_out_12_3_0,
  output     [2:0]    port_state_out_12_3_1,
  output     [2:0]    port_state_out_12_3_2,
  output     [2:0]    port_state_out_12_3_3,
  output     [2:0]    port_state_out_12_3_4,
  output     [2:0]    port_state_out_12_3_5,
  output     [2:0]    port_state_out_12_3_6,
  output     [2:0]    port_state_out_12_3_7,
  output     [2:0]    port_state_out_13_0_0,
  output     [2:0]    port_state_out_13_0_1,
  output     [2:0]    port_state_out_13_0_2,
  output     [2:0]    port_state_out_13_0_3,
  output     [2:0]    port_state_out_13_0_4,
  output     [2:0]    port_state_out_13_0_5,
  output     [2:0]    port_state_out_13_0_6,
  output     [2:0]    port_state_out_13_0_7,
  output     [2:0]    port_state_out_13_1_0,
  output     [2:0]    port_state_out_13_1_1,
  output     [2:0]    port_state_out_13_1_2,
  output     [2:0]    port_state_out_13_1_3,
  output     [2:0]    port_state_out_13_1_4,
  output     [2:0]    port_state_out_13_1_5,
  output     [2:0]    port_state_out_13_1_6,
  output     [2:0]    port_state_out_13_1_7,
  output     [2:0]    port_state_out_13_2_0,
  output     [2:0]    port_state_out_13_2_1,
  output     [2:0]    port_state_out_13_2_2,
  output     [2:0]    port_state_out_13_2_3,
  output     [2:0]    port_state_out_13_2_4,
  output     [2:0]    port_state_out_13_2_5,
  output     [2:0]    port_state_out_13_2_6,
  output     [2:0]    port_state_out_13_2_7,
  output     [2:0]    port_state_out_13_3_0,
  output     [2:0]    port_state_out_13_3_1,
  output     [2:0]    port_state_out_13_3_2,
  output     [2:0]    port_state_out_13_3_3,
  output     [2:0]    port_state_out_13_3_4,
  output     [2:0]    port_state_out_13_3_5,
  output     [2:0]    port_state_out_13_3_6,
  output     [2:0]    port_state_out_13_3_7,
  output     [2:0]    port_state_out_14_0_0,
  output     [2:0]    port_state_out_14_0_1,
  output     [2:0]    port_state_out_14_0_2,
  output     [2:0]    port_state_out_14_0_3,
  output     [2:0]    port_state_out_14_0_4,
  output     [2:0]    port_state_out_14_0_5,
  output     [2:0]    port_state_out_14_0_6,
  output     [2:0]    port_state_out_14_0_7,
  output     [2:0]    port_state_out_14_1_0,
  output     [2:0]    port_state_out_14_1_1,
  output     [2:0]    port_state_out_14_1_2,
  output     [2:0]    port_state_out_14_1_3,
  output     [2:0]    port_state_out_14_1_4,
  output     [2:0]    port_state_out_14_1_5,
  output     [2:0]    port_state_out_14_1_6,
  output     [2:0]    port_state_out_14_1_7,
  output     [2:0]    port_state_out_14_2_0,
  output     [2:0]    port_state_out_14_2_1,
  output     [2:0]    port_state_out_14_2_2,
  output     [2:0]    port_state_out_14_2_3,
  output     [2:0]    port_state_out_14_2_4,
  output     [2:0]    port_state_out_14_2_5,
  output     [2:0]    port_state_out_14_2_6,
  output     [2:0]    port_state_out_14_2_7,
  output     [2:0]    port_state_out_14_3_0,
  output     [2:0]    port_state_out_14_3_1,
  output     [2:0]    port_state_out_14_3_2,
  output     [2:0]    port_state_out_14_3_3,
  output     [2:0]    port_state_out_14_3_4,
  output     [2:0]    port_state_out_14_3_5,
  output     [2:0]    port_state_out_14_3_6,
  output     [2:0]    port_state_out_14_3_7,
  output     [2:0]    port_state_out_15_0_0,
  output     [2:0]    port_state_out_15_0_1,
  output     [2:0]    port_state_out_15_0_2,
  output     [2:0]    port_state_out_15_0_3,
  output     [2:0]    port_state_out_15_0_4,
  output     [2:0]    port_state_out_15_0_5,
  output     [2:0]    port_state_out_15_0_6,
  output     [2:0]    port_state_out_15_0_7,
  output     [2:0]    port_state_out_15_1_0,
  output     [2:0]    port_state_out_15_1_1,
  output     [2:0]    port_state_out_15_1_2,
  output     [2:0]    port_state_out_15_1_3,
  output     [2:0]    port_state_out_15_1_4,
  output     [2:0]    port_state_out_15_1_5,
  output     [2:0]    port_state_out_15_1_6,
  output     [2:0]    port_state_out_15_1_7,
  output     [2:0]    port_state_out_15_2_0,
  output     [2:0]    port_state_out_15_2_1,
  output     [2:0]    port_state_out_15_2_2,
  output     [2:0]    port_state_out_15_2_3,
  output     [2:0]    port_state_out_15_2_4,
  output     [2:0]    port_state_out_15_2_5,
  output     [2:0]    port_state_out_15_2_6,
  output     [2:0]    port_state_out_15_2_7,
  output     [2:0]    port_state_out_15_3_0,
  output     [2:0]    port_state_out_15_3_1,
  output     [2:0]    port_state_out_15_3_2,
  output     [2:0]    port_state_out_15_3_3,
  output     [2:0]    port_state_out_15_3_4,
  output     [2:0]    port_state_out_15_3_5,
  output     [2:0]    port_state_out_15_3_6,
  output     [2:0]    port_state_out_15_3_7
);


  assign port_state_out_0_0_0 = (port_state_in_0_0_0 ^ port_key_0_0_0);
  assign port_state_out_0_0_1 = (port_state_in_0_0_1 ^ port_key_0_0_1);
  assign port_state_out_0_0_2 = (port_state_in_0_0_2 ^ port_key_0_0_2);
  assign port_state_out_0_0_3 = (port_state_in_0_0_3 ^ port_key_0_0_3);
  assign port_state_out_0_0_4 = (port_state_in_0_0_4 ^ port_key_0_0_4);
  assign port_state_out_0_0_5 = (port_state_in_0_0_5 ^ port_key_0_0_5);
  assign port_state_out_0_0_6 = (port_state_in_0_0_6 ^ port_key_0_0_6);
  assign port_state_out_0_0_7 = (port_state_in_0_0_7 ^ port_key_0_0_7);
  assign port_state_out_0_1_0 = (port_state_in_0_1_0 ^ port_key_0_1_0);
  assign port_state_out_0_1_1 = (port_state_in_0_1_1 ^ port_key_0_1_1);
  assign port_state_out_0_1_2 = (port_state_in_0_1_2 ^ port_key_0_1_2);
  assign port_state_out_0_1_3 = (port_state_in_0_1_3 ^ port_key_0_1_3);
  assign port_state_out_0_1_4 = (port_state_in_0_1_4 ^ port_key_0_1_4);
  assign port_state_out_0_1_5 = (port_state_in_0_1_5 ^ port_key_0_1_5);
  assign port_state_out_0_1_6 = (port_state_in_0_1_6 ^ port_key_0_1_6);
  assign port_state_out_0_1_7 = (port_state_in_0_1_7 ^ port_key_0_1_7);
  assign port_state_out_0_2_0 = (port_state_in_0_2_0 ^ port_key_0_2_0);
  assign port_state_out_0_2_1 = (port_state_in_0_2_1 ^ port_key_0_2_1);
  assign port_state_out_0_2_2 = (port_state_in_0_2_2 ^ port_key_0_2_2);
  assign port_state_out_0_2_3 = (port_state_in_0_2_3 ^ port_key_0_2_3);
  assign port_state_out_0_2_4 = (port_state_in_0_2_4 ^ port_key_0_2_4);
  assign port_state_out_0_2_5 = (port_state_in_0_2_5 ^ port_key_0_2_5);
  assign port_state_out_0_2_6 = (port_state_in_0_2_6 ^ port_key_0_2_6);
  assign port_state_out_0_2_7 = (port_state_in_0_2_7 ^ port_key_0_2_7);
  assign port_state_out_0_3_0 = (port_state_in_0_3_0 ^ port_key_0_3_0);
  assign port_state_out_0_3_1 = (port_state_in_0_3_1 ^ port_key_0_3_1);
  assign port_state_out_0_3_2 = (port_state_in_0_3_2 ^ port_key_0_3_2);
  assign port_state_out_0_3_3 = (port_state_in_0_3_3 ^ port_key_0_3_3);
  assign port_state_out_0_3_4 = (port_state_in_0_3_4 ^ port_key_0_3_4);
  assign port_state_out_0_3_5 = (port_state_in_0_3_5 ^ port_key_0_3_5);
  assign port_state_out_0_3_6 = (port_state_in_0_3_6 ^ port_key_0_3_6);
  assign port_state_out_0_3_7 = (port_state_in_0_3_7 ^ port_key_0_3_7);
  assign port_state_out_1_0_0 = (port_state_in_1_0_0 ^ port_key_1_0_0);
  assign port_state_out_1_0_1 = (port_state_in_1_0_1 ^ port_key_1_0_1);
  assign port_state_out_1_0_2 = (port_state_in_1_0_2 ^ port_key_1_0_2);
  assign port_state_out_1_0_3 = (port_state_in_1_0_3 ^ port_key_1_0_3);
  assign port_state_out_1_0_4 = (port_state_in_1_0_4 ^ port_key_1_0_4);
  assign port_state_out_1_0_5 = (port_state_in_1_0_5 ^ port_key_1_0_5);
  assign port_state_out_1_0_6 = (port_state_in_1_0_6 ^ port_key_1_0_6);
  assign port_state_out_1_0_7 = (port_state_in_1_0_7 ^ port_key_1_0_7);
  assign port_state_out_1_1_0 = (port_state_in_1_1_0 ^ port_key_1_1_0);
  assign port_state_out_1_1_1 = (port_state_in_1_1_1 ^ port_key_1_1_1);
  assign port_state_out_1_1_2 = (port_state_in_1_1_2 ^ port_key_1_1_2);
  assign port_state_out_1_1_3 = (port_state_in_1_1_3 ^ port_key_1_1_3);
  assign port_state_out_1_1_4 = (port_state_in_1_1_4 ^ port_key_1_1_4);
  assign port_state_out_1_1_5 = (port_state_in_1_1_5 ^ port_key_1_1_5);
  assign port_state_out_1_1_6 = (port_state_in_1_1_6 ^ port_key_1_1_6);
  assign port_state_out_1_1_7 = (port_state_in_1_1_7 ^ port_key_1_1_7);
  assign port_state_out_1_2_0 = (port_state_in_1_2_0 ^ port_key_1_2_0);
  assign port_state_out_1_2_1 = (port_state_in_1_2_1 ^ port_key_1_2_1);
  assign port_state_out_1_2_2 = (port_state_in_1_2_2 ^ port_key_1_2_2);
  assign port_state_out_1_2_3 = (port_state_in_1_2_3 ^ port_key_1_2_3);
  assign port_state_out_1_2_4 = (port_state_in_1_2_4 ^ port_key_1_2_4);
  assign port_state_out_1_2_5 = (port_state_in_1_2_5 ^ port_key_1_2_5);
  assign port_state_out_1_2_6 = (port_state_in_1_2_6 ^ port_key_1_2_6);
  assign port_state_out_1_2_7 = (port_state_in_1_2_7 ^ port_key_1_2_7);
  assign port_state_out_1_3_0 = (port_state_in_1_3_0 ^ port_key_1_3_0);
  assign port_state_out_1_3_1 = (port_state_in_1_3_1 ^ port_key_1_3_1);
  assign port_state_out_1_3_2 = (port_state_in_1_3_2 ^ port_key_1_3_2);
  assign port_state_out_1_3_3 = (port_state_in_1_3_3 ^ port_key_1_3_3);
  assign port_state_out_1_3_4 = (port_state_in_1_3_4 ^ port_key_1_3_4);
  assign port_state_out_1_3_5 = (port_state_in_1_3_5 ^ port_key_1_3_5);
  assign port_state_out_1_3_6 = (port_state_in_1_3_6 ^ port_key_1_3_6);
  assign port_state_out_1_3_7 = (port_state_in_1_3_7 ^ port_key_1_3_7);
  assign port_state_out_2_0_0 = (port_state_in_2_0_0 ^ port_key_2_0_0);
  assign port_state_out_2_0_1 = (port_state_in_2_0_1 ^ port_key_2_0_1);
  assign port_state_out_2_0_2 = (port_state_in_2_0_2 ^ port_key_2_0_2);
  assign port_state_out_2_0_3 = (port_state_in_2_0_3 ^ port_key_2_0_3);
  assign port_state_out_2_0_4 = (port_state_in_2_0_4 ^ port_key_2_0_4);
  assign port_state_out_2_0_5 = (port_state_in_2_0_5 ^ port_key_2_0_5);
  assign port_state_out_2_0_6 = (port_state_in_2_0_6 ^ port_key_2_0_6);
  assign port_state_out_2_0_7 = (port_state_in_2_0_7 ^ port_key_2_0_7);
  assign port_state_out_2_1_0 = (port_state_in_2_1_0 ^ port_key_2_1_0);
  assign port_state_out_2_1_1 = (port_state_in_2_1_1 ^ port_key_2_1_1);
  assign port_state_out_2_1_2 = (port_state_in_2_1_2 ^ port_key_2_1_2);
  assign port_state_out_2_1_3 = (port_state_in_2_1_3 ^ port_key_2_1_3);
  assign port_state_out_2_1_4 = (port_state_in_2_1_4 ^ port_key_2_1_4);
  assign port_state_out_2_1_5 = (port_state_in_2_1_5 ^ port_key_2_1_5);
  assign port_state_out_2_1_6 = (port_state_in_2_1_6 ^ port_key_2_1_6);
  assign port_state_out_2_1_7 = (port_state_in_2_1_7 ^ port_key_2_1_7);
  assign port_state_out_2_2_0 = (port_state_in_2_2_0 ^ port_key_2_2_0);
  assign port_state_out_2_2_1 = (port_state_in_2_2_1 ^ port_key_2_2_1);
  assign port_state_out_2_2_2 = (port_state_in_2_2_2 ^ port_key_2_2_2);
  assign port_state_out_2_2_3 = (port_state_in_2_2_3 ^ port_key_2_2_3);
  assign port_state_out_2_2_4 = (port_state_in_2_2_4 ^ port_key_2_2_4);
  assign port_state_out_2_2_5 = (port_state_in_2_2_5 ^ port_key_2_2_5);
  assign port_state_out_2_2_6 = (port_state_in_2_2_6 ^ port_key_2_2_6);
  assign port_state_out_2_2_7 = (port_state_in_2_2_7 ^ port_key_2_2_7);
  assign port_state_out_2_3_0 = (port_state_in_2_3_0 ^ port_key_2_3_0);
  assign port_state_out_2_3_1 = (port_state_in_2_3_1 ^ port_key_2_3_1);
  assign port_state_out_2_3_2 = (port_state_in_2_3_2 ^ port_key_2_3_2);
  assign port_state_out_2_3_3 = (port_state_in_2_3_3 ^ port_key_2_3_3);
  assign port_state_out_2_3_4 = (port_state_in_2_3_4 ^ port_key_2_3_4);
  assign port_state_out_2_3_5 = (port_state_in_2_3_5 ^ port_key_2_3_5);
  assign port_state_out_2_3_6 = (port_state_in_2_3_6 ^ port_key_2_3_6);
  assign port_state_out_2_3_7 = (port_state_in_2_3_7 ^ port_key_2_3_7);
  assign port_state_out_3_0_0 = (port_state_in_3_0_0 ^ port_key_3_0_0);
  assign port_state_out_3_0_1 = (port_state_in_3_0_1 ^ port_key_3_0_1);
  assign port_state_out_3_0_2 = (port_state_in_3_0_2 ^ port_key_3_0_2);
  assign port_state_out_3_0_3 = (port_state_in_3_0_3 ^ port_key_3_0_3);
  assign port_state_out_3_0_4 = (port_state_in_3_0_4 ^ port_key_3_0_4);
  assign port_state_out_3_0_5 = (port_state_in_3_0_5 ^ port_key_3_0_5);
  assign port_state_out_3_0_6 = (port_state_in_3_0_6 ^ port_key_3_0_6);
  assign port_state_out_3_0_7 = (port_state_in_3_0_7 ^ port_key_3_0_7);
  assign port_state_out_3_1_0 = (port_state_in_3_1_0 ^ port_key_3_1_0);
  assign port_state_out_3_1_1 = (port_state_in_3_1_1 ^ port_key_3_1_1);
  assign port_state_out_3_1_2 = (port_state_in_3_1_2 ^ port_key_3_1_2);
  assign port_state_out_3_1_3 = (port_state_in_3_1_3 ^ port_key_3_1_3);
  assign port_state_out_3_1_4 = (port_state_in_3_1_4 ^ port_key_3_1_4);
  assign port_state_out_3_1_5 = (port_state_in_3_1_5 ^ port_key_3_1_5);
  assign port_state_out_3_1_6 = (port_state_in_3_1_6 ^ port_key_3_1_6);
  assign port_state_out_3_1_7 = (port_state_in_3_1_7 ^ port_key_3_1_7);
  assign port_state_out_3_2_0 = (port_state_in_3_2_0 ^ port_key_3_2_0);
  assign port_state_out_3_2_1 = (port_state_in_3_2_1 ^ port_key_3_2_1);
  assign port_state_out_3_2_2 = (port_state_in_3_2_2 ^ port_key_3_2_2);
  assign port_state_out_3_2_3 = (port_state_in_3_2_3 ^ port_key_3_2_3);
  assign port_state_out_3_2_4 = (port_state_in_3_2_4 ^ port_key_3_2_4);
  assign port_state_out_3_2_5 = (port_state_in_3_2_5 ^ port_key_3_2_5);
  assign port_state_out_3_2_6 = (port_state_in_3_2_6 ^ port_key_3_2_6);
  assign port_state_out_3_2_7 = (port_state_in_3_2_7 ^ port_key_3_2_7);
  assign port_state_out_3_3_0 = (port_state_in_3_3_0 ^ port_key_3_3_0);
  assign port_state_out_3_3_1 = (port_state_in_3_3_1 ^ port_key_3_3_1);
  assign port_state_out_3_3_2 = (port_state_in_3_3_2 ^ port_key_3_3_2);
  assign port_state_out_3_3_3 = (port_state_in_3_3_3 ^ port_key_3_3_3);
  assign port_state_out_3_3_4 = (port_state_in_3_3_4 ^ port_key_3_3_4);
  assign port_state_out_3_3_5 = (port_state_in_3_3_5 ^ port_key_3_3_5);
  assign port_state_out_3_3_6 = (port_state_in_3_3_6 ^ port_key_3_3_6);
  assign port_state_out_3_3_7 = (port_state_in_3_3_7 ^ port_key_3_3_7);
  assign port_state_out_4_0_0 = (port_state_in_4_0_0 ^ port_key_4_0_0);
  assign port_state_out_4_0_1 = (port_state_in_4_0_1 ^ port_key_4_0_1);
  assign port_state_out_4_0_2 = (port_state_in_4_0_2 ^ port_key_4_0_2);
  assign port_state_out_4_0_3 = (port_state_in_4_0_3 ^ port_key_4_0_3);
  assign port_state_out_4_0_4 = (port_state_in_4_0_4 ^ port_key_4_0_4);
  assign port_state_out_4_0_5 = (port_state_in_4_0_5 ^ port_key_4_0_5);
  assign port_state_out_4_0_6 = (port_state_in_4_0_6 ^ port_key_4_0_6);
  assign port_state_out_4_0_7 = (port_state_in_4_0_7 ^ port_key_4_0_7);
  assign port_state_out_4_1_0 = (port_state_in_4_1_0 ^ port_key_4_1_0);
  assign port_state_out_4_1_1 = (port_state_in_4_1_1 ^ port_key_4_1_1);
  assign port_state_out_4_1_2 = (port_state_in_4_1_2 ^ port_key_4_1_2);
  assign port_state_out_4_1_3 = (port_state_in_4_1_3 ^ port_key_4_1_3);
  assign port_state_out_4_1_4 = (port_state_in_4_1_4 ^ port_key_4_1_4);
  assign port_state_out_4_1_5 = (port_state_in_4_1_5 ^ port_key_4_1_5);
  assign port_state_out_4_1_6 = (port_state_in_4_1_6 ^ port_key_4_1_6);
  assign port_state_out_4_1_7 = (port_state_in_4_1_7 ^ port_key_4_1_7);
  assign port_state_out_4_2_0 = (port_state_in_4_2_0 ^ port_key_4_2_0);
  assign port_state_out_4_2_1 = (port_state_in_4_2_1 ^ port_key_4_2_1);
  assign port_state_out_4_2_2 = (port_state_in_4_2_2 ^ port_key_4_2_2);
  assign port_state_out_4_2_3 = (port_state_in_4_2_3 ^ port_key_4_2_3);
  assign port_state_out_4_2_4 = (port_state_in_4_2_4 ^ port_key_4_2_4);
  assign port_state_out_4_2_5 = (port_state_in_4_2_5 ^ port_key_4_2_5);
  assign port_state_out_4_2_6 = (port_state_in_4_2_6 ^ port_key_4_2_6);
  assign port_state_out_4_2_7 = (port_state_in_4_2_7 ^ port_key_4_2_7);
  assign port_state_out_4_3_0 = (port_state_in_4_3_0 ^ port_key_4_3_0);
  assign port_state_out_4_3_1 = (port_state_in_4_3_1 ^ port_key_4_3_1);
  assign port_state_out_4_3_2 = (port_state_in_4_3_2 ^ port_key_4_3_2);
  assign port_state_out_4_3_3 = (port_state_in_4_3_3 ^ port_key_4_3_3);
  assign port_state_out_4_3_4 = (port_state_in_4_3_4 ^ port_key_4_3_4);
  assign port_state_out_4_3_5 = (port_state_in_4_3_5 ^ port_key_4_3_5);
  assign port_state_out_4_3_6 = (port_state_in_4_3_6 ^ port_key_4_3_6);
  assign port_state_out_4_3_7 = (port_state_in_4_3_7 ^ port_key_4_3_7);
  assign port_state_out_5_0_0 = (port_state_in_5_0_0 ^ port_key_5_0_0);
  assign port_state_out_5_0_1 = (port_state_in_5_0_1 ^ port_key_5_0_1);
  assign port_state_out_5_0_2 = (port_state_in_5_0_2 ^ port_key_5_0_2);
  assign port_state_out_5_0_3 = (port_state_in_5_0_3 ^ port_key_5_0_3);
  assign port_state_out_5_0_4 = (port_state_in_5_0_4 ^ port_key_5_0_4);
  assign port_state_out_5_0_5 = (port_state_in_5_0_5 ^ port_key_5_0_5);
  assign port_state_out_5_0_6 = (port_state_in_5_0_6 ^ port_key_5_0_6);
  assign port_state_out_5_0_7 = (port_state_in_5_0_7 ^ port_key_5_0_7);
  assign port_state_out_5_1_0 = (port_state_in_5_1_0 ^ port_key_5_1_0);
  assign port_state_out_5_1_1 = (port_state_in_5_1_1 ^ port_key_5_1_1);
  assign port_state_out_5_1_2 = (port_state_in_5_1_2 ^ port_key_5_1_2);
  assign port_state_out_5_1_3 = (port_state_in_5_1_3 ^ port_key_5_1_3);
  assign port_state_out_5_1_4 = (port_state_in_5_1_4 ^ port_key_5_1_4);
  assign port_state_out_5_1_5 = (port_state_in_5_1_5 ^ port_key_5_1_5);
  assign port_state_out_5_1_6 = (port_state_in_5_1_6 ^ port_key_5_1_6);
  assign port_state_out_5_1_7 = (port_state_in_5_1_7 ^ port_key_5_1_7);
  assign port_state_out_5_2_0 = (port_state_in_5_2_0 ^ port_key_5_2_0);
  assign port_state_out_5_2_1 = (port_state_in_5_2_1 ^ port_key_5_2_1);
  assign port_state_out_5_2_2 = (port_state_in_5_2_2 ^ port_key_5_2_2);
  assign port_state_out_5_2_3 = (port_state_in_5_2_3 ^ port_key_5_2_3);
  assign port_state_out_5_2_4 = (port_state_in_5_2_4 ^ port_key_5_2_4);
  assign port_state_out_5_2_5 = (port_state_in_5_2_5 ^ port_key_5_2_5);
  assign port_state_out_5_2_6 = (port_state_in_5_2_6 ^ port_key_5_2_6);
  assign port_state_out_5_2_7 = (port_state_in_5_2_7 ^ port_key_5_2_7);
  assign port_state_out_5_3_0 = (port_state_in_5_3_0 ^ port_key_5_3_0);
  assign port_state_out_5_3_1 = (port_state_in_5_3_1 ^ port_key_5_3_1);
  assign port_state_out_5_3_2 = (port_state_in_5_3_2 ^ port_key_5_3_2);
  assign port_state_out_5_3_3 = (port_state_in_5_3_3 ^ port_key_5_3_3);
  assign port_state_out_5_3_4 = (port_state_in_5_3_4 ^ port_key_5_3_4);
  assign port_state_out_5_3_5 = (port_state_in_5_3_5 ^ port_key_5_3_5);
  assign port_state_out_5_3_6 = (port_state_in_5_3_6 ^ port_key_5_3_6);
  assign port_state_out_5_3_7 = (port_state_in_5_3_7 ^ port_key_5_3_7);
  assign port_state_out_6_0_0 = (port_state_in_6_0_0 ^ port_key_6_0_0);
  assign port_state_out_6_0_1 = (port_state_in_6_0_1 ^ port_key_6_0_1);
  assign port_state_out_6_0_2 = (port_state_in_6_0_2 ^ port_key_6_0_2);
  assign port_state_out_6_0_3 = (port_state_in_6_0_3 ^ port_key_6_0_3);
  assign port_state_out_6_0_4 = (port_state_in_6_0_4 ^ port_key_6_0_4);
  assign port_state_out_6_0_5 = (port_state_in_6_0_5 ^ port_key_6_0_5);
  assign port_state_out_6_0_6 = (port_state_in_6_0_6 ^ port_key_6_0_6);
  assign port_state_out_6_0_7 = (port_state_in_6_0_7 ^ port_key_6_0_7);
  assign port_state_out_6_1_0 = (port_state_in_6_1_0 ^ port_key_6_1_0);
  assign port_state_out_6_1_1 = (port_state_in_6_1_1 ^ port_key_6_1_1);
  assign port_state_out_6_1_2 = (port_state_in_6_1_2 ^ port_key_6_1_2);
  assign port_state_out_6_1_3 = (port_state_in_6_1_3 ^ port_key_6_1_3);
  assign port_state_out_6_1_4 = (port_state_in_6_1_4 ^ port_key_6_1_4);
  assign port_state_out_6_1_5 = (port_state_in_6_1_5 ^ port_key_6_1_5);
  assign port_state_out_6_1_6 = (port_state_in_6_1_6 ^ port_key_6_1_6);
  assign port_state_out_6_1_7 = (port_state_in_6_1_7 ^ port_key_6_1_7);
  assign port_state_out_6_2_0 = (port_state_in_6_2_0 ^ port_key_6_2_0);
  assign port_state_out_6_2_1 = (port_state_in_6_2_1 ^ port_key_6_2_1);
  assign port_state_out_6_2_2 = (port_state_in_6_2_2 ^ port_key_6_2_2);
  assign port_state_out_6_2_3 = (port_state_in_6_2_3 ^ port_key_6_2_3);
  assign port_state_out_6_2_4 = (port_state_in_6_2_4 ^ port_key_6_2_4);
  assign port_state_out_6_2_5 = (port_state_in_6_2_5 ^ port_key_6_2_5);
  assign port_state_out_6_2_6 = (port_state_in_6_2_6 ^ port_key_6_2_6);
  assign port_state_out_6_2_7 = (port_state_in_6_2_7 ^ port_key_6_2_7);
  assign port_state_out_6_3_0 = (port_state_in_6_3_0 ^ port_key_6_3_0);
  assign port_state_out_6_3_1 = (port_state_in_6_3_1 ^ port_key_6_3_1);
  assign port_state_out_6_3_2 = (port_state_in_6_3_2 ^ port_key_6_3_2);
  assign port_state_out_6_3_3 = (port_state_in_6_3_3 ^ port_key_6_3_3);
  assign port_state_out_6_3_4 = (port_state_in_6_3_4 ^ port_key_6_3_4);
  assign port_state_out_6_3_5 = (port_state_in_6_3_5 ^ port_key_6_3_5);
  assign port_state_out_6_3_6 = (port_state_in_6_3_6 ^ port_key_6_3_6);
  assign port_state_out_6_3_7 = (port_state_in_6_3_7 ^ port_key_6_3_7);
  assign port_state_out_7_0_0 = (port_state_in_7_0_0 ^ port_key_7_0_0);
  assign port_state_out_7_0_1 = (port_state_in_7_0_1 ^ port_key_7_0_1);
  assign port_state_out_7_0_2 = (port_state_in_7_0_2 ^ port_key_7_0_2);
  assign port_state_out_7_0_3 = (port_state_in_7_0_3 ^ port_key_7_0_3);
  assign port_state_out_7_0_4 = (port_state_in_7_0_4 ^ port_key_7_0_4);
  assign port_state_out_7_0_5 = (port_state_in_7_0_5 ^ port_key_7_0_5);
  assign port_state_out_7_0_6 = (port_state_in_7_0_6 ^ port_key_7_0_6);
  assign port_state_out_7_0_7 = (port_state_in_7_0_7 ^ port_key_7_0_7);
  assign port_state_out_7_1_0 = (port_state_in_7_1_0 ^ port_key_7_1_0);
  assign port_state_out_7_1_1 = (port_state_in_7_1_1 ^ port_key_7_1_1);
  assign port_state_out_7_1_2 = (port_state_in_7_1_2 ^ port_key_7_1_2);
  assign port_state_out_7_1_3 = (port_state_in_7_1_3 ^ port_key_7_1_3);
  assign port_state_out_7_1_4 = (port_state_in_7_1_4 ^ port_key_7_1_4);
  assign port_state_out_7_1_5 = (port_state_in_7_1_5 ^ port_key_7_1_5);
  assign port_state_out_7_1_6 = (port_state_in_7_1_6 ^ port_key_7_1_6);
  assign port_state_out_7_1_7 = (port_state_in_7_1_7 ^ port_key_7_1_7);
  assign port_state_out_7_2_0 = (port_state_in_7_2_0 ^ port_key_7_2_0);
  assign port_state_out_7_2_1 = (port_state_in_7_2_1 ^ port_key_7_2_1);
  assign port_state_out_7_2_2 = (port_state_in_7_2_2 ^ port_key_7_2_2);
  assign port_state_out_7_2_3 = (port_state_in_7_2_3 ^ port_key_7_2_3);
  assign port_state_out_7_2_4 = (port_state_in_7_2_4 ^ port_key_7_2_4);
  assign port_state_out_7_2_5 = (port_state_in_7_2_5 ^ port_key_7_2_5);
  assign port_state_out_7_2_6 = (port_state_in_7_2_6 ^ port_key_7_2_6);
  assign port_state_out_7_2_7 = (port_state_in_7_2_7 ^ port_key_7_2_7);
  assign port_state_out_7_3_0 = (port_state_in_7_3_0 ^ port_key_7_3_0);
  assign port_state_out_7_3_1 = (port_state_in_7_3_1 ^ port_key_7_3_1);
  assign port_state_out_7_3_2 = (port_state_in_7_3_2 ^ port_key_7_3_2);
  assign port_state_out_7_3_3 = (port_state_in_7_3_3 ^ port_key_7_3_3);
  assign port_state_out_7_3_4 = (port_state_in_7_3_4 ^ port_key_7_3_4);
  assign port_state_out_7_3_5 = (port_state_in_7_3_5 ^ port_key_7_3_5);
  assign port_state_out_7_3_6 = (port_state_in_7_3_6 ^ port_key_7_3_6);
  assign port_state_out_7_3_7 = (port_state_in_7_3_7 ^ port_key_7_3_7);
  assign port_state_out_8_0_0 = (port_state_in_8_0_0 ^ port_key_8_0_0);
  assign port_state_out_8_0_1 = (port_state_in_8_0_1 ^ port_key_8_0_1);
  assign port_state_out_8_0_2 = (port_state_in_8_0_2 ^ port_key_8_0_2);
  assign port_state_out_8_0_3 = (port_state_in_8_0_3 ^ port_key_8_0_3);
  assign port_state_out_8_0_4 = (port_state_in_8_0_4 ^ port_key_8_0_4);
  assign port_state_out_8_0_5 = (port_state_in_8_0_5 ^ port_key_8_0_5);
  assign port_state_out_8_0_6 = (port_state_in_8_0_6 ^ port_key_8_0_6);
  assign port_state_out_8_0_7 = (port_state_in_8_0_7 ^ port_key_8_0_7);
  assign port_state_out_8_1_0 = (port_state_in_8_1_0 ^ port_key_8_1_0);
  assign port_state_out_8_1_1 = (port_state_in_8_1_1 ^ port_key_8_1_1);
  assign port_state_out_8_1_2 = (port_state_in_8_1_2 ^ port_key_8_1_2);
  assign port_state_out_8_1_3 = (port_state_in_8_1_3 ^ port_key_8_1_3);
  assign port_state_out_8_1_4 = (port_state_in_8_1_4 ^ port_key_8_1_4);
  assign port_state_out_8_1_5 = (port_state_in_8_1_5 ^ port_key_8_1_5);
  assign port_state_out_8_1_6 = (port_state_in_8_1_6 ^ port_key_8_1_6);
  assign port_state_out_8_1_7 = (port_state_in_8_1_7 ^ port_key_8_1_7);
  assign port_state_out_8_2_0 = (port_state_in_8_2_0 ^ port_key_8_2_0);
  assign port_state_out_8_2_1 = (port_state_in_8_2_1 ^ port_key_8_2_1);
  assign port_state_out_8_2_2 = (port_state_in_8_2_2 ^ port_key_8_2_2);
  assign port_state_out_8_2_3 = (port_state_in_8_2_3 ^ port_key_8_2_3);
  assign port_state_out_8_2_4 = (port_state_in_8_2_4 ^ port_key_8_2_4);
  assign port_state_out_8_2_5 = (port_state_in_8_2_5 ^ port_key_8_2_5);
  assign port_state_out_8_2_6 = (port_state_in_8_2_6 ^ port_key_8_2_6);
  assign port_state_out_8_2_7 = (port_state_in_8_2_7 ^ port_key_8_2_7);
  assign port_state_out_8_3_0 = (port_state_in_8_3_0 ^ port_key_8_3_0);
  assign port_state_out_8_3_1 = (port_state_in_8_3_1 ^ port_key_8_3_1);
  assign port_state_out_8_3_2 = (port_state_in_8_3_2 ^ port_key_8_3_2);
  assign port_state_out_8_3_3 = (port_state_in_8_3_3 ^ port_key_8_3_3);
  assign port_state_out_8_3_4 = (port_state_in_8_3_4 ^ port_key_8_3_4);
  assign port_state_out_8_3_5 = (port_state_in_8_3_5 ^ port_key_8_3_5);
  assign port_state_out_8_3_6 = (port_state_in_8_3_6 ^ port_key_8_3_6);
  assign port_state_out_8_3_7 = (port_state_in_8_3_7 ^ port_key_8_3_7);
  assign port_state_out_9_0_0 = (port_state_in_9_0_0 ^ port_key_9_0_0);
  assign port_state_out_9_0_1 = (port_state_in_9_0_1 ^ port_key_9_0_1);
  assign port_state_out_9_0_2 = (port_state_in_9_0_2 ^ port_key_9_0_2);
  assign port_state_out_9_0_3 = (port_state_in_9_0_3 ^ port_key_9_0_3);
  assign port_state_out_9_0_4 = (port_state_in_9_0_4 ^ port_key_9_0_4);
  assign port_state_out_9_0_5 = (port_state_in_9_0_5 ^ port_key_9_0_5);
  assign port_state_out_9_0_6 = (port_state_in_9_0_6 ^ port_key_9_0_6);
  assign port_state_out_9_0_7 = (port_state_in_9_0_7 ^ port_key_9_0_7);
  assign port_state_out_9_1_0 = (port_state_in_9_1_0 ^ port_key_9_1_0);
  assign port_state_out_9_1_1 = (port_state_in_9_1_1 ^ port_key_9_1_1);
  assign port_state_out_9_1_2 = (port_state_in_9_1_2 ^ port_key_9_1_2);
  assign port_state_out_9_1_3 = (port_state_in_9_1_3 ^ port_key_9_1_3);
  assign port_state_out_9_1_4 = (port_state_in_9_1_4 ^ port_key_9_1_4);
  assign port_state_out_9_1_5 = (port_state_in_9_1_5 ^ port_key_9_1_5);
  assign port_state_out_9_1_6 = (port_state_in_9_1_6 ^ port_key_9_1_6);
  assign port_state_out_9_1_7 = (port_state_in_9_1_7 ^ port_key_9_1_7);
  assign port_state_out_9_2_0 = (port_state_in_9_2_0 ^ port_key_9_2_0);
  assign port_state_out_9_2_1 = (port_state_in_9_2_1 ^ port_key_9_2_1);
  assign port_state_out_9_2_2 = (port_state_in_9_2_2 ^ port_key_9_2_2);
  assign port_state_out_9_2_3 = (port_state_in_9_2_3 ^ port_key_9_2_3);
  assign port_state_out_9_2_4 = (port_state_in_9_2_4 ^ port_key_9_2_4);
  assign port_state_out_9_2_5 = (port_state_in_9_2_5 ^ port_key_9_2_5);
  assign port_state_out_9_2_6 = (port_state_in_9_2_6 ^ port_key_9_2_6);
  assign port_state_out_9_2_7 = (port_state_in_9_2_7 ^ port_key_9_2_7);
  assign port_state_out_9_3_0 = (port_state_in_9_3_0 ^ port_key_9_3_0);
  assign port_state_out_9_3_1 = (port_state_in_9_3_1 ^ port_key_9_3_1);
  assign port_state_out_9_3_2 = (port_state_in_9_3_2 ^ port_key_9_3_2);
  assign port_state_out_9_3_3 = (port_state_in_9_3_3 ^ port_key_9_3_3);
  assign port_state_out_9_3_4 = (port_state_in_9_3_4 ^ port_key_9_3_4);
  assign port_state_out_9_3_5 = (port_state_in_9_3_5 ^ port_key_9_3_5);
  assign port_state_out_9_3_6 = (port_state_in_9_3_6 ^ port_key_9_3_6);
  assign port_state_out_9_3_7 = (port_state_in_9_3_7 ^ port_key_9_3_7);
  assign port_state_out_10_0_0 = (port_state_in_10_0_0 ^ port_key_10_0_0);
  assign port_state_out_10_0_1 = (port_state_in_10_0_1 ^ port_key_10_0_1);
  assign port_state_out_10_0_2 = (port_state_in_10_0_2 ^ port_key_10_0_2);
  assign port_state_out_10_0_3 = (port_state_in_10_0_3 ^ port_key_10_0_3);
  assign port_state_out_10_0_4 = (port_state_in_10_0_4 ^ port_key_10_0_4);
  assign port_state_out_10_0_5 = (port_state_in_10_0_5 ^ port_key_10_0_5);
  assign port_state_out_10_0_6 = (port_state_in_10_0_6 ^ port_key_10_0_6);
  assign port_state_out_10_0_7 = (port_state_in_10_0_7 ^ port_key_10_0_7);
  assign port_state_out_10_1_0 = (port_state_in_10_1_0 ^ port_key_10_1_0);
  assign port_state_out_10_1_1 = (port_state_in_10_1_1 ^ port_key_10_1_1);
  assign port_state_out_10_1_2 = (port_state_in_10_1_2 ^ port_key_10_1_2);
  assign port_state_out_10_1_3 = (port_state_in_10_1_3 ^ port_key_10_1_3);
  assign port_state_out_10_1_4 = (port_state_in_10_1_4 ^ port_key_10_1_4);
  assign port_state_out_10_1_5 = (port_state_in_10_1_5 ^ port_key_10_1_5);
  assign port_state_out_10_1_6 = (port_state_in_10_1_6 ^ port_key_10_1_6);
  assign port_state_out_10_1_7 = (port_state_in_10_1_7 ^ port_key_10_1_7);
  assign port_state_out_10_2_0 = (port_state_in_10_2_0 ^ port_key_10_2_0);
  assign port_state_out_10_2_1 = (port_state_in_10_2_1 ^ port_key_10_2_1);
  assign port_state_out_10_2_2 = (port_state_in_10_2_2 ^ port_key_10_2_2);
  assign port_state_out_10_2_3 = (port_state_in_10_2_3 ^ port_key_10_2_3);
  assign port_state_out_10_2_4 = (port_state_in_10_2_4 ^ port_key_10_2_4);
  assign port_state_out_10_2_5 = (port_state_in_10_2_5 ^ port_key_10_2_5);
  assign port_state_out_10_2_6 = (port_state_in_10_2_6 ^ port_key_10_2_6);
  assign port_state_out_10_2_7 = (port_state_in_10_2_7 ^ port_key_10_2_7);
  assign port_state_out_10_3_0 = (port_state_in_10_3_0 ^ port_key_10_3_0);
  assign port_state_out_10_3_1 = (port_state_in_10_3_1 ^ port_key_10_3_1);
  assign port_state_out_10_3_2 = (port_state_in_10_3_2 ^ port_key_10_3_2);
  assign port_state_out_10_3_3 = (port_state_in_10_3_3 ^ port_key_10_3_3);
  assign port_state_out_10_3_4 = (port_state_in_10_3_4 ^ port_key_10_3_4);
  assign port_state_out_10_3_5 = (port_state_in_10_3_5 ^ port_key_10_3_5);
  assign port_state_out_10_3_6 = (port_state_in_10_3_6 ^ port_key_10_3_6);
  assign port_state_out_10_3_7 = (port_state_in_10_3_7 ^ port_key_10_3_7);
  assign port_state_out_11_0_0 = (port_state_in_11_0_0 ^ port_key_11_0_0);
  assign port_state_out_11_0_1 = (port_state_in_11_0_1 ^ port_key_11_0_1);
  assign port_state_out_11_0_2 = (port_state_in_11_0_2 ^ port_key_11_0_2);
  assign port_state_out_11_0_3 = (port_state_in_11_0_3 ^ port_key_11_0_3);
  assign port_state_out_11_0_4 = (port_state_in_11_0_4 ^ port_key_11_0_4);
  assign port_state_out_11_0_5 = (port_state_in_11_0_5 ^ port_key_11_0_5);
  assign port_state_out_11_0_6 = (port_state_in_11_0_6 ^ port_key_11_0_6);
  assign port_state_out_11_0_7 = (port_state_in_11_0_7 ^ port_key_11_0_7);
  assign port_state_out_11_1_0 = (port_state_in_11_1_0 ^ port_key_11_1_0);
  assign port_state_out_11_1_1 = (port_state_in_11_1_1 ^ port_key_11_1_1);
  assign port_state_out_11_1_2 = (port_state_in_11_1_2 ^ port_key_11_1_2);
  assign port_state_out_11_1_3 = (port_state_in_11_1_3 ^ port_key_11_1_3);
  assign port_state_out_11_1_4 = (port_state_in_11_1_4 ^ port_key_11_1_4);
  assign port_state_out_11_1_5 = (port_state_in_11_1_5 ^ port_key_11_1_5);
  assign port_state_out_11_1_6 = (port_state_in_11_1_6 ^ port_key_11_1_6);
  assign port_state_out_11_1_7 = (port_state_in_11_1_7 ^ port_key_11_1_7);
  assign port_state_out_11_2_0 = (port_state_in_11_2_0 ^ port_key_11_2_0);
  assign port_state_out_11_2_1 = (port_state_in_11_2_1 ^ port_key_11_2_1);
  assign port_state_out_11_2_2 = (port_state_in_11_2_2 ^ port_key_11_2_2);
  assign port_state_out_11_2_3 = (port_state_in_11_2_3 ^ port_key_11_2_3);
  assign port_state_out_11_2_4 = (port_state_in_11_2_4 ^ port_key_11_2_4);
  assign port_state_out_11_2_5 = (port_state_in_11_2_5 ^ port_key_11_2_5);
  assign port_state_out_11_2_6 = (port_state_in_11_2_6 ^ port_key_11_2_6);
  assign port_state_out_11_2_7 = (port_state_in_11_2_7 ^ port_key_11_2_7);
  assign port_state_out_11_3_0 = (port_state_in_11_3_0 ^ port_key_11_3_0);
  assign port_state_out_11_3_1 = (port_state_in_11_3_1 ^ port_key_11_3_1);
  assign port_state_out_11_3_2 = (port_state_in_11_3_2 ^ port_key_11_3_2);
  assign port_state_out_11_3_3 = (port_state_in_11_3_3 ^ port_key_11_3_3);
  assign port_state_out_11_3_4 = (port_state_in_11_3_4 ^ port_key_11_3_4);
  assign port_state_out_11_3_5 = (port_state_in_11_3_5 ^ port_key_11_3_5);
  assign port_state_out_11_3_6 = (port_state_in_11_3_6 ^ port_key_11_3_6);
  assign port_state_out_11_3_7 = (port_state_in_11_3_7 ^ port_key_11_3_7);
  assign port_state_out_12_0_0 = (port_state_in_12_0_0 ^ port_key_12_0_0);
  assign port_state_out_12_0_1 = (port_state_in_12_0_1 ^ port_key_12_0_1);
  assign port_state_out_12_0_2 = (port_state_in_12_0_2 ^ port_key_12_0_2);
  assign port_state_out_12_0_3 = (port_state_in_12_0_3 ^ port_key_12_0_3);
  assign port_state_out_12_0_4 = (port_state_in_12_0_4 ^ port_key_12_0_4);
  assign port_state_out_12_0_5 = (port_state_in_12_0_5 ^ port_key_12_0_5);
  assign port_state_out_12_0_6 = (port_state_in_12_0_6 ^ port_key_12_0_6);
  assign port_state_out_12_0_7 = (port_state_in_12_0_7 ^ port_key_12_0_7);
  assign port_state_out_12_1_0 = (port_state_in_12_1_0 ^ port_key_12_1_0);
  assign port_state_out_12_1_1 = (port_state_in_12_1_1 ^ port_key_12_1_1);
  assign port_state_out_12_1_2 = (port_state_in_12_1_2 ^ port_key_12_1_2);
  assign port_state_out_12_1_3 = (port_state_in_12_1_3 ^ port_key_12_1_3);
  assign port_state_out_12_1_4 = (port_state_in_12_1_4 ^ port_key_12_1_4);
  assign port_state_out_12_1_5 = (port_state_in_12_1_5 ^ port_key_12_1_5);
  assign port_state_out_12_1_6 = (port_state_in_12_1_6 ^ port_key_12_1_6);
  assign port_state_out_12_1_7 = (port_state_in_12_1_7 ^ port_key_12_1_7);
  assign port_state_out_12_2_0 = (port_state_in_12_2_0 ^ port_key_12_2_0);
  assign port_state_out_12_2_1 = (port_state_in_12_2_1 ^ port_key_12_2_1);
  assign port_state_out_12_2_2 = (port_state_in_12_2_2 ^ port_key_12_2_2);
  assign port_state_out_12_2_3 = (port_state_in_12_2_3 ^ port_key_12_2_3);
  assign port_state_out_12_2_4 = (port_state_in_12_2_4 ^ port_key_12_2_4);
  assign port_state_out_12_2_5 = (port_state_in_12_2_5 ^ port_key_12_2_5);
  assign port_state_out_12_2_6 = (port_state_in_12_2_6 ^ port_key_12_2_6);
  assign port_state_out_12_2_7 = (port_state_in_12_2_7 ^ port_key_12_2_7);
  assign port_state_out_12_3_0 = (port_state_in_12_3_0 ^ port_key_12_3_0);
  assign port_state_out_12_3_1 = (port_state_in_12_3_1 ^ port_key_12_3_1);
  assign port_state_out_12_3_2 = (port_state_in_12_3_2 ^ port_key_12_3_2);
  assign port_state_out_12_3_3 = (port_state_in_12_3_3 ^ port_key_12_3_3);
  assign port_state_out_12_3_4 = (port_state_in_12_3_4 ^ port_key_12_3_4);
  assign port_state_out_12_3_5 = (port_state_in_12_3_5 ^ port_key_12_3_5);
  assign port_state_out_12_3_6 = (port_state_in_12_3_6 ^ port_key_12_3_6);
  assign port_state_out_12_3_7 = (port_state_in_12_3_7 ^ port_key_12_3_7);
  assign port_state_out_13_0_0 = (port_state_in_13_0_0 ^ port_key_13_0_0);
  assign port_state_out_13_0_1 = (port_state_in_13_0_1 ^ port_key_13_0_1);
  assign port_state_out_13_0_2 = (port_state_in_13_0_2 ^ port_key_13_0_2);
  assign port_state_out_13_0_3 = (port_state_in_13_0_3 ^ port_key_13_0_3);
  assign port_state_out_13_0_4 = (port_state_in_13_0_4 ^ port_key_13_0_4);
  assign port_state_out_13_0_5 = (port_state_in_13_0_5 ^ port_key_13_0_5);
  assign port_state_out_13_0_6 = (port_state_in_13_0_6 ^ port_key_13_0_6);
  assign port_state_out_13_0_7 = (port_state_in_13_0_7 ^ port_key_13_0_7);
  assign port_state_out_13_1_0 = (port_state_in_13_1_0 ^ port_key_13_1_0);
  assign port_state_out_13_1_1 = (port_state_in_13_1_1 ^ port_key_13_1_1);
  assign port_state_out_13_1_2 = (port_state_in_13_1_2 ^ port_key_13_1_2);
  assign port_state_out_13_1_3 = (port_state_in_13_1_3 ^ port_key_13_1_3);
  assign port_state_out_13_1_4 = (port_state_in_13_1_4 ^ port_key_13_1_4);
  assign port_state_out_13_1_5 = (port_state_in_13_1_5 ^ port_key_13_1_5);
  assign port_state_out_13_1_6 = (port_state_in_13_1_6 ^ port_key_13_1_6);
  assign port_state_out_13_1_7 = (port_state_in_13_1_7 ^ port_key_13_1_7);
  assign port_state_out_13_2_0 = (port_state_in_13_2_0 ^ port_key_13_2_0);
  assign port_state_out_13_2_1 = (port_state_in_13_2_1 ^ port_key_13_2_1);
  assign port_state_out_13_2_2 = (port_state_in_13_2_2 ^ port_key_13_2_2);
  assign port_state_out_13_2_3 = (port_state_in_13_2_3 ^ port_key_13_2_3);
  assign port_state_out_13_2_4 = (port_state_in_13_2_4 ^ port_key_13_2_4);
  assign port_state_out_13_2_5 = (port_state_in_13_2_5 ^ port_key_13_2_5);
  assign port_state_out_13_2_6 = (port_state_in_13_2_6 ^ port_key_13_2_6);
  assign port_state_out_13_2_7 = (port_state_in_13_2_7 ^ port_key_13_2_7);
  assign port_state_out_13_3_0 = (port_state_in_13_3_0 ^ port_key_13_3_0);
  assign port_state_out_13_3_1 = (port_state_in_13_3_1 ^ port_key_13_3_1);
  assign port_state_out_13_3_2 = (port_state_in_13_3_2 ^ port_key_13_3_2);
  assign port_state_out_13_3_3 = (port_state_in_13_3_3 ^ port_key_13_3_3);
  assign port_state_out_13_3_4 = (port_state_in_13_3_4 ^ port_key_13_3_4);
  assign port_state_out_13_3_5 = (port_state_in_13_3_5 ^ port_key_13_3_5);
  assign port_state_out_13_3_6 = (port_state_in_13_3_6 ^ port_key_13_3_6);
  assign port_state_out_13_3_7 = (port_state_in_13_3_7 ^ port_key_13_3_7);
  assign port_state_out_14_0_0 = (port_state_in_14_0_0 ^ port_key_14_0_0);
  assign port_state_out_14_0_1 = (port_state_in_14_0_1 ^ port_key_14_0_1);
  assign port_state_out_14_0_2 = (port_state_in_14_0_2 ^ port_key_14_0_2);
  assign port_state_out_14_0_3 = (port_state_in_14_0_3 ^ port_key_14_0_3);
  assign port_state_out_14_0_4 = (port_state_in_14_0_4 ^ port_key_14_0_4);
  assign port_state_out_14_0_5 = (port_state_in_14_0_5 ^ port_key_14_0_5);
  assign port_state_out_14_0_6 = (port_state_in_14_0_6 ^ port_key_14_0_6);
  assign port_state_out_14_0_7 = (port_state_in_14_0_7 ^ port_key_14_0_7);
  assign port_state_out_14_1_0 = (port_state_in_14_1_0 ^ port_key_14_1_0);
  assign port_state_out_14_1_1 = (port_state_in_14_1_1 ^ port_key_14_1_1);
  assign port_state_out_14_1_2 = (port_state_in_14_1_2 ^ port_key_14_1_2);
  assign port_state_out_14_1_3 = (port_state_in_14_1_3 ^ port_key_14_1_3);
  assign port_state_out_14_1_4 = (port_state_in_14_1_4 ^ port_key_14_1_4);
  assign port_state_out_14_1_5 = (port_state_in_14_1_5 ^ port_key_14_1_5);
  assign port_state_out_14_1_6 = (port_state_in_14_1_6 ^ port_key_14_1_6);
  assign port_state_out_14_1_7 = (port_state_in_14_1_7 ^ port_key_14_1_7);
  assign port_state_out_14_2_0 = (port_state_in_14_2_0 ^ port_key_14_2_0);
  assign port_state_out_14_2_1 = (port_state_in_14_2_1 ^ port_key_14_2_1);
  assign port_state_out_14_2_2 = (port_state_in_14_2_2 ^ port_key_14_2_2);
  assign port_state_out_14_2_3 = (port_state_in_14_2_3 ^ port_key_14_2_3);
  assign port_state_out_14_2_4 = (port_state_in_14_2_4 ^ port_key_14_2_4);
  assign port_state_out_14_2_5 = (port_state_in_14_2_5 ^ port_key_14_2_5);
  assign port_state_out_14_2_6 = (port_state_in_14_2_6 ^ port_key_14_2_6);
  assign port_state_out_14_2_7 = (port_state_in_14_2_7 ^ port_key_14_2_7);
  assign port_state_out_14_3_0 = (port_state_in_14_3_0 ^ port_key_14_3_0);
  assign port_state_out_14_3_1 = (port_state_in_14_3_1 ^ port_key_14_3_1);
  assign port_state_out_14_3_2 = (port_state_in_14_3_2 ^ port_key_14_3_2);
  assign port_state_out_14_3_3 = (port_state_in_14_3_3 ^ port_key_14_3_3);
  assign port_state_out_14_3_4 = (port_state_in_14_3_4 ^ port_key_14_3_4);
  assign port_state_out_14_3_5 = (port_state_in_14_3_5 ^ port_key_14_3_5);
  assign port_state_out_14_3_6 = (port_state_in_14_3_6 ^ port_key_14_3_6);
  assign port_state_out_14_3_7 = (port_state_in_14_3_7 ^ port_key_14_3_7);
  assign port_state_out_15_0_0 = (port_state_in_15_0_0 ^ port_key_15_0_0);
  assign port_state_out_15_0_1 = (port_state_in_15_0_1 ^ port_key_15_0_1);
  assign port_state_out_15_0_2 = (port_state_in_15_0_2 ^ port_key_15_0_2);
  assign port_state_out_15_0_3 = (port_state_in_15_0_3 ^ port_key_15_0_3);
  assign port_state_out_15_0_4 = (port_state_in_15_0_4 ^ port_key_15_0_4);
  assign port_state_out_15_0_5 = (port_state_in_15_0_5 ^ port_key_15_0_5);
  assign port_state_out_15_0_6 = (port_state_in_15_0_6 ^ port_key_15_0_6);
  assign port_state_out_15_0_7 = (port_state_in_15_0_7 ^ port_key_15_0_7);
  assign port_state_out_15_1_0 = (port_state_in_15_1_0 ^ port_key_15_1_0);
  assign port_state_out_15_1_1 = (port_state_in_15_1_1 ^ port_key_15_1_1);
  assign port_state_out_15_1_2 = (port_state_in_15_1_2 ^ port_key_15_1_2);
  assign port_state_out_15_1_3 = (port_state_in_15_1_3 ^ port_key_15_1_3);
  assign port_state_out_15_1_4 = (port_state_in_15_1_4 ^ port_key_15_1_4);
  assign port_state_out_15_1_5 = (port_state_in_15_1_5 ^ port_key_15_1_5);
  assign port_state_out_15_1_6 = (port_state_in_15_1_6 ^ port_key_15_1_6);
  assign port_state_out_15_1_7 = (port_state_in_15_1_7 ^ port_key_15_1_7);
  assign port_state_out_15_2_0 = (port_state_in_15_2_0 ^ port_key_15_2_0);
  assign port_state_out_15_2_1 = (port_state_in_15_2_1 ^ port_key_15_2_1);
  assign port_state_out_15_2_2 = (port_state_in_15_2_2 ^ port_key_15_2_2);
  assign port_state_out_15_2_3 = (port_state_in_15_2_3 ^ port_key_15_2_3);
  assign port_state_out_15_2_4 = (port_state_in_15_2_4 ^ port_key_15_2_4);
  assign port_state_out_15_2_5 = (port_state_in_15_2_5 ^ port_key_15_2_5);
  assign port_state_out_15_2_6 = (port_state_in_15_2_6 ^ port_key_15_2_6);
  assign port_state_out_15_2_7 = (port_state_in_15_2_7 ^ port_key_15_2_7);
  assign port_state_out_15_3_0 = (port_state_in_15_3_0 ^ port_key_15_3_0);
  assign port_state_out_15_3_1 = (port_state_in_15_3_1 ^ port_key_15_3_1);
  assign port_state_out_15_3_2 = (port_state_in_15_3_2 ^ port_key_15_3_2);
  assign port_state_out_15_3_3 = (port_state_in_15_3_3 ^ port_key_15_3_3);
  assign port_state_out_15_3_4 = (port_state_in_15_3_4 ^ port_key_15_3_4);
  assign port_state_out_15_3_5 = (port_state_in_15_3_5 ^ port_key_15_3_5);
  assign port_state_out_15_3_6 = (port_state_in_15_3_6 ^ port_key_15_3_6);
  assign port_state_out_15_3_7 = (port_state_in_15_3_7 ^ port_key_15_3_7);

endmodule

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

//Mul3 replaced by Mul3

//Mul2 replaced by Mul2

module Mul3 (
  input      [2:0]    port_byte_in_0,
  input      [2:0]    port_byte_in_1,
  input      [2:0]    port_byte_in_2,
  input      [2:0]    port_byte_in_3,
  input      [2:0]    port_byte_in_4,
  input      [2:0]    port_byte_in_5,
  input      [2:0]    port_byte_in_6,
  input      [2:0]    port_byte_in_7,
  output     [2:0]    port_byte_out_0,
  output     [2:0]    port_byte_out_1,
  output     [2:0]    port_byte_out_2,
  output     [2:0]    port_byte_out_3,
  output     [2:0]    port_byte_out_4,
  output     [2:0]    port_byte_out_5,
  output     [2:0]    port_byte_out_6,
  output     [2:0]    port_byte_out_7
);


  assign port_byte_out_7 = (port_byte_in_7 ^ port_byte_in_6);
  assign port_byte_out_6 = (port_byte_in_6 ^ port_byte_in_5);
  assign port_byte_out_5 = (port_byte_in_5 ^ port_byte_in_4);
  assign port_byte_out_4 = ((port_byte_in_7 ^ port_byte_in_4) ^ port_byte_in_3);
  assign port_byte_out_3 = ((port_byte_in_7 ^ port_byte_in_3) ^ port_byte_in_2);
  assign port_byte_out_2 = (port_byte_in_2 ^ port_byte_in_1);
  assign port_byte_out_1 = ((port_byte_in_7 ^ port_byte_in_1) ^ port_byte_in_0);
  assign port_byte_out_0 = (port_byte_in_7 ^ port_byte_in_0);

endmodule

module Mul2 (
  input      [2:0]    port_byte_in_0,
  input      [2:0]    port_byte_in_1,
  input      [2:0]    port_byte_in_2,
  input      [2:0]    port_byte_in_3,
  input      [2:0]    port_byte_in_4,
  input      [2:0]    port_byte_in_5,
  input      [2:0]    port_byte_in_6,
  input      [2:0]    port_byte_in_7,
  output     [2:0]    port_byte_out_0,
  output     [2:0]    port_byte_out_1,
  output     [2:0]    port_byte_out_2,
  output     [2:0]    port_byte_out_3,
  output     [2:0]    port_byte_out_4,
  output     [2:0]    port_byte_out_5,
  output     [2:0]    port_byte_out_6,
  output     [2:0]    port_byte_out_7
);


  assign port_byte_out_7 = port_byte_in_6;
  assign port_byte_out_6 = port_byte_in_5;
  assign port_byte_out_5 = port_byte_in_4;
  assign port_byte_out_4 = (port_byte_in_7 ^ port_byte_in_3);
  assign port_byte_out_3 = (port_byte_in_7 ^ port_byte_in_2);
  assign port_byte_out_2 = port_byte_in_1;
  assign port_byte_out_1 = (port_byte_in_7 ^ port_byte_in_0);
  assign port_byte_out_0 = port_byte_in_7;

endmodule

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_Inv_TI replaced by Addition_Inv_TI

module Addition_Inv_TI (
  input      [2:0]    port_x0_0,
  input      [2:0]    port_x0_1,
  input      [2:0]    port_x0_2,
  input      [2:0]    port_x0_3,
  input      [2:0]    port_x1_0,
  input      [2:0]    port_x1_1,
  input      [2:0]    port_x1_2,
  input      [2:0]    port_x1_3,
  output reg [2:0]    port_y_0,
  output reg [2:0]    port_y_1,
  output reg [2:0]    port_y_2,
  output reg [2:0]    port_y_3
);


  always @(*) begin
    port_y_0[0] = (! (port_x0_0[0] ^ port_x1_0[0]));
    port_y_0[1] = (! (port_x0_0[1] ^ port_x1_0[1]));
    port_y_0[2] = (! (port_x0_0[2] ^ port_x1_0[2]));
  end

  always @(*) begin
    port_y_1[0] = (port_x0_1[0] ^ port_x1_1[0]);
    port_y_1[1] = (port_x0_1[1] ^ port_x1_1[1]);
    port_y_1[2] = (port_x0_1[2] ^ port_x1_1[2]);
  end

  always @(*) begin
    port_y_2[0] = (port_x0_2[0] ^ port_x1_2[0]);
    port_y_2[1] = (port_x0_2[1] ^ port_x1_2[1]);
    port_y_2[2] = (port_x0_2[2] ^ port_x1_2[2]);
  end

  always @(*) begin
    port_y_3[0] = (port_x0_3[0] ^ port_x1_3[0]);
    port_y_3[1] = (port_x0_3[1] ^ port_x1_3[1]);
    port_y_3[2] = (port_x0_3[2] ^ port_x1_3[2]);
  end


endmodule

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

//Multiplication_TI_noReg replaced by Multiplication_TI_noReg

module Multiplication_TI_noReg (
  input      [2:0]    port_x0_0,
  input      [2:0]    port_x0_1,
  input      [2:0]    port_x0_2,
  input      [2:0]    port_x0_3,
  input      [2:0]    port_x1_0,
  input      [2:0]    port_x1_1,
  input      [2:0]    port_x1_2,
  input      [2:0]    port_x1_3,
  output     [2:0]    port_y_0,
  output     [2:0]    port_y_1,
  output     [2:0]    port_y_2,
  output     [2:0]    port_y_3
);

  reg        [2:0]    _zz_port_y_0;
  reg        [2:0]    _zz_port_y_1;
  reg        [2:0]    _zz_port_y_2;
  reg        [2:0]    _zz_port_y_3;

  always @(*) begin
    _zz_port_y_0[0] = (((((port_x0_1[0] ^ port_x0_2[0]) ^ port_x0_3[0]) && (port_x1_1[0] ^ port_x1_2[0])) ^ port_x1_3[0]) ^ port_x1_2[0]);
    _zz_port_y_0[1] = (((((port_x0_1[1] ^ port_x0_2[1]) ^ port_x0_3[1]) && (port_x1_1[1] ^ port_x1_2[1])) ^ port_x1_3[1]) ^ port_x1_2[1]);
    _zz_port_y_0[2] = (((((port_x0_1[2] ^ port_x0_2[2]) ^ port_x0_3[2]) && (port_x1_1[2] ^ port_x1_2[2])) ^ port_x1_3[2]) ^ port_x1_2[2]);
  end

  always @(*) begin
    _zz_port_y_1[0] = ((((port_x0_0[0] ^ port_x0_2[0]) && (port_x1_0[0] ^ port_x1_3[0])) ^ (port_x0_0[0] && port_x1_2[0])) ^ port_x0_3[0]);
    _zz_port_y_1[1] = ((((port_x0_0[1] ^ port_x0_2[1]) && (port_x1_0[1] ^ port_x1_3[1])) ^ (port_x0_0[1] && port_x1_2[1])) ^ port_x0_3[1]);
    _zz_port_y_1[2] = ((((port_x0_0[2] ^ port_x0_2[2]) && (port_x1_0[2] ^ port_x1_3[2])) ^ (port_x0_0[2] && port_x1_2[2])) ^ port_x0_3[2]);
  end

  always @(*) begin
    _zz_port_y_2[0] = ((((port_x0_1[0] ^ port_x0_3[0]) && (port_x1_0[0] ^ port_x1_3[0])) ^ port_x0_3[0]) ^ port_x1_3[0]);
    _zz_port_y_2[1] = ((((port_x0_1[1] ^ port_x0_3[1]) && (port_x1_0[1] ^ port_x1_3[1])) ^ port_x0_3[1]) ^ port_x1_3[1]);
    _zz_port_y_2[2] = ((((port_x0_1[2] ^ port_x0_3[2]) && (port_x1_0[2] ^ port_x1_3[2])) ^ port_x0_3[2]) ^ port_x1_3[2]);
  end

  always @(*) begin
    _zz_port_y_3[0] = ((port_x0_0[0] && port_x1_1[0]) ^ port_x1_2[0]);
    _zz_port_y_3[1] = ((port_x0_0[1] && port_x1_1[1]) ^ port_x1_2[1]);
    _zz_port_y_3[2] = ((port_x0_0[2] && port_x1_1[2]) ^ port_x1_2[2]);
  end

  assign port_y_0 = _zz_port_y_0;
  assign port_y_1 = _zz_port_y_1;
  assign port_y_2 = _zz_port_y_2;
  assign port_y_3 = _zz_port_y_3;

endmodule

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

//Multiplication_TI replaced by Multiplication_TI

module Multiplication_TI (
  input      [2:0]    port_x0_0,
  input      [2:0]    port_x0_1,
  input      [2:0]    port_x0_2,
  input      [2:0]    port_x0_3,
  input      [2:0]    port_x1_0,
  input      [2:0]    port_x1_1,
  input      [2:0]    port_x1_2,
  input      [2:0]    port_x1_3,
  output     [2:0]    port_y_0,
  output     [2:0]    port_y_1,
  output     [2:0]    port_y_2,
  output     [2:0]    port_y_3,
  input               clk,
  input               reset
);

  wire                majority_4608_port_o;
  wire                majority_4609_port_o;
  wire                majority_4610_port_o;
  wire                majority_4611_port_o;
  wire                majority_4612_port_o;
  wire                majority_4613_port_o;
  wire                majority_4614_port_o;
  wire                majority_4615_port_o;
  wire                majority_4616_port_o;
  wire                majority_4617_port_o;
  wire                majority_4618_port_o;
  wire                majority_4619_port_o;
  reg        [2:0]    _zz_port_i;
  reg        [2:0]    _zz_port_i_1;
  reg        [2:0]    _zz_port_i_2;
  reg        [2:0]    _zz_port_i_3;
  reg        [2:0]    _zz_port_y_0;
  reg        [2:0]    _zz_port_y_1;
  reg        [2:0]    _zz_port_y_2;
  reg        [2:0]    _zz_port_y_3;

  Majority majority_4608 (
    .port_i (_zz_port_i[2:0]     ), //i
    .port_o (majority_4608_port_o)  //o
  );
  Majority majority_4609 (
    .port_i (_zz_port_i_1[2:0]   ), //i
    .port_o (majority_4609_port_o)  //o
  );
  Majority majority_4610 (
    .port_i (_zz_port_i_2[2:0]   ), //i
    .port_o (majority_4610_port_o)  //o
  );
  Majority majority_4611 (
    .port_i (_zz_port_i_3[2:0]   ), //i
    .port_o (majority_4611_port_o)  //o
  );
  Majority majority_4612 (
    .port_i (_zz_port_i[2:0]     ), //i
    .port_o (majority_4612_port_o)  //o
  );
  Majority majority_4613 (
    .port_i (_zz_port_i_1[2:0]   ), //i
    .port_o (majority_4613_port_o)  //o
  );
  Majority majority_4614 (
    .port_i (_zz_port_i_2[2:0]   ), //i
    .port_o (majority_4614_port_o)  //o
  );
  Majority majority_4615 (
    .port_i (_zz_port_i_3[2:0]   ), //i
    .port_o (majority_4615_port_o)  //o
  );
  Majority majority_4616 (
    .port_i (_zz_port_i[2:0]     ), //i
    .port_o (majority_4616_port_o)  //o
  );
  Majority majority_4617 (
    .port_i (_zz_port_i_1[2:0]   ), //i
    .port_o (majority_4617_port_o)  //o
  );
  Majority majority_4618 (
    .port_i (_zz_port_i_2[2:0]   ), //i
    .port_o (majority_4618_port_o)  //o
  );
  Majority majority_4619 (
    .port_i (_zz_port_i_3[2:0]   ), //i
    .port_o (majority_4619_port_o)  //o
  );
  always @(*) begin
    _zz_port_i[0] = (((((port_x0_1[0] ^ port_x0_2[0]) ^ port_x0_3[0]) && (port_x1_1[0] ^ port_x1_2[0])) ^ port_x1_3[0]) ^ port_x1_2[0]);
    _zz_port_i[1] = (((((port_x0_1[1] ^ port_x0_2[1]) ^ port_x0_3[1]) && (port_x1_1[1] ^ port_x1_2[1])) ^ port_x1_3[1]) ^ port_x1_2[1]);
    _zz_port_i[2] = (((((port_x0_1[2] ^ port_x0_2[2]) ^ port_x0_3[2]) && (port_x1_1[2] ^ port_x1_2[2])) ^ port_x1_3[2]) ^ port_x1_2[2]);
  end

  always @(*) begin
    _zz_port_i_1[0] = ((((port_x0_0[0] ^ port_x0_2[0]) && (port_x1_0[0] ^ port_x1_3[0])) ^ (port_x0_0[0] && port_x1_2[0])) ^ port_x0_3[0]);
    _zz_port_i_1[1] = ((((port_x0_0[1] ^ port_x0_2[1]) && (port_x1_0[1] ^ port_x1_3[1])) ^ (port_x0_0[1] && port_x1_2[1])) ^ port_x0_3[1]);
    _zz_port_i_1[2] = ((((port_x0_0[2] ^ port_x0_2[2]) && (port_x1_0[2] ^ port_x1_3[2])) ^ (port_x0_0[2] && port_x1_2[2])) ^ port_x0_3[2]);
  end

  always @(*) begin
    _zz_port_i_2[0] = ((((port_x0_1[0] ^ port_x0_3[0]) && (port_x1_0[0] ^ port_x1_3[0])) ^ port_x0_3[0]) ^ port_x1_3[0]);
    _zz_port_i_2[1] = ((((port_x0_1[1] ^ port_x0_3[1]) && (port_x1_0[1] ^ port_x1_3[1])) ^ port_x0_3[1]) ^ port_x1_3[1]);
    _zz_port_i_2[2] = ((((port_x0_1[2] ^ port_x0_3[2]) && (port_x1_0[2] ^ port_x1_3[2])) ^ port_x0_3[2]) ^ port_x1_3[2]);
  end

  always @(*) begin
    _zz_port_i_3[0] = ((port_x0_0[0] && port_x1_1[0]) ^ port_x1_2[0]);
    _zz_port_i_3[1] = ((port_x0_0[1] && port_x1_1[1]) ^ port_x1_2[1]);
    _zz_port_i_3[2] = ((port_x0_0[2] && port_x1_1[2]) ^ port_x1_2[2]);
  end

  assign port_y_0 = _zz_port_y_0;
  assign port_y_1 = _zz_port_y_1;
  assign port_y_2 = _zz_port_y_2;
  assign port_y_3 = _zz_port_y_3;
  always @(posedge clk) begin
    _zz_port_y_0[0] <= majority_4608_port_o;
    _zz_port_y_1[0] <= majority_4609_port_o;
    _zz_port_y_2[0] <= majority_4610_port_o;
    _zz_port_y_3[0] <= majority_4611_port_o;
    _zz_port_y_0[1] <= majority_4612_port_o;
    _zz_port_y_1[1] <= majority_4613_port_o;
    _zz_port_y_2[1] <= majority_4614_port_o;
    _zz_port_y_3[1] <= majority_4615_port_o;
    _zz_port_y_0[2] <= majority_4616_port_o;
    _zz_port_y_1[2] <= majority_4617_port_o;
    _zz_port_y_2[2] <= majority_4618_port_o;
    _zz_port_y_3[2] <= majority_4619_port_o;
  end


endmodule

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

//Addition_TI replaced by Addition_TI

module Addition_TI (
  input      [2:0]    port_x0_0,
  input      [2:0]    port_x0_1,
  input      [2:0]    port_x0_2,
  input      [2:0]    port_x0_3,
  input      [2:0]    port_x1_0,
  input      [2:0]    port_x1_1,
  input      [2:0]    port_x1_2,
  input      [2:0]    port_x1_3,
  output reg [2:0]    port_y_0,
  output reg [2:0]    port_y_1,
  output reg [2:0]    port_y_2,
  output reg [2:0]    port_y_3
);


  always @(*) begin
    port_y_0[0] = (port_x0_0[0] ^ port_x1_0[0]);
    port_y_0[1] = (port_x0_0[1] ^ port_x1_0[1]);
    port_y_0[2] = (port_x0_0[2] ^ port_x1_0[2]);
  end

  always @(*) begin
    port_y_1[0] = (port_x0_1[0] ^ port_x1_1[0]);
    port_y_1[1] = (port_x0_1[1] ^ port_x1_1[1]);
    port_y_1[2] = (port_x0_1[2] ^ port_x1_1[2]);
  end

  always @(*) begin
    port_y_2[0] = (port_x0_2[0] ^ port_x1_2[0]);
    port_y_2[1] = (port_x0_2[1] ^ port_x1_2[1]);
    port_y_2[2] = (port_x0_2[2] ^ port_x1_2[2]);
  end

  always @(*) begin
    port_y_3[0] = (port_x0_3[0] ^ port_x1_3[0]);
    port_y_3[1] = (port_x0_3[1] ^ port_x1_3[1]);
    port_y_3[2] = (port_x0_3[2] ^ port_x1_3[2]);
  end


endmodule

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

//Majority replaced by Majority

module Majority (
  input      [2:0]    port_i,
  output              port_o
);

  wire       [2:0]    _zz_port_o;
  wire                _zz_port_o_1;
  wire                _zz_port_o_2;
  wire                _zz_port_o_3;

  assign _zz_port_o = port_i;
  assign _zz_port_o_1 = _zz_port_o[0];
  assign _zz_port_o_2 = _zz_port_o[1];
  assign _zz_port_o_3 = _zz_port_o[2];
  assign port_o = (((1'b0 || ((1'b1 && _zz_port_o_1) && _zz_port_o_2)) || ((1'b1 && _zz_port_o_1) && _zz_port_o_3)) || ((1'b1 && _zz_port_o_2) && _zz_port_o_3));

endmodule
